-- File created by Bench2VHDL
-- Name: s35932
-- File: bench/s35932.bench
-- Timestamp: 2019-05-21T22:08:29.492009
--
-- Original File
-- =============
--	# s35932
--	# 35 inputs
--	# 320 outputs
--	# 1728 D-type flipflops
--	# 3861 inverters
--	# 12204 gates (4032 ANDs + 7020 NANDs + 1152 ORs + 0 NORs)
--	
--	INPUT(DATA_0_31)
--	INPUT(DATA_0_30)
--	INPUT(DATA_0_29)
--	INPUT(DATA_0_28)
--	INPUT(DATA_0_27)
--	INPUT(DATA_0_26)
--	INPUT(DATA_0_25)
--	INPUT(DATA_0_24)
--	INPUT(DATA_0_23)
--	INPUT(DATA_0_22)
--	INPUT(DATA_0_21)
--	INPUT(DATA_0_20)
--	INPUT(DATA_0_19)
--	INPUT(DATA_0_18)
--	INPUT(DATA_0_17)
--	INPUT(DATA_0_16)
--	INPUT(DATA_0_15)
--	INPUT(DATA_0_14)
--	INPUT(DATA_0_13)
--	INPUT(DATA_0_12)
--	INPUT(DATA_0_11)
--	INPUT(DATA_0_10)
--	INPUT(DATA_0_9)
--	INPUT(DATA_0_8)
--	INPUT(DATA_0_7)
--	INPUT(DATA_0_6)
--	INPUT(DATA_0_5)
--	INPUT(DATA_0_4)
--	INPUT(DATA_0_3)
--	INPUT(DATA_0_2)
--	INPUT(DATA_0_1)
--	INPUT(DATA_0_0)
--	INPUT(RESET)
--	INPUT(TM1)
--	INPUT(TM0)
--	
--	OUTPUT(DATA_9_31)
--	OUTPUT(DATA_9_30)
--	OUTPUT(DATA_9_29)
--	OUTPUT(DATA_9_28)
--	OUTPUT(DATA_9_27)
--	OUTPUT(DATA_9_26)
--	OUTPUT(DATA_9_25)
--	OUTPUT(DATA_9_24)
--	OUTPUT(DATA_9_23)
--	OUTPUT(DATA_9_22)
--	OUTPUT(DATA_9_21)
--	OUTPUT(DATA_9_20)
--	OUTPUT(DATA_9_19)
--	OUTPUT(DATA_9_18)
--	OUTPUT(DATA_9_17)
--	OUTPUT(DATA_9_16)
--	OUTPUT(DATA_9_15)
--	OUTPUT(DATA_9_14)
--	OUTPUT(DATA_9_13)
--	OUTPUT(DATA_9_12)
--	OUTPUT(DATA_9_11)
--	OUTPUT(DATA_9_10)
--	OUTPUT(DATA_9_9)
--	OUTPUT(DATA_9_8)
--	OUTPUT(DATA_9_7)
--	OUTPUT(DATA_9_6)
--	OUTPUT(DATA_9_5)
--	OUTPUT(DATA_9_4)
--	OUTPUT(DATA_9_3)
--	OUTPUT(DATA_9_2)
--	OUTPUT(DATA_9_1)
--	OUTPUT(DATA_9_0)
--	OUTPUT(CRC_OUT_9_0)
--	OUTPUT(CRC_OUT_9_1)
--	OUTPUT(CRC_OUT_9_2)
--	OUTPUT(CRC_OUT_9_3)
--	OUTPUT(CRC_OUT_9_4)
--	OUTPUT(CRC_OUT_9_5)
--	OUTPUT(CRC_OUT_9_6)
--	OUTPUT(CRC_OUT_9_7)
--	OUTPUT(CRC_OUT_9_8)
--	OUTPUT(CRC_OUT_9_9)
--	OUTPUT(CRC_OUT_9_10)
--	OUTPUT(CRC_OUT_9_11)
--	OUTPUT(CRC_OUT_9_12)
--	OUTPUT(CRC_OUT_9_13)
--	OUTPUT(CRC_OUT_9_14)
--	OUTPUT(CRC_OUT_9_15)
--	OUTPUT(CRC_OUT_9_16)
--	OUTPUT(CRC_OUT_9_17)
--	OUTPUT(CRC_OUT_9_18)
--	OUTPUT(CRC_OUT_9_19)
--	OUTPUT(CRC_OUT_9_20)
--	OUTPUT(CRC_OUT_9_21)
--	OUTPUT(CRC_OUT_9_22)
--	OUTPUT(CRC_OUT_9_23)
--	OUTPUT(CRC_OUT_9_24)
--	OUTPUT(CRC_OUT_9_25)
--	OUTPUT(CRC_OUT_9_26)
--	OUTPUT(CRC_OUT_9_27)
--	OUTPUT(CRC_OUT_9_28)
--	OUTPUT(CRC_OUT_9_29)
--	OUTPUT(CRC_OUT_9_30)
--	OUTPUT(CRC_OUT_9_31)
--	OUTPUT(CRC_OUT_8_0)
--	OUTPUT(CRC_OUT_8_1)
--	OUTPUT(CRC_OUT_8_2)
--	OUTPUT(CRC_OUT_8_3)
--	OUTPUT(CRC_OUT_8_4)
--	OUTPUT(CRC_OUT_8_5)
--	OUTPUT(CRC_OUT_8_6)
--	OUTPUT(CRC_OUT_8_7)
--	OUTPUT(CRC_OUT_8_8)
--	OUTPUT(CRC_OUT_8_9)
--	OUTPUT(CRC_OUT_8_10)
--	OUTPUT(CRC_OUT_8_11)
--	OUTPUT(CRC_OUT_8_12)
--	OUTPUT(CRC_OUT_8_13)
--	OUTPUT(CRC_OUT_8_14)
--	OUTPUT(CRC_OUT_8_15)
--	OUTPUT(CRC_OUT_8_16)
--	OUTPUT(CRC_OUT_8_17)
--	OUTPUT(CRC_OUT_8_18)
--	OUTPUT(CRC_OUT_8_19)
--	OUTPUT(CRC_OUT_8_20)
--	OUTPUT(CRC_OUT_8_21)
--	OUTPUT(CRC_OUT_8_22)
--	OUTPUT(CRC_OUT_8_23)
--	OUTPUT(CRC_OUT_8_24)
--	OUTPUT(CRC_OUT_8_25)
--	OUTPUT(CRC_OUT_8_26)
--	OUTPUT(CRC_OUT_8_27)
--	OUTPUT(CRC_OUT_8_28)
--	OUTPUT(CRC_OUT_8_29)
--	OUTPUT(CRC_OUT_8_30)
--	OUTPUT(CRC_OUT_8_31)
--	OUTPUT(CRC_OUT_7_0)
--	OUTPUT(CRC_OUT_7_1)
--	OUTPUT(CRC_OUT_7_2)
--	OUTPUT(CRC_OUT_7_3)
--	OUTPUT(CRC_OUT_7_4)
--	OUTPUT(CRC_OUT_7_5)
--	OUTPUT(CRC_OUT_7_6)
--	OUTPUT(CRC_OUT_7_7)
--	OUTPUT(CRC_OUT_7_8)
--	OUTPUT(CRC_OUT_7_9)
--	OUTPUT(CRC_OUT_7_10)
--	OUTPUT(CRC_OUT_7_11)
--	OUTPUT(CRC_OUT_7_12)
--	OUTPUT(CRC_OUT_7_13)
--	OUTPUT(CRC_OUT_7_14)
--	OUTPUT(CRC_OUT_7_15)
--	OUTPUT(CRC_OUT_7_16)
--	OUTPUT(CRC_OUT_7_17)
--	OUTPUT(CRC_OUT_7_18)
--	OUTPUT(CRC_OUT_7_19)
--	OUTPUT(CRC_OUT_7_20)
--	OUTPUT(CRC_OUT_7_21)
--	OUTPUT(CRC_OUT_7_22)
--	OUTPUT(CRC_OUT_7_23)
--	OUTPUT(CRC_OUT_7_24)
--	OUTPUT(CRC_OUT_7_25)
--	OUTPUT(CRC_OUT_7_26)
--	OUTPUT(CRC_OUT_7_27)
--	OUTPUT(CRC_OUT_7_28)
--	OUTPUT(CRC_OUT_7_29)
--	OUTPUT(CRC_OUT_7_30)
--	OUTPUT(CRC_OUT_7_31)
--	OUTPUT(CRC_OUT_6_0)
--	OUTPUT(CRC_OUT_6_1)
--	OUTPUT(CRC_OUT_6_2)
--	OUTPUT(CRC_OUT_6_3)
--	OUTPUT(CRC_OUT_6_4)
--	OUTPUT(CRC_OUT_6_5)
--	OUTPUT(CRC_OUT_6_6)
--	OUTPUT(CRC_OUT_6_7)
--	OUTPUT(CRC_OUT_6_8)
--	OUTPUT(CRC_OUT_6_9)
--	OUTPUT(CRC_OUT_6_10)
--	OUTPUT(CRC_OUT_6_11)
--	OUTPUT(CRC_OUT_6_12)
--	OUTPUT(CRC_OUT_6_13)
--	OUTPUT(CRC_OUT_6_14)
--	OUTPUT(CRC_OUT_6_15)
--	OUTPUT(CRC_OUT_6_16)
--	OUTPUT(CRC_OUT_6_17)
--	OUTPUT(CRC_OUT_6_18)
--	OUTPUT(CRC_OUT_6_19)
--	OUTPUT(CRC_OUT_6_20)
--	OUTPUT(CRC_OUT_6_21)
--	OUTPUT(CRC_OUT_6_22)
--	OUTPUT(CRC_OUT_6_23)
--	OUTPUT(CRC_OUT_6_24)
--	OUTPUT(CRC_OUT_6_25)
--	OUTPUT(CRC_OUT_6_26)
--	OUTPUT(CRC_OUT_6_27)
--	OUTPUT(CRC_OUT_6_28)
--	OUTPUT(CRC_OUT_6_29)
--	OUTPUT(CRC_OUT_6_30)
--	OUTPUT(CRC_OUT_6_31)
--	OUTPUT(CRC_OUT_5_0)
--	OUTPUT(CRC_OUT_5_1)
--	OUTPUT(CRC_OUT_5_2)
--	OUTPUT(CRC_OUT_5_3)
--	OUTPUT(CRC_OUT_5_4)
--	OUTPUT(CRC_OUT_5_5)
--	OUTPUT(CRC_OUT_5_6)
--	OUTPUT(CRC_OUT_5_7)
--	OUTPUT(CRC_OUT_5_8)
--	OUTPUT(CRC_OUT_5_9)
--	OUTPUT(CRC_OUT_5_10)
--	OUTPUT(CRC_OUT_5_11)
--	OUTPUT(CRC_OUT_5_12)
--	OUTPUT(CRC_OUT_5_13)
--	OUTPUT(CRC_OUT_5_14)
--	OUTPUT(CRC_OUT_5_15)
--	OUTPUT(CRC_OUT_5_16)
--	OUTPUT(CRC_OUT_5_17)
--	OUTPUT(CRC_OUT_5_18)
--	OUTPUT(CRC_OUT_5_19)
--	OUTPUT(CRC_OUT_5_20)
--	OUTPUT(CRC_OUT_5_21)
--	OUTPUT(CRC_OUT_5_22)
--	OUTPUT(CRC_OUT_5_23)
--	OUTPUT(CRC_OUT_5_24)
--	OUTPUT(CRC_OUT_5_25)
--	OUTPUT(CRC_OUT_5_26)
--	OUTPUT(CRC_OUT_5_27)
--	OUTPUT(CRC_OUT_5_28)
--	OUTPUT(CRC_OUT_5_29)
--	OUTPUT(CRC_OUT_5_30)
--	OUTPUT(CRC_OUT_5_31)
--	OUTPUT(CRC_OUT_4_0)
--	OUTPUT(CRC_OUT_4_1)
--	OUTPUT(CRC_OUT_4_2)
--	OUTPUT(CRC_OUT_4_3)
--	OUTPUT(CRC_OUT_4_4)
--	OUTPUT(CRC_OUT_4_5)
--	OUTPUT(CRC_OUT_4_6)
--	OUTPUT(CRC_OUT_4_7)
--	OUTPUT(CRC_OUT_4_8)
--	OUTPUT(CRC_OUT_4_9)
--	OUTPUT(CRC_OUT_4_10)
--	OUTPUT(CRC_OUT_4_11)
--	OUTPUT(CRC_OUT_4_12)
--	OUTPUT(CRC_OUT_4_13)
--	OUTPUT(CRC_OUT_4_14)
--	OUTPUT(CRC_OUT_4_15)
--	OUTPUT(CRC_OUT_4_16)
--	OUTPUT(CRC_OUT_4_17)
--	OUTPUT(CRC_OUT_4_18)
--	OUTPUT(CRC_OUT_4_19)
--	OUTPUT(CRC_OUT_4_20)
--	OUTPUT(CRC_OUT_4_21)
--	OUTPUT(CRC_OUT_4_22)
--	OUTPUT(CRC_OUT_4_23)
--	OUTPUT(CRC_OUT_4_24)
--	OUTPUT(CRC_OUT_4_25)
--	OUTPUT(CRC_OUT_4_26)
--	OUTPUT(CRC_OUT_4_27)
--	OUTPUT(CRC_OUT_4_28)
--	OUTPUT(CRC_OUT_4_29)
--	OUTPUT(CRC_OUT_4_30)
--	OUTPUT(CRC_OUT_4_31)
--	OUTPUT(CRC_OUT_3_0)
--	OUTPUT(CRC_OUT_3_1)
--	OUTPUT(CRC_OUT_3_2)
--	OUTPUT(CRC_OUT_3_3)
--	OUTPUT(CRC_OUT_3_4)
--	OUTPUT(CRC_OUT_3_5)
--	OUTPUT(CRC_OUT_3_6)
--	OUTPUT(CRC_OUT_3_7)
--	OUTPUT(CRC_OUT_3_8)
--	OUTPUT(CRC_OUT_3_9)
--	OUTPUT(CRC_OUT_3_10)
--	OUTPUT(CRC_OUT_3_11)
--	OUTPUT(CRC_OUT_3_12)
--	OUTPUT(CRC_OUT_3_13)
--	OUTPUT(CRC_OUT_3_14)
--	OUTPUT(CRC_OUT_3_15)
--	OUTPUT(CRC_OUT_3_16)
--	OUTPUT(CRC_OUT_3_17)
--	OUTPUT(CRC_OUT_3_18)
--	OUTPUT(CRC_OUT_3_19)
--	OUTPUT(CRC_OUT_3_20)
--	OUTPUT(CRC_OUT_3_21)
--	OUTPUT(CRC_OUT_3_22)
--	OUTPUT(CRC_OUT_3_23)
--	OUTPUT(CRC_OUT_3_24)
--	OUTPUT(CRC_OUT_3_25)
--	OUTPUT(CRC_OUT_3_26)
--	OUTPUT(CRC_OUT_3_27)
--	OUTPUT(CRC_OUT_3_28)
--	OUTPUT(CRC_OUT_3_29)
--	OUTPUT(CRC_OUT_3_30)
--	OUTPUT(CRC_OUT_3_31)
--	OUTPUT(CRC_OUT_2_0)
--	OUTPUT(CRC_OUT_2_1)
--	OUTPUT(CRC_OUT_2_2)
--	OUTPUT(CRC_OUT_2_3)
--	OUTPUT(CRC_OUT_2_4)
--	OUTPUT(CRC_OUT_2_5)
--	OUTPUT(CRC_OUT_2_6)
--	OUTPUT(CRC_OUT_2_7)
--	OUTPUT(CRC_OUT_2_8)
--	OUTPUT(CRC_OUT_2_9)
--	OUTPUT(CRC_OUT_2_10)
--	OUTPUT(CRC_OUT_2_11)
--	OUTPUT(CRC_OUT_2_12)
--	OUTPUT(CRC_OUT_2_13)
--	OUTPUT(CRC_OUT_2_14)
--	OUTPUT(CRC_OUT_2_15)
--	OUTPUT(CRC_OUT_2_16)
--	OUTPUT(CRC_OUT_2_17)
--	OUTPUT(CRC_OUT_2_18)
--	OUTPUT(CRC_OUT_2_19)
--	OUTPUT(CRC_OUT_2_20)
--	OUTPUT(CRC_OUT_2_21)
--	OUTPUT(CRC_OUT_2_22)
--	OUTPUT(CRC_OUT_2_23)
--	OUTPUT(CRC_OUT_2_24)
--	OUTPUT(CRC_OUT_2_25)
--	OUTPUT(CRC_OUT_2_26)
--	OUTPUT(CRC_OUT_2_27)
--	OUTPUT(CRC_OUT_2_28)
--	OUTPUT(CRC_OUT_2_29)
--	OUTPUT(CRC_OUT_2_30)
--	OUTPUT(CRC_OUT_2_31)
--	OUTPUT(CRC_OUT_1_0)
--	OUTPUT(CRC_OUT_1_1)
--	OUTPUT(CRC_OUT_1_2)
--	OUTPUT(CRC_OUT_1_3)
--	OUTPUT(CRC_OUT_1_4)
--	OUTPUT(CRC_OUT_1_5)
--	OUTPUT(CRC_OUT_1_6)
--	OUTPUT(CRC_OUT_1_7)
--	OUTPUT(CRC_OUT_1_8)
--	OUTPUT(CRC_OUT_1_9)
--	OUTPUT(CRC_OUT_1_10)
--	OUTPUT(CRC_OUT_1_11)
--	OUTPUT(CRC_OUT_1_12)
--	OUTPUT(CRC_OUT_1_13)
--	OUTPUT(CRC_OUT_1_14)
--	OUTPUT(CRC_OUT_1_15)
--	OUTPUT(CRC_OUT_1_16)
--	OUTPUT(CRC_OUT_1_17)
--	OUTPUT(CRC_OUT_1_18)
--	OUTPUT(CRC_OUT_1_19)
--	OUTPUT(CRC_OUT_1_20)
--	OUTPUT(CRC_OUT_1_21)
--	OUTPUT(CRC_OUT_1_22)
--	OUTPUT(CRC_OUT_1_23)
--	OUTPUT(CRC_OUT_1_24)
--	OUTPUT(CRC_OUT_1_25)
--	OUTPUT(CRC_OUT_1_26)
--	OUTPUT(CRC_OUT_1_27)
--	OUTPUT(CRC_OUT_1_28)
--	OUTPUT(CRC_OUT_1_29)
--	OUTPUT(CRC_OUT_1_30)
--	OUTPUT(CRC_OUT_1_31)
--	
--	WX485 = DFF(WX484)
--	WX487 = DFF(WX486)
--	WX489 = DFF(WX488)
--	WX491 = DFF(WX490)
--	WX493 = DFF(WX492)
--	WX495 = DFF(WX494)
--	WX497 = DFF(WX496)
--	WX499 = DFF(WX498)
--	WX501 = DFF(WX500)
--	WX503 = DFF(WX502)
--	WX505 = DFF(WX504)
--	WX507 = DFF(WX506)
--	WX509 = DFF(WX508)
--	WX511 = DFF(WX510)
--	WX513 = DFF(WX512)
--	WX515 = DFF(WX514)
--	WX517 = DFF(WX516)
--	WX519 = DFF(WX518)
--	WX521 = DFF(WX520)
--	WX523 = DFF(WX522)
--	WX525 = DFF(WX524)
--	WX527 = DFF(WX526)
--	WX529 = DFF(WX528)
--	WX531 = DFF(WX530)
--	WX533 = DFF(WX532)
--	WX535 = DFF(WX534)
--	WX537 = DFF(WX536)
--	WX539 = DFF(WX538)
--	WX541 = DFF(WX540)
--	WX543 = DFF(WX542)
--	WX545 = DFF(WX544)
--	WX547 = DFF(WX546)
--	WX645 = DFF(WX644)
--	WX647 = DFF(WX646)
--	WX649 = DFF(WX648)
--	WX651 = DFF(WX650)
--	WX653 = DFF(WX652)
--	WX655 = DFF(WX654)
--	WX657 = DFF(WX656)
--	WX659 = DFF(WX658)
--	WX661 = DFF(WX660)
--	WX663 = DFF(WX662)
--	WX665 = DFF(WX664)
--	WX667 = DFF(WX666)
--	WX669 = DFF(WX668)
--	WX671 = DFF(WX670)
--	WX673 = DFF(WX672)
--	WX675 = DFF(WX674)
--	WX677 = DFF(WX676)
--	WX679 = DFF(WX678)
--	WX681 = DFF(WX680)
--	WX683 = DFF(WX682)
--	WX685 = DFF(WX684)
--	WX687 = DFF(WX686)
--	WX689 = DFF(WX688)
--	WX691 = DFF(WX690)
--	WX693 = DFF(WX692)
--	WX695 = DFF(WX694)
--	WX697 = DFF(WX696)
--	WX699 = DFF(WX698)
--	WX701 = DFF(WX700)
--	WX703 = DFF(WX702)
--	WX705 = DFF(WX704)
--	WX707 = DFF(WX706)
--	WX709 = DFF(WX708)
--	WX711 = DFF(WX710)
--	WX713 = DFF(WX712)
--	WX715 = DFF(WX714)
--	WX717 = DFF(WX716)
--	WX719 = DFF(WX718)
--	WX721 = DFF(WX720)
--	WX723 = DFF(WX722)
--	WX725 = DFF(WX724)
--	WX727 = DFF(WX726)
--	WX729 = DFF(WX728)
--	WX731 = DFF(WX730)
--	WX733 = DFF(WX732)
--	WX735 = DFF(WX734)
--	WX737 = DFF(WX736)
--	WX739 = DFF(WX738)
--	WX741 = DFF(WX740)
--	WX743 = DFF(WX742)
--	WX745 = DFF(WX744)
--	WX747 = DFF(WX746)
--	WX749 = DFF(WX748)
--	WX751 = DFF(WX750)
--	WX753 = DFF(WX752)
--	WX755 = DFF(WX754)
--	WX757 = DFF(WX756)
--	WX759 = DFF(WX758)
--	WX761 = DFF(WX760)
--	WX763 = DFF(WX762)
--	WX765 = DFF(WX764)
--	WX767 = DFF(WX766)
--	WX769 = DFF(WX768)
--	WX771 = DFF(WX770)
--	WX773 = DFF(WX772)
--	WX775 = DFF(WX774)
--	WX777 = DFF(WX776)
--	WX779 = DFF(WX778)
--	WX781 = DFF(WX780)
--	WX783 = DFF(WX782)
--	WX785 = DFF(WX784)
--	WX787 = DFF(WX786)
--	WX789 = DFF(WX788)
--	WX791 = DFF(WX790)
--	WX793 = DFF(WX792)
--	WX795 = DFF(WX794)
--	WX797 = DFF(WX796)
--	WX799 = DFF(WX798)
--	WX801 = DFF(WX800)
--	WX803 = DFF(WX802)
--	WX805 = DFF(WX804)
--	WX807 = DFF(WX806)
--	WX809 = DFF(WX808)
--	WX811 = DFF(WX810)
--	WX813 = DFF(WX812)
--	WX815 = DFF(WX814)
--	WX817 = DFF(WX816)
--	WX819 = DFF(WX818)
--	WX821 = DFF(WX820)
--	WX823 = DFF(WX822)
--	WX825 = DFF(WX824)
--	WX827 = DFF(WX826)
--	WX829 = DFF(WX828)
--	WX831 = DFF(WX830)
--	WX833 = DFF(WX832)
--	WX835 = DFF(WX834)
--	WX837 = DFF(WX836)
--	WX839 = DFF(WX838)
--	WX841 = DFF(WX840)
--	WX843 = DFF(WX842)
--	WX845 = DFF(WX844)
--	WX847 = DFF(WX846)
--	WX849 = DFF(WX848)
--	WX851 = DFF(WX850)
--	WX853 = DFF(WX852)
--	WX855 = DFF(WX854)
--	WX857 = DFF(WX856)
--	WX859 = DFF(WX858)
--	WX861 = DFF(WX860)
--	WX863 = DFF(WX862)
--	WX865 = DFF(WX864)
--	WX867 = DFF(WX866)
--	WX869 = DFF(WX868)
--	WX871 = DFF(WX870)
--	WX873 = DFF(WX872)
--	WX875 = DFF(WX874)
--	WX877 = DFF(WX876)
--	WX879 = DFF(WX878)
--	WX881 = DFF(WX880)
--	WX883 = DFF(WX882)
--	WX885 = DFF(WX884)
--	WX887 = DFF(WX886)
--	WX889 = DFF(WX888)
--	WX891 = DFF(WX890)
--	WX893 = DFF(WX892)
--	WX895 = DFF(WX894)
--	WX897 = DFF(WX896)
--	WX899 = DFF(WX898)
--	CRC_OUT_9_0 = DFF(WX1264)
--	CRC_OUT_9_1 = DFF(WX1266)
--	CRC_OUT_9_2 = DFF(WX1268)
--	CRC_OUT_9_3 = DFF(WX1270)
--	CRC_OUT_9_4 = DFF(WX1272)
--	CRC_OUT_9_5 = DFF(WX1274)
--	CRC_OUT_9_6 = DFF(WX1276)
--	CRC_OUT_9_7 = DFF(WX1278)
--	CRC_OUT_9_8 = DFF(WX1280)
--	CRC_OUT_9_9 = DFF(WX1282)
--	CRC_OUT_9_10 = DFF(WX1284)
--	CRC_OUT_9_11 = DFF(WX1286)
--	CRC_OUT_9_12 = DFF(WX1288)
--	CRC_OUT_9_13 = DFF(WX1290)
--	CRC_OUT_9_14 = DFF(WX1292)
--	CRC_OUT_9_15 = DFF(WX1294)
--	CRC_OUT_9_16 = DFF(WX1296)
--	CRC_OUT_9_17 = DFF(WX1298)
--	CRC_OUT_9_18 = DFF(WX1300)
--	CRC_OUT_9_19 = DFF(WX1302)
--	CRC_OUT_9_20 = DFF(WX1304)
--	CRC_OUT_9_21 = DFF(WX1306)
--	CRC_OUT_9_22 = DFF(WX1308)
--	CRC_OUT_9_23 = DFF(WX1310)
--	CRC_OUT_9_24 = DFF(WX1312)
--	CRC_OUT_9_25 = DFF(WX1314)
--	CRC_OUT_9_26 = DFF(WX1316)
--	CRC_OUT_9_27 = DFF(WX1318)
--	CRC_OUT_9_28 = DFF(WX1320)
--	CRC_OUT_9_29 = DFF(WX1322)
--	CRC_OUT_9_30 = DFF(WX1324)
--	CRC_OUT_9_31 = DFF(WX1326)
--	WX1778 = DFF(WX1777)
--	WX1780 = DFF(WX1779)
--	WX1782 = DFF(WX1781)
--	WX1784 = DFF(WX1783)
--	WX1786 = DFF(WX1785)
--	WX1788 = DFF(WX1787)
--	WX1790 = DFF(WX1789)
--	WX1792 = DFF(WX1791)
--	WX1794 = DFF(WX1793)
--	WX1796 = DFF(WX1795)
--	WX1798 = DFF(WX1797)
--	WX1800 = DFF(WX1799)
--	WX1802 = DFF(WX1801)
--	WX1804 = DFF(WX1803)
--	WX1806 = DFF(WX1805)
--	WX1808 = DFF(WX1807)
--	WX1810 = DFF(WX1809)
--	WX1812 = DFF(WX1811)
--	WX1814 = DFF(WX1813)
--	WX1816 = DFF(WX1815)
--	WX1818 = DFF(WX1817)
--	WX1820 = DFF(WX1819)
--	WX1822 = DFF(WX1821)
--	WX1824 = DFF(WX1823)
--	WX1826 = DFF(WX1825)
--	WX1828 = DFF(WX1827)
--	WX1830 = DFF(WX1829)
--	WX1832 = DFF(WX1831)
--	WX1834 = DFF(WX1833)
--	WX1836 = DFF(WX1835)
--	WX1838 = DFF(WX1837)
--	WX1840 = DFF(WX1839)
--	WX1938 = DFF(WX1937)
--	WX1940 = DFF(WX1939)
--	WX1942 = DFF(WX1941)
--	WX1944 = DFF(WX1943)
--	WX1946 = DFF(WX1945)
--	WX1948 = DFF(WX1947)
--	WX1950 = DFF(WX1949)
--	WX1952 = DFF(WX1951)
--	WX1954 = DFF(WX1953)
--	WX1956 = DFF(WX1955)
--	WX1958 = DFF(WX1957)
--	WX1960 = DFF(WX1959)
--	WX1962 = DFF(WX1961)
--	WX1964 = DFF(WX1963)
--	WX1966 = DFF(WX1965)
--	WX1968 = DFF(WX1967)
--	WX1970 = DFF(WX1969)
--	WX1972 = DFF(WX1971)
--	WX1974 = DFF(WX1973)
--	WX1976 = DFF(WX1975)
--	WX1978 = DFF(WX1977)
--	WX1980 = DFF(WX1979)
--	WX1982 = DFF(WX1981)
--	WX1984 = DFF(WX1983)
--	WX1986 = DFF(WX1985)
--	WX1988 = DFF(WX1987)
--	WX1990 = DFF(WX1989)
--	WX1992 = DFF(WX1991)
--	WX1994 = DFF(WX1993)
--	WX1996 = DFF(WX1995)
--	WX1998 = DFF(WX1997)
--	WX2000 = DFF(WX1999)
--	WX2002 = DFF(WX2001)
--	WX2004 = DFF(WX2003)
--	WX2006 = DFF(WX2005)
--	WX2008 = DFF(WX2007)
--	WX2010 = DFF(WX2009)
--	WX2012 = DFF(WX2011)
--	WX2014 = DFF(WX2013)
--	WX2016 = DFF(WX2015)
--	WX2018 = DFF(WX2017)
--	WX2020 = DFF(WX2019)
--	WX2022 = DFF(WX2021)
--	WX2024 = DFF(WX2023)
--	WX2026 = DFF(WX2025)
--	WX2028 = DFF(WX2027)
--	WX2030 = DFF(WX2029)
--	WX2032 = DFF(WX2031)
--	WX2034 = DFF(WX2033)
--	WX2036 = DFF(WX2035)
--	WX2038 = DFF(WX2037)
--	WX2040 = DFF(WX2039)
--	WX2042 = DFF(WX2041)
--	WX2044 = DFF(WX2043)
--	WX2046 = DFF(WX2045)
--	WX2048 = DFF(WX2047)
--	WX2050 = DFF(WX2049)
--	WX2052 = DFF(WX2051)
--	WX2054 = DFF(WX2053)
--	WX2056 = DFF(WX2055)
--	WX2058 = DFF(WX2057)
--	WX2060 = DFF(WX2059)
--	WX2062 = DFF(WX2061)
--	WX2064 = DFF(WX2063)
--	WX2066 = DFF(WX2065)
--	WX2068 = DFF(WX2067)
--	WX2070 = DFF(WX2069)
--	WX2072 = DFF(WX2071)
--	WX2074 = DFF(WX2073)
--	WX2076 = DFF(WX2075)
--	WX2078 = DFF(WX2077)
--	WX2080 = DFF(WX2079)
--	WX2082 = DFF(WX2081)
--	WX2084 = DFF(WX2083)
--	WX2086 = DFF(WX2085)
--	WX2088 = DFF(WX2087)
--	WX2090 = DFF(WX2089)
--	WX2092 = DFF(WX2091)
--	WX2094 = DFF(WX2093)
--	WX2096 = DFF(WX2095)
--	WX2098 = DFF(WX2097)
--	WX2100 = DFF(WX2099)
--	WX2102 = DFF(WX2101)
--	WX2104 = DFF(WX2103)
--	WX2106 = DFF(WX2105)
--	WX2108 = DFF(WX2107)
--	WX2110 = DFF(WX2109)
--	WX2112 = DFF(WX2111)
--	WX2114 = DFF(WX2113)
--	WX2116 = DFF(WX2115)
--	WX2118 = DFF(WX2117)
--	WX2120 = DFF(WX2119)
--	WX2122 = DFF(WX2121)
--	WX2124 = DFF(WX2123)
--	WX2126 = DFF(WX2125)
--	WX2128 = DFF(WX2127)
--	WX2130 = DFF(WX2129)
--	WX2132 = DFF(WX2131)
--	WX2134 = DFF(WX2133)
--	WX2136 = DFF(WX2135)
--	WX2138 = DFF(WX2137)
--	WX2140 = DFF(WX2139)
--	WX2142 = DFF(WX2141)
--	WX2144 = DFF(WX2143)
--	WX2146 = DFF(WX2145)
--	WX2148 = DFF(WX2147)
--	WX2150 = DFF(WX2149)
--	WX2152 = DFF(WX2151)
--	WX2154 = DFF(WX2153)
--	WX2156 = DFF(WX2155)
--	WX2158 = DFF(WX2157)
--	WX2160 = DFF(WX2159)
--	WX2162 = DFF(WX2161)
--	WX2164 = DFF(WX2163)
--	WX2166 = DFF(WX2165)
--	WX2168 = DFF(WX2167)
--	WX2170 = DFF(WX2169)
--	WX2172 = DFF(WX2171)
--	WX2174 = DFF(WX2173)
--	WX2176 = DFF(WX2175)
--	WX2178 = DFF(WX2177)
--	WX2180 = DFF(WX2179)
--	WX2182 = DFF(WX2181)
--	WX2184 = DFF(WX2183)
--	WX2186 = DFF(WX2185)
--	WX2188 = DFF(WX2187)
--	WX2190 = DFF(WX2189)
--	WX2192 = DFF(WX2191)
--	CRC_OUT_8_0 = DFF(WX2557)
--	CRC_OUT_8_1 = DFF(WX2559)
--	CRC_OUT_8_2 = DFF(WX2561)
--	CRC_OUT_8_3 = DFF(WX2563)
--	CRC_OUT_8_4 = DFF(WX2565)
--	CRC_OUT_8_5 = DFF(WX2567)
--	CRC_OUT_8_6 = DFF(WX2569)
--	CRC_OUT_8_7 = DFF(WX2571)
--	CRC_OUT_8_8 = DFF(WX2573)
--	CRC_OUT_8_9 = DFF(WX2575)
--	CRC_OUT_8_10 = DFF(WX2577)
--	CRC_OUT_8_11 = DFF(WX2579)
--	CRC_OUT_8_12 = DFF(WX2581)
--	CRC_OUT_8_13 = DFF(WX2583)
--	CRC_OUT_8_14 = DFF(WX2585)
--	CRC_OUT_8_15 = DFF(WX2587)
--	CRC_OUT_8_16 = DFF(WX2589)
--	CRC_OUT_8_17 = DFF(WX2591)
--	CRC_OUT_8_18 = DFF(WX2593)
--	CRC_OUT_8_19 = DFF(WX2595)
--	CRC_OUT_8_20 = DFF(WX2597)
--	CRC_OUT_8_21 = DFF(WX2599)
--	CRC_OUT_8_22 = DFF(WX2601)
--	CRC_OUT_8_23 = DFF(WX2603)
--	CRC_OUT_8_24 = DFF(WX2605)
--	CRC_OUT_8_25 = DFF(WX2607)
--	CRC_OUT_8_26 = DFF(WX2609)
--	CRC_OUT_8_27 = DFF(WX2611)
--	CRC_OUT_8_28 = DFF(WX2613)
--	CRC_OUT_8_29 = DFF(WX2615)
--	CRC_OUT_8_30 = DFF(WX2617)
--	CRC_OUT_8_31 = DFF(WX2619)
--	WX3071 = DFF(WX3070)
--	WX3073 = DFF(WX3072)
--	WX3075 = DFF(WX3074)
--	WX3077 = DFF(WX3076)
--	WX3079 = DFF(WX3078)
--	WX3081 = DFF(WX3080)
--	WX3083 = DFF(WX3082)
--	WX3085 = DFF(WX3084)
--	WX3087 = DFF(WX3086)
--	WX3089 = DFF(WX3088)
--	WX3091 = DFF(WX3090)
--	WX3093 = DFF(WX3092)
--	WX3095 = DFF(WX3094)
--	WX3097 = DFF(WX3096)
--	WX3099 = DFF(WX3098)
--	WX3101 = DFF(WX3100)
--	WX3103 = DFF(WX3102)
--	WX3105 = DFF(WX3104)
--	WX3107 = DFF(WX3106)
--	WX3109 = DFF(WX3108)
--	WX3111 = DFF(WX3110)
--	WX3113 = DFF(WX3112)
--	WX3115 = DFF(WX3114)
--	WX3117 = DFF(WX3116)
--	WX3119 = DFF(WX3118)
--	WX3121 = DFF(WX3120)
--	WX3123 = DFF(WX3122)
--	WX3125 = DFF(WX3124)
--	WX3127 = DFF(WX3126)
--	WX3129 = DFF(WX3128)
--	WX3131 = DFF(WX3130)
--	WX3133 = DFF(WX3132)
--	WX3231 = DFF(WX3230)
--	WX3233 = DFF(WX3232)
--	WX3235 = DFF(WX3234)
--	WX3237 = DFF(WX3236)
--	WX3239 = DFF(WX3238)
--	WX3241 = DFF(WX3240)
--	WX3243 = DFF(WX3242)
--	WX3245 = DFF(WX3244)
--	WX3247 = DFF(WX3246)
--	WX3249 = DFF(WX3248)
--	WX3251 = DFF(WX3250)
--	WX3253 = DFF(WX3252)
--	WX3255 = DFF(WX3254)
--	WX3257 = DFF(WX3256)
--	WX3259 = DFF(WX3258)
--	WX3261 = DFF(WX3260)
--	WX3263 = DFF(WX3262)
--	WX3265 = DFF(WX3264)
--	WX3267 = DFF(WX3266)
--	WX3269 = DFF(WX3268)
--	WX3271 = DFF(WX3270)
--	WX3273 = DFF(WX3272)
--	WX3275 = DFF(WX3274)
--	WX3277 = DFF(WX3276)
--	WX3279 = DFF(WX3278)
--	WX3281 = DFF(WX3280)
--	WX3283 = DFF(WX3282)
--	WX3285 = DFF(WX3284)
--	WX3287 = DFF(WX3286)
--	WX3289 = DFF(WX3288)
--	WX3291 = DFF(WX3290)
--	WX3293 = DFF(WX3292)
--	WX3295 = DFF(WX3294)
--	WX3297 = DFF(WX3296)
--	WX3299 = DFF(WX3298)
--	WX3301 = DFF(WX3300)
--	WX3303 = DFF(WX3302)
--	WX3305 = DFF(WX3304)
--	WX3307 = DFF(WX3306)
--	WX3309 = DFF(WX3308)
--	WX3311 = DFF(WX3310)
--	WX3313 = DFF(WX3312)
--	WX3315 = DFF(WX3314)
--	WX3317 = DFF(WX3316)
--	WX3319 = DFF(WX3318)
--	WX3321 = DFF(WX3320)
--	WX3323 = DFF(WX3322)
--	WX3325 = DFF(WX3324)
--	WX3327 = DFF(WX3326)
--	WX3329 = DFF(WX3328)
--	WX3331 = DFF(WX3330)
--	WX3333 = DFF(WX3332)
--	WX3335 = DFF(WX3334)
--	WX3337 = DFF(WX3336)
--	WX3339 = DFF(WX3338)
--	WX3341 = DFF(WX3340)
--	WX3343 = DFF(WX3342)
--	WX3345 = DFF(WX3344)
--	WX3347 = DFF(WX3346)
--	WX3349 = DFF(WX3348)
--	WX3351 = DFF(WX3350)
--	WX3353 = DFF(WX3352)
--	WX3355 = DFF(WX3354)
--	WX3357 = DFF(WX3356)
--	WX3359 = DFF(WX3358)
--	WX3361 = DFF(WX3360)
--	WX3363 = DFF(WX3362)
--	WX3365 = DFF(WX3364)
--	WX3367 = DFF(WX3366)
--	WX3369 = DFF(WX3368)
--	WX3371 = DFF(WX3370)
--	WX3373 = DFF(WX3372)
--	WX3375 = DFF(WX3374)
--	WX3377 = DFF(WX3376)
--	WX3379 = DFF(WX3378)
--	WX3381 = DFF(WX3380)
--	WX3383 = DFF(WX3382)
--	WX3385 = DFF(WX3384)
--	WX3387 = DFF(WX3386)
--	WX3389 = DFF(WX3388)
--	WX3391 = DFF(WX3390)
--	WX3393 = DFF(WX3392)
--	WX3395 = DFF(WX3394)
--	WX3397 = DFF(WX3396)
--	WX3399 = DFF(WX3398)
--	WX3401 = DFF(WX3400)
--	WX3403 = DFF(WX3402)
--	WX3405 = DFF(WX3404)
--	WX3407 = DFF(WX3406)
--	WX3409 = DFF(WX3408)
--	WX3411 = DFF(WX3410)
--	WX3413 = DFF(WX3412)
--	WX3415 = DFF(WX3414)
--	WX3417 = DFF(WX3416)
--	WX3419 = DFF(WX3418)
--	WX3421 = DFF(WX3420)
--	WX3423 = DFF(WX3422)
--	WX3425 = DFF(WX3424)
--	WX3427 = DFF(WX3426)
--	WX3429 = DFF(WX3428)
--	WX3431 = DFF(WX3430)
--	WX3433 = DFF(WX3432)
--	WX3435 = DFF(WX3434)
--	WX3437 = DFF(WX3436)
--	WX3439 = DFF(WX3438)
--	WX3441 = DFF(WX3440)
--	WX3443 = DFF(WX3442)
--	WX3445 = DFF(WX3444)
--	WX3447 = DFF(WX3446)
--	WX3449 = DFF(WX3448)
--	WX3451 = DFF(WX3450)
--	WX3453 = DFF(WX3452)
--	WX3455 = DFF(WX3454)
--	WX3457 = DFF(WX3456)
--	WX3459 = DFF(WX3458)
--	WX3461 = DFF(WX3460)
--	WX3463 = DFF(WX3462)
--	WX3465 = DFF(WX3464)
--	WX3467 = DFF(WX3466)
--	WX3469 = DFF(WX3468)
--	WX3471 = DFF(WX3470)
--	WX3473 = DFF(WX3472)
--	WX3475 = DFF(WX3474)
--	WX3477 = DFF(WX3476)
--	WX3479 = DFF(WX3478)
--	WX3481 = DFF(WX3480)
--	WX3483 = DFF(WX3482)
--	WX3485 = DFF(WX3484)
--	CRC_OUT_7_0 = DFF(WX3850)
--	CRC_OUT_7_1 = DFF(WX3852)
--	CRC_OUT_7_2 = DFF(WX3854)
--	CRC_OUT_7_3 = DFF(WX3856)
--	CRC_OUT_7_4 = DFF(WX3858)
--	CRC_OUT_7_5 = DFF(WX3860)
--	CRC_OUT_7_6 = DFF(WX3862)
--	CRC_OUT_7_7 = DFF(WX3864)
--	CRC_OUT_7_8 = DFF(WX3866)
--	CRC_OUT_7_9 = DFF(WX3868)
--	CRC_OUT_7_10 = DFF(WX3870)
--	CRC_OUT_7_11 = DFF(WX3872)
--	CRC_OUT_7_12 = DFF(WX3874)
--	CRC_OUT_7_13 = DFF(WX3876)
--	CRC_OUT_7_14 = DFF(WX3878)
--	CRC_OUT_7_15 = DFF(WX3880)
--	CRC_OUT_7_16 = DFF(WX3882)
--	CRC_OUT_7_17 = DFF(WX3884)
--	CRC_OUT_7_18 = DFF(WX3886)
--	CRC_OUT_7_19 = DFF(WX3888)
--	CRC_OUT_7_20 = DFF(WX3890)
--	CRC_OUT_7_21 = DFF(WX3892)
--	CRC_OUT_7_22 = DFF(WX3894)
--	CRC_OUT_7_23 = DFF(WX3896)
--	CRC_OUT_7_24 = DFF(WX3898)
--	CRC_OUT_7_25 = DFF(WX3900)
--	CRC_OUT_7_26 = DFF(WX3902)
--	CRC_OUT_7_27 = DFF(WX3904)
--	CRC_OUT_7_28 = DFF(WX3906)
--	CRC_OUT_7_29 = DFF(WX3908)
--	CRC_OUT_7_30 = DFF(WX3910)
--	CRC_OUT_7_31 = DFF(WX3912)
--	WX4364 = DFF(WX4363)
--	WX4366 = DFF(WX4365)
--	WX4368 = DFF(WX4367)
--	WX4370 = DFF(WX4369)
--	WX4372 = DFF(WX4371)
--	WX4374 = DFF(WX4373)
--	WX4376 = DFF(WX4375)
--	WX4378 = DFF(WX4377)
--	WX4380 = DFF(WX4379)
--	WX4382 = DFF(WX4381)
--	WX4384 = DFF(WX4383)
--	WX4386 = DFF(WX4385)
--	WX4388 = DFF(WX4387)
--	WX4390 = DFF(WX4389)
--	WX4392 = DFF(WX4391)
--	WX4394 = DFF(WX4393)
--	WX4396 = DFF(WX4395)
--	WX4398 = DFF(WX4397)
--	WX4400 = DFF(WX4399)
--	WX4402 = DFF(WX4401)
--	WX4404 = DFF(WX4403)
--	WX4406 = DFF(WX4405)
--	WX4408 = DFF(WX4407)
--	WX4410 = DFF(WX4409)
--	WX4412 = DFF(WX4411)
--	WX4414 = DFF(WX4413)
--	WX4416 = DFF(WX4415)
--	WX4418 = DFF(WX4417)
--	WX4420 = DFF(WX4419)
--	WX4422 = DFF(WX4421)
--	WX4424 = DFF(WX4423)
--	WX4426 = DFF(WX4425)
--	WX4524 = DFF(WX4523)
--	WX4526 = DFF(WX4525)
--	WX4528 = DFF(WX4527)
--	WX4530 = DFF(WX4529)
--	WX4532 = DFF(WX4531)
--	WX4534 = DFF(WX4533)
--	WX4536 = DFF(WX4535)
--	WX4538 = DFF(WX4537)
--	WX4540 = DFF(WX4539)
--	WX4542 = DFF(WX4541)
--	WX4544 = DFF(WX4543)
--	WX4546 = DFF(WX4545)
--	WX4548 = DFF(WX4547)
--	WX4550 = DFF(WX4549)
--	WX4552 = DFF(WX4551)
--	WX4554 = DFF(WX4553)
--	WX4556 = DFF(WX4555)
--	WX4558 = DFF(WX4557)
--	WX4560 = DFF(WX4559)
--	WX4562 = DFF(WX4561)
--	WX4564 = DFF(WX4563)
--	WX4566 = DFF(WX4565)
--	WX4568 = DFF(WX4567)
--	WX4570 = DFF(WX4569)
--	WX4572 = DFF(WX4571)
--	WX4574 = DFF(WX4573)
--	WX4576 = DFF(WX4575)
--	WX4578 = DFF(WX4577)
--	WX4580 = DFF(WX4579)
--	WX4582 = DFF(WX4581)
--	WX4584 = DFF(WX4583)
--	WX4586 = DFF(WX4585)
--	WX4588 = DFF(WX4587)
--	WX4590 = DFF(WX4589)
--	WX4592 = DFF(WX4591)
--	WX4594 = DFF(WX4593)
--	WX4596 = DFF(WX4595)
--	WX4598 = DFF(WX4597)
--	WX4600 = DFF(WX4599)
--	WX4602 = DFF(WX4601)
--	WX4604 = DFF(WX4603)
--	WX4606 = DFF(WX4605)
--	WX4608 = DFF(WX4607)
--	WX4610 = DFF(WX4609)
--	WX4612 = DFF(WX4611)
--	WX4614 = DFF(WX4613)
--	WX4616 = DFF(WX4615)
--	WX4618 = DFF(WX4617)
--	WX4620 = DFF(WX4619)
--	WX4622 = DFF(WX4621)
--	WX4624 = DFF(WX4623)
--	WX4626 = DFF(WX4625)
--	WX4628 = DFF(WX4627)
--	WX4630 = DFF(WX4629)
--	WX4632 = DFF(WX4631)
--	WX4634 = DFF(WX4633)
--	WX4636 = DFF(WX4635)
--	WX4638 = DFF(WX4637)
--	WX4640 = DFF(WX4639)
--	WX4642 = DFF(WX4641)
--	WX4644 = DFF(WX4643)
--	WX4646 = DFF(WX4645)
--	WX4648 = DFF(WX4647)
--	WX4650 = DFF(WX4649)
--	WX4652 = DFF(WX4651)
--	WX4654 = DFF(WX4653)
--	WX4656 = DFF(WX4655)
--	WX4658 = DFF(WX4657)
--	WX4660 = DFF(WX4659)
--	WX4662 = DFF(WX4661)
--	WX4664 = DFF(WX4663)
--	WX4666 = DFF(WX4665)
--	WX4668 = DFF(WX4667)
--	WX4670 = DFF(WX4669)
--	WX4672 = DFF(WX4671)
--	WX4674 = DFF(WX4673)
--	WX4676 = DFF(WX4675)
--	WX4678 = DFF(WX4677)
--	WX4680 = DFF(WX4679)
--	WX4682 = DFF(WX4681)
--	WX4684 = DFF(WX4683)
--	WX4686 = DFF(WX4685)
--	WX4688 = DFF(WX4687)
--	WX4690 = DFF(WX4689)
--	WX4692 = DFF(WX4691)
--	WX4694 = DFF(WX4693)
--	WX4696 = DFF(WX4695)
--	WX4698 = DFF(WX4697)
--	WX4700 = DFF(WX4699)
--	WX4702 = DFF(WX4701)
--	WX4704 = DFF(WX4703)
--	WX4706 = DFF(WX4705)
--	WX4708 = DFF(WX4707)
--	WX4710 = DFF(WX4709)
--	WX4712 = DFF(WX4711)
--	WX4714 = DFF(WX4713)
--	WX4716 = DFF(WX4715)
--	WX4718 = DFF(WX4717)
--	WX4720 = DFF(WX4719)
--	WX4722 = DFF(WX4721)
--	WX4724 = DFF(WX4723)
--	WX4726 = DFF(WX4725)
--	WX4728 = DFF(WX4727)
--	WX4730 = DFF(WX4729)
--	WX4732 = DFF(WX4731)
--	WX4734 = DFF(WX4733)
--	WX4736 = DFF(WX4735)
--	WX4738 = DFF(WX4737)
--	WX4740 = DFF(WX4739)
--	WX4742 = DFF(WX4741)
--	WX4744 = DFF(WX4743)
--	WX4746 = DFF(WX4745)
--	WX4748 = DFF(WX4747)
--	WX4750 = DFF(WX4749)
--	WX4752 = DFF(WX4751)
--	WX4754 = DFF(WX4753)
--	WX4756 = DFF(WX4755)
--	WX4758 = DFF(WX4757)
--	WX4760 = DFF(WX4759)
--	WX4762 = DFF(WX4761)
--	WX4764 = DFF(WX4763)
--	WX4766 = DFF(WX4765)
--	WX4768 = DFF(WX4767)
--	WX4770 = DFF(WX4769)
--	WX4772 = DFF(WX4771)
--	WX4774 = DFF(WX4773)
--	WX4776 = DFF(WX4775)
--	WX4778 = DFF(WX4777)
--	CRC_OUT_6_0 = DFF(WX5143)
--	CRC_OUT_6_1 = DFF(WX5145)
--	CRC_OUT_6_2 = DFF(WX5147)
--	CRC_OUT_6_3 = DFF(WX5149)
--	CRC_OUT_6_4 = DFF(WX5151)
--	CRC_OUT_6_5 = DFF(WX5153)
--	CRC_OUT_6_6 = DFF(WX5155)
--	CRC_OUT_6_7 = DFF(WX5157)
--	CRC_OUT_6_8 = DFF(WX5159)
--	CRC_OUT_6_9 = DFF(WX5161)
--	CRC_OUT_6_10 = DFF(WX5163)
--	CRC_OUT_6_11 = DFF(WX5165)
--	CRC_OUT_6_12 = DFF(WX5167)
--	CRC_OUT_6_13 = DFF(WX5169)
--	CRC_OUT_6_14 = DFF(WX5171)
--	CRC_OUT_6_15 = DFF(WX5173)
--	CRC_OUT_6_16 = DFF(WX5175)
--	CRC_OUT_6_17 = DFF(WX5177)
--	CRC_OUT_6_18 = DFF(WX5179)
--	CRC_OUT_6_19 = DFF(WX5181)
--	CRC_OUT_6_20 = DFF(WX5183)
--	CRC_OUT_6_21 = DFF(WX5185)
--	CRC_OUT_6_22 = DFF(WX5187)
--	CRC_OUT_6_23 = DFF(WX5189)
--	CRC_OUT_6_24 = DFF(WX5191)
--	CRC_OUT_6_25 = DFF(WX5193)
--	CRC_OUT_6_26 = DFF(WX5195)
--	CRC_OUT_6_27 = DFF(WX5197)
--	CRC_OUT_6_28 = DFF(WX5199)
--	CRC_OUT_6_29 = DFF(WX5201)
--	CRC_OUT_6_30 = DFF(WX5203)
--	CRC_OUT_6_31 = DFF(WX5205)
--	WX5657 = DFF(WX5656)
--	WX5659 = DFF(WX5658)
--	WX5661 = DFF(WX5660)
--	WX5663 = DFF(WX5662)
--	WX5665 = DFF(WX5664)
--	WX5667 = DFF(WX5666)
--	WX5669 = DFF(WX5668)
--	WX5671 = DFF(WX5670)
--	WX5673 = DFF(WX5672)
--	WX5675 = DFF(WX5674)
--	WX5677 = DFF(WX5676)
--	WX5679 = DFF(WX5678)
--	WX5681 = DFF(WX5680)
--	WX5683 = DFF(WX5682)
--	WX5685 = DFF(WX5684)
--	WX5687 = DFF(WX5686)
--	WX5689 = DFF(WX5688)
--	WX5691 = DFF(WX5690)
--	WX5693 = DFF(WX5692)
--	WX5695 = DFF(WX5694)
--	WX5697 = DFF(WX5696)
--	WX5699 = DFF(WX5698)
--	WX5701 = DFF(WX5700)
--	WX5703 = DFF(WX5702)
--	WX5705 = DFF(WX5704)
--	WX5707 = DFF(WX5706)
--	WX5709 = DFF(WX5708)
--	WX5711 = DFF(WX5710)
--	WX5713 = DFF(WX5712)
--	WX5715 = DFF(WX5714)
--	WX5717 = DFF(WX5716)
--	WX5719 = DFF(WX5718)
--	WX5817 = DFF(WX5816)
--	WX5819 = DFF(WX5818)
--	WX5821 = DFF(WX5820)
--	WX5823 = DFF(WX5822)
--	WX5825 = DFF(WX5824)
--	WX5827 = DFF(WX5826)
--	WX5829 = DFF(WX5828)
--	WX5831 = DFF(WX5830)
--	WX5833 = DFF(WX5832)
--	WX5835 = DFF(WX5834)
--	WX5837 = DFF(WX5836)
--	WX5839 = DFF(WX5838)
--	WX5841 = DFF(WX5840)
--	WX5843 = DFF(WX5842)
--	WX5845 = DFF(WX5844)
--	WX5847 = DFF(WX5846)
--	WX5849 = DFF(WX5848)
--	WX5851 = DFF(WX5850)
--	WX5853 = DFF(WX5852)
--	WX5855 = DFF(WX5854)
--	WX5857 = DFF(WX5856)
--	WX5859 = DFF(WX5858)
--	WX5861 = DFF(WX5860)
--	WX5863 = DFF(WX5862)
--	WX5865 = DFF(WX5864)
--	WX5867 = DFF(WX5866)
--	WX5869 = DFF(WX5868)
--	WX5871 = DFF(WX5870)
--	WX5873 = DFF(WX5872)
--	WX5875 = DFF(WX5874)
--	WX5877 = DFF(WX5876)
--	WX5879 = DFF(WX5878)
--	WX5881 = DFF(WX5880)
--	WX5883 = DFF(WX5882)
--	WX5885 = DFF(WX5884)
--	WX5887 = DFF(WX5886)
--	WX5889 = DFF(WX5888)
--	WX5891 = DFF(WX5890)
--	WX5893 = DFF(WX5892)
--	WX5895 = DFF(WX5894)
--	WX5897 = DFF(WX5896)
--	WX5899 = DFF(WX5898)
--	WX5901 = DFF(WX5900)
--	WX5903 = DFF(WX5902)
--	WX5905 = DFF(WX5904)
--	WX5907 = DFF(WX5906)
--	WX5909 = DFF(WX5908)
--	WX5911 = DFF(WX5910)
--	WX5913 = DFF(WX5912)
--	WX5915 = DFF(WX5914)
--	WX5917 = DFF(WX5916)
--	WX5919 = DFF(WX5918)
--	WX5921 = DFF(WX5920)
--	WX5923 = DFF(WX5922)
--	WX5925 = DFF(WX5924)
--	WX5927 = DFF(WX5926)
--	WX5929 = DFF(WX5928)
--	WX5931 = DFF(WX5930)
--	WX5933 = DFF(WX5932)
--	WX5935 = DFF(WX5934)
--	WX5937 = DFF(WX5936)
--	WX5939 = DFF(WX5938)
--	WX5941 = DFF(WX5940)
--	WX5943 = DFF(WX5942)
--	WX5945 = DFF(WX5944)
--	WX5947 = DFF(WX5946)
--	WX5949 = DFF(WX5948)
--	WX5951 = DFF(WX5950)
--	WX5953 = DFF(WX5952)
--	WX5955 = DFF(WX5954)
--	WX5957 = DFF(WX5956)
--	WX5959 = DFF(WX5958)
--	WX5961 = DFF(WX5960)
--	WX5963 = DFF(WX5962)
--	WX5965 = DFF(WX5964)
--	WX5967 = DFF(WX5966)
--	WX5969 = DFF(WX5968)
--	WX5971 = DFF(WX5970)
--	WX5973 = DFF(WX5972)
--	WX5975 = DFF(WX5974)
--	WX5977 = DFF(WX5976)
--	WX5979 = DFF(WX5978)
--	WX5981 = DFF(WX5980)
--	WX5983 = DFF(WX5982)
--	WX5985 = DFF(WX5984)
--	WX5987 = DFF(WX5986)
--	WX5989 = DFF(WX5988)
--	WX5991 = DFF(WX5990)
--	WX5993 = DFF(WX5992)
--	WX5995 = DFF(WX5994)
--	WX5997 = DFF(WX5996)
--	WX5999 = DFF(WX5998)
--	WX6001 = DFF(WX6000)
--	WX6003 = DFF(WX6002)
--	WX6005 = DFF(WX6004)
--	WX6007 = DFF(WX6006)
--	WX6009 = DFF(WX6008)
--	WX6011 = DFF(WX6010)
--	WX6013 = DFF(WX6012)
--	WX6015 = DFF(WX6014)
--	WX6017 = DFF(WX6016)
--	WX6019 = DFF(WX6018)
--	WX6021 = DFF(WX6020)
--	WX6023 = DFF(WX6022)
--	WX6025 = DFF(WX6024)
--	WX6027 = DFF(WX6026)
--	WX6029 = DFF(WX6028)
--	WX6031 = DFF(WX6030)
--	WX6033 = DFF(WX6032)
--	WX6035 = DFF(WX6034)
--	WX6037 = DFF(WX6036)
--	WX6039 = DFF(WX6038)
--	WX6041 = DFF(WX6040)
--	WX6043 = DFF(WX6042)
--	WX6045 = DFF(WX6044)
--	WX6047 = DFF(WX6046)
--	WX6049 = DFF(WX6048)
--	WX6051 = DFF(WX6050)
--	WX6053 = DFF(WX6052)
--	WX6055 = DFF(WX6054)
--	WX6057 = DFF(WX6056)
--	WX6059 = DFF(WX6058)
--	WX6061 = DFF(WX6060)
--	WX6063 = DFF(WX6062)
--	WX6065 = DFF(WX6064)
--	WX6067 = DFF(WX6066)
--	WX6069 = DFF(WX6068)
--	WX6071 = DFF(WX6070)
--	CRC_OUT_5_0 = DFF(WX6436)
--	CRC_OUT_5_1 = DFF(WX6438)
--	CRC_OUT_5_2 = DFF(WX6440)
--	CRC_OUT_5_3 = DFF(WX6442)
--	CRC_OUT_5_4 = DFF(WX6444)
--	CRC_OUT_5_5 = DFF(WX6446)
--	CRC_OUT_5_6 = DFF(WX6448)
--	CRC_OUT_5_7 = DFF(WX6450)
--	CRC_OUT_5_8 = DFF(WX6452)
--	CRC_OUT_5_9 = DFF(WX6454)
--	CRC_OUT_5_10 = DFF(WX6456)
--	CRC_OUT_5_11 = DFF(WX6458)
--	CRC_OUT_5_12 = DFF(WX6460)
--	CRC_OUT_5_13 = DFF(WX6462)
--	CRC_OUT_5_14 = DFF(WX6464)
--	CRC_OUT_5_15 = DFF(WX6466)
--	CRC_OUT_5_16 = DFF(WX6468)
--	CRC_OUT_5_17 = DFF(WX6470)
--	CRC_OUT_5_18 = DFF(WX6472)
--	CRC_OUT_5_19 = DFF(WX6474)
--	CRC_OUT_5_20 = DFF(WX6476)
--	CRC_OUT_5_21 = DFF(WX6478)
--	CRC_OUT_5_22 = DFF(WX6480)
--	CRC_OUT_5_23 = DFF(WX6482)
--	CRC_OUT_5_24 = DFF(WX6484)
--	CRC_OUT_5_25 = DFF(WX6486)
--	CRC_OUT_5_26 = DFF(WX6488)
--	CRC_OUT_5_27 = DFF(WX6490)
--	CRC_OUT_5_28 = DFF(WX6492)
--	CRC_OUT_5_29 = DFF(WX6494)
--	CRC_OUT_5_30 = DFF(WX6496)
--	CRC_OUT_5_31 = DFF(WX6498)
--	WX6950 = DFF(WX6949)
--	WX6952 = DFF(WX6951)
--	WX6954 = DFF(WX6953)
--	WX6956 = DFF(WX6955)
--	WX6958 = DFF(WX6957)
--	WX6960 = DFF(WX6959)
--	WX6962 = DFF(WX6961)
--	WX6964 = DFF(WX6963)
--	WX6966 = DFF(WX6965)
--	WX6968 = DFF(WX6967)
--	WX6970 = DFF(WX6969)
--	WX6972 = DFF(WX6971)
--	WX6974 = DFF(WX6973)
--	WX6976 = DFF(WX6975)
--	WX6978 = DFF(WX6977)
--	WX6980 = DFF(WX6979)
--	WX6982 = DFF(WX6981)
--	WX6984 = DFF(WX6983)
--	WX6986 = DFF(WX6985)
--	WX6988 = DFF(WX6987)
--	WX6990 = DFF(WX6989)
--	WX6992 = DFF(WX6991)
--	WX6994 = DFF(WX6993)
--	WX6996 = DFF(WX6995)
--	WX6998 = DFF(WX6997)
--	WX7000 = DFF(WX6999)
--	WX7002 = DFF(WX7001)
--	WX7004 = DFF(WX7003)
--	WX7006 = DFF(WX7005)
--	WX7008 = DFF(WX7007)
--	WX7010 = DFF(WX7009)
--	WX7012 = DFF(WX7011)
--	WX7110 = DFF(WX7109)
--	WX7112 = DFF(WX7111)
--	WX7114 = DFF(WX7113)
--	WX7116 = DFF(WX7115)
--	WX7118 = DFF(WX7117)
--	WX7120 = DFF(WX7119)
--	WX7122 = DFF(WX7121)
--	WX7124 = DFF(WX7123)
--	WX7126 = DFF(WX7125)
--	WX7128 = DFF(WX7127)
--	WX7130 = DFF(WX7129)
--	WX7132 = DFF(WX7131)
--	WX7134 = DFF(WX7133)
--	WX7136 = DFF(WX7135)
--	WX7138 = DFF(WX7137)
--	WX7140 = DFF(WX7139)
--	WX7142 = DFF(WX7141)
--	WX7144 = DFF(WX7143)
--	WX7146 = DFF(WX7145)
--	WX7148 = DFF(WX7147)
--	WX7150 = DFF(WX7149)
--	WX7152 = DFF(WX7151)
--	WX7154 = DFF(WX7153)
--	WX7156 = DFF(WX7155)
--	WX7158 = DFF(WX7157)
--	WX7160 = DFF(WX7159)
--	WX7162 = DFF(WX7161)
--	WX7164 = DFF(WX7163)
--	WX7166 = DFF(WX7165)
--	WX7168 = DFF(WX7167)
--	WX7170 = DFF(WX7169)
--	WX7172 = DFF(WX7171)
--	WX7174 = DFF(WX7173)
--	WX7176 = DFF(WX7175)
--	WX7178 = DFF(WX7177)
--	WX7180 = DFF(WX7179)
--	WX7182 = DFF(WX7181)
--	WX7184 = DFF(WX7183)
--	WX7186 = DFF(WX7185)
--	WX7188 = DFF(WX7187)
--	WX7190 = DFF(WX7189)
--	WX7192 = DFF(WX7191)
--	WX7194 = DFF(WX7193)
--	WX7196 = DFF(WX7195)
--	WX7198 = DFF(WX7197)
--	WX7200 = DFF(WX7199)
--	WX7202 = DFF(WX7201)
--	WX7204 = DFF(WX7203)
--	WX7206 = DFF(WX7205)
--	WX7208 = DFF(WX7207)
--	WX7210 = DFF(WX7209)
--	WX7212 = DFF(WX7211)
--	WX7214 = DFF(WX7213)
--	WX7216 = DFF(WX7215)
--	WX7218 = DFF(WX7217)
--	WX7220 = DFF(WX7219)
--	WX7222 = DFF(WX7221)
--	WX7224 = DFF(WX7223)
--	WX7226 = DFF(WX7225)
--	WX7228 = DFF(WX7227)
--	WX7230 = DFF(WX7229)
--	WX7232 = DFF(WX7231)
--	WX7234 = DFF(WX7233)
--	WX7236 = DFF(WX7235)
--	WX7238 = DFF(WX7237)
--	WX7240 = DFF(WX7239)
--	WX7242 = DFF(WX7241)
--	WX7244 = DFF(WX7243)
--	WX7246 = DFF(WX7245)
--	WX7248 = DFF(WX7247)
--	WX7250 = DFF(WX7249)
--	WX7252 = DFF(WX7251)
--	WX7254 = DFF(WX7253)
--	WX7256 = DFF(WX7255)
--	WX7258 = DFF(WX7257)
--	WX7260 = DFF(WX7259)
--	WX7262 = DFF(WX7261)
--	WX7264 = DFF(WX7263)
--	WX7266 = DFF(WX7265)
--	WX7268 = DFF(WX7267)
--	WX7270 = DFF(WX7269)
--	WX7272 = DFF(WX7271)
--	WX7274 = DFF(WX7273)
--	WX7276 = DFF(WX7275)
--	WX7278 = DFF(WX7277)
--	WX7280 = DFF(WX7279)
--	WX7282 = DFF(WX7281)
--	WX7284 = DFF(WX7283)
--	WX7286 = DFF(WX7285)
--	WX7288 = DFF(WX7287)
--	WX7290 = DFF(WX7289)
--	WX7292 = DFF(WX7291)
--	WX7294 = DFF(WX7293)
--	WX7296 = DFF(WX7295)
--	WX7298 = DFF(WX7297)
--	WX7300 = DFF(WX7299)
--	WX7302 = DFF(WX7301)
--	WX7304 = DFF(WX7303)
--	WX7306 = DFF(WX7305)
--	WX7308 = DFF(WX7307)
--	WX7310 = DFF(WX7309)
--	WX7312 = DFF(WX7311)
--	WX7314 = DFF(WX7313)
--	WX7316 = DFF(WX7315)
--	WX7318 = DFF(WX7317)
--	WX7320 = DFF(WX7319)
--	WX7322 = DFF(WX7321)
--	WX7324 = DFF(WX7323)
--	WX7326 = DFF(WX7325)
--	WX7328 = DFF(WX7327)
--	WX7330 = DFF(WX7329)
--	WX7332 = DFF(WX7331)
--	WX7334 = DFF(WX7333)
--	WX7336 = DFF(WX7335)
--	WX7338 = DFF(WX7337)
--	WX7340 = DFF(WX7339)
--	WX7342 = DFF(WX7341)
--	WX7344 = DFF(WX7343)
--	WX7346 = DFF(WX7345)
--	WX7348 = DFF(WX7347)
--	WX7350 = DFF(WX7349)
--	WX7352 = DFF(WX7351)
--	WX7354 = DFF(WX7353)
--	WX7356 = DFF(WX7355)
--	WX7358 = DFF(WX7357)
--	WX7360 = DFF(WX7359)
--	WX7362 = DFF(WX7361)
--	WX7364 = DFF(WX7363)
--	CRC_OUT_4_0 = DFF(WX7729)
--	CRC_OUT_4_1 = DFF(WX7731)
--	CRC_OUT_4_2 = DFF(WX7733)
--	CRC_OUT_4_3 = DFF(WX7735)
--	CRC_OUT_4_4 = DFF(WX7737)
--	CRC_OUT_4_5 = DFF(WX7739)
--	CRC_OUT_4_6 = DFF(WX7741)
--	CRC_OUT_4_7 = DFF(WX7743)
--	CRC_OUT_4_8 = DFF(WX7745)
--	CRC_OUT_4_9 = DFF(WX7747)
--	CRC_OUT_4_10 = DFF(WX7749)
--	CRC_OUT_4_11 = DFF(WX7751)
--	CRC_OUT_4_12 = DFF(WX7753)
--	CRC_OUT_4_13 = DFF(WX7755)
--	CRC_OUT_4_14 = DFF(WX7757)
--	CRC_OUT_4_15 = DFF(WX7759)
--	CRC_OUT_4_16 = DFF(WX7761)
--	CRC_OUT_4_17 = DFF(WX7763)
--	CRC_OUT_4_18 = DFF(WX7765)
--	CRC_OUT_4_19 = DFF(WX7767)
--	CRC_OUT_4_20 = DFF(WX7769)
--	CRC_OUT_4_21 = DFF(WX7771)
--	CRC_OUT_4_22 = DFF(WX7773)
--	CRC_OUT_4_23 = DFF(WX7775)
--	CRC_OUT_4_24 = DFF(WX7777)
--	CRC_OUT_4_25 = DFF(WX7779)
--	CRC_OUT_4_26 = DFF(WX7781)
--	CRC_OUT_4_27 = DFF(WX7783)
--	CRC_OUT_4_28 = DFF(WX7785)
--	CRC_OUT_4_29 = DFF(WX7787)
--	CRC_OUT_4_30 = DFF(WX7789)
--	CRC_OUT_4_31 = DFF(WX7791)
--	WX8243 = DFF(WX8242)
--	WX8245 = DFF(WX8244)
--	WX8247 = DFF(WX8246)
--	WX8249 = DFF(WX8248)
--	WX8251 = DFF(WX8250)
--	WX8253 = DFF(WX8252)
--	WX8255 = DFF(WX8254)
--	WX8257 = DFF(WX8256)
--	WX8259 = DFF(WX8258)
--	WX8261 = DFF(WX8260)
--	WX8263 = DFF(WX8262)
--	WX8265 = DFF(WX8264)
--	WX8267 = DFF(WX8266)
--	WX8269 = DFF(WX8268)
--	WX8271 = DFF(WX8270)
--	WX8273 = DFF(WX8272)
--	WX8275 = DFF(WX8274)
--	WX8277 = DFF(WX8276)
--	WX8279 = DFF(WX8278)
--	WX8281 = DFF(WX8280)
--	WX8283 = DFF(WX8282)
--	WX8285 = DFF(WX8284)
--	WX8287 = DFF(WX8286)
--	WX8289 = DFF(WX8288)
--	WX8291 = DFF(WX8290)
--	WX8293 = DFF(WX8292)
--	WX8295 = DFF(WX8294)
--	WX8297 = DFF(WX8296)
--	WX8299 = DFF(WX8298)
--	WX8301 = DFF(WX8300)
--	WX8303 = DFF(WX8302)
--	WX8305 = DFF(WX8304)
--	WX8403 = DFF(WX8402)
--	WX8405 = DFF(WX8404)
--	WX8407 = DFF(WX8406)
--	WX8409 = DFF(WX8408)
--	WX8411 = DFF(WX8410)
--	WX8413 = DFF(WX8412)
--	WX8415 = DFF(WX8414)
--	WX8417 = DFF(WX8416)
--	WX8419 = DFF(WX8418)
--	WX8421 = DFF(WX8420)
--	WX8423 = DFF(WX8422)
--	WX8425 = DFF(WX8424)
--	WX8427 = DFF(WX8426)
--	WX8429 = DFF(WX8428)
--	WX8431 = DFF(WX8430)
--	WX8433 = DFF(WX8432)
--	WX8435 = DFF(WX8434)
--	WX8437 = DFF(WX8436)
--	WX8439 = DFF(WX8438)
--	WX8441 = DFF(WX8440)
--	WX8443 = DFF(WX8442)
--	WX8445 = DFF(WX8444)
--	WX8447 = DFF(WX8446)
--	WX8449 = DFF(WX8448)
--	WX8451 = DFF(WX8450)
--	WX8453 = DFF(WX8452)
--	WX8455 = DFF(WX8454)
--	WX8457 = DFF(WX8456)
--	WX8459 = DFF(WX8458)
--	WX8461 = DFF(WX8460)
--	WX8463 = DFF(WX8462)
--	WX8465 = DFF(WX8464)
--	WX8467 = DFF(WX8466)
--	WX8469 = DFF(WX8468)
--	WX8471 = DFF(WX8470)
--	WX8473 = DFF(WX8472)
--	WX8475 = DFF(WX8474)
--	WX8477 = DFF(WX8476)
--	WX8479 = DFF(WX8478)
--	WX8481 = DFF(WX8480)
--	WX8483 = DFF(WX8482)
--	WX8485 = DFF(WX8484)
--	WX8487 = DFF(WX8486)
--	WX8489 = DFF(WX8488)
--	WX8491 = DFF(WX8490)
--	WX8493 = DFF(WX8492)
--	WX8495 = DFF(WX8494)
--	WX8497 = DFF(WX8496)
--	WX8499 = DFF(WX8498)
--	WX8501 = DFF(WX8500)
--	WX8503 = DFF(WX8502)
--	WX8505 = DFF(WX8504)
--	WX8507 = DFF(WX8506)
--	WX8509 = DFF(WX8508)
--	WX8511 = DFF(WX8510)
--	WX8513 = DFF(WX8512)
--	WX8515 = DFF(WX8514)
--	WX8517 = DFF(WX8516)
--	WX8519 = DFF(WX8518)
--	WX8521 = DFF(WX8520)
--	WX8523 = DFF(WX8522)
--	WX8525 = DFF(WX8524)
--	WX8527 = DFF(WX8526)
--	WX8529 = DFF(WX8528)
--	WX8531 = DFF(WX8530)
--	WX8533 = DFF(WX8532)
--	WX8535 = DFF(WX8534)
--	WX8537 = DFF(WX8536)
--	WX8539 = DFF(WX8538)
--	WX8541 = DFF(WX8540)
--	WX8543 = DFF(WX8542)
--	WX8545 = DFF(WX8544)
--	WX8547 = DFF(WX8546)
--	WX8549 = DFF(WX8548)
--	WX8551 = DFF(WX8550)
--	WX8553 = DFF(WX8552)
--	WX8555 = DFF(WX8554)
--	WX8557 = DFF(WX8556)
--	WX8559 = DFF(WX8558)
--	WX8561 = DFF(WX8560)
--	WX8563 = DFF(WX8562)
--	WX8565 = DFF(WX8564)
--	WX8567 = DFF(WX8566)
--	WX8569 = DFF(WX8568)
--	WX8571 = DFF(WX8570)
--	WX8573 = DFF(WX8572)
--	WX8575 = DFF(WX8574)
--	WX8577 = DFF(WX8576)
--	WX8579 = DFF(WX8578)
--	WX8581 = DFF(WX8580)
--	WX8583 = DFF(WX8582)
--	WX8585 = DFF(WX8584)
--	WX8587 = DFF(WX8586)
--	WX8589 = DFF(WX8588)
--	WX8591 = DFF(WX8590)
--	WX8593 = DFF(WX8592)
--	WX8595 = DFF(WX8594)
--	WX8597 = DFF(WX8596)
--	WX8599 = DFF(WX8598)
--	WX8601 = DFF(WX8600)
--	WX8603 = DFF(WX8602)
--	WX8605 = DFF(WX8604)
--	WX8607 = DFF(WX8606)
--	WX8609 = DFF(WX8608)
--	WX8611 = DFF(WX8610)
--	WX8613 = DFF(WX8612)
--	WX8615 = DFF(WX8614)
--	WX8617 = DFF(WX8616)
--	WX8619 = DFF(WX8618)
--	WX8621 = DFF(WX8620)
--	WX8623 = DFF(WX8622)
--	WX8625 = DFF(WX8624)
--	WX8627 = DFF(WX8626)
--	WX8629 = DFF(WX8628)
--	WX8631 = DFF(WX8630)
--	WX8633 = DFF(WX8632)
--	WX8635 = DFF(WX8634)
--	WX8637 = DFF(WX8636)
--	WX8639 = DFF(WX8638)
--	WX8641 = DFF(WX8640)
--	WX8643 = DFF(WX8642)
--	WX8645 = DFF(WX8644)
--	WX8647 = DFF(WX8646)
--	WX8649 = DFF(WX8648)
--	WX8651 = DFF(WX8650)
--	WX8653 = DFF(WX8652)
--	WX8655 = DFF(WX8654)
--	WX8657 = DFF(WX8656)
--	CRC_OUT_3_0 = DFF(WX9022)
--	CRC_OUT_3_1 = DFF(WX9024)
--	CRC_OUT_3_2 = DFF(WX9026)
--	CRC_OUT_3_3 = DFF(WX9028)
--	CRC_OUT_3_4 = DFF(WX9030)
--	CRC_OUT_3_5 = DFF(WX9032)
--	CRC_OUT_3_6 = DFF(WX9034)
--	CRC_OUT_3_7 = DFF(WX9036)
--	CRC_OUT_3_8 = DFF(WX9038)
--	CRC_OUT_3_9 = DFF(WX9040)
--	CRC_OUT_3_10 = DFF(WX9042)
--	CRC_OUT_3_11 = DFF(WX9044)
--	CRC_OUT_3_12 = DFF(WX9046)
--	CRC_OUT_3_13 = DFF(WX9048)
--	CRC_OUT_3_14 = DFF(WX9050)
--	CRC_OUT_3_15 = DFF(WX9052)
--	CRC_OUT_3_16 = DFF(WX9054)
--	CRC_OUT_3_17 = DFF(WX9056)
--	CRC_OUT_3_18 = DFF(WX9058)
--	CRC_OUT_3_19 = DFF(WX9060)
--	CRC_OUT_3_20 = DFF(WX9062)
--	CRC_OUT_3_21 = DFF(WX9064)
--	CRC_OUT_3_22 = DFF(WX9066)
--	CRC_OUT_3_23 = DFF(WX9068)
--	CRC_OUT_3_24 = DFF(WX9070)
--	CRC_OUT_3_25 = DFF(WX9072)
--	CRC_OUT_3_26 = DFF(WX9074)
--	CRC_OUT_3_27 = DFF(WX9076)
--	CRC_OUT_3_28 = DFF(WX9078)
--	CRC_OUT_3_29 = DFF(WX9080)
--	CRC_OUT_3_30 = DFF(WX9082)
--	CRC_OUT_3_31 = DFF(WX9084)
--	WX9536 = DFF(WX9535)
--	WX9538 = DFF(WX9537)
--	WX9540 = DFF(WX9539)
--	WX9542 = DFF(WX9541)
--	WX9544 = DFF(WX9543)
--	WX9546 = DFF(WX9545)
--	WX9548 = DFF(WX9547)
--	WX9550 = DFF(WX9549)
--	WX9552 = DFF(WX9551)
--	WX9554 = DFF(WX9553)
--	WX9556 = DFF(WX9555)
--	WX9558 = DFF(WX9557)
--	WX9560 = DFF(WX9559)
--	WX9562 = DFF(WX9561)
--	WX9564 = DFF(WX9563)
--	WX9566 = DFF(WX9565)
--	WX9568 = DFF(WX9567)
--	WX9570 = DFF(WX9569)
--	WX9572 = DFF(WX9571)
--	WX9574 = DFF(WX9573)
--	WX9576 = DFF(WX9575)
--	WX9578 = DFF(WX9577)
--	WX9580 = DFF(WX9579)
--	WX9582 = DFF(WX9581)
--	WX9584 = DFF(WX9583)
--	WX9586 = DFF(WX9585)
--	WX9588 = DFF(WX9587)
--	WX9590 = DFF(WX9589)
--	WX9592 = DFF(WX9591)
--	WX9594 = DFF(WX9593)
--	WX9596 = DFF(WX9595)
--	WX9598 = DFF(WX9597)
--	WX9696 = DFF(WX9695)
--	WX9698 = DFF(WX9697)
--	WX9700 = DFF(WX9699)
--	WX9702 = DFF(WX9701)
--	WX9704 = DFF(WX9703)
--	WX9706 = DFF(WX9705)
--	WX9708 = DFF(WX9707)
--	WX9710 = DFF(WX9709)
--	WX9712 = DFF(WX9711)
--	WX9714 = DFF(WX9713)
--	WX9716 = DFF(WX9715)
--	WX9718 = DFF(WX9717)
--	WX9720 = DFF(WX9719)
--	WX9722 = DFF(WX9721)
--	WX9724 = DFF(WX9723)
--	WX9726 = DFF(WX9725)
--	WX9728 = DFF(WX9727)
--	WX9730 = DFF(WX9729)
--	WX9732 = DFF(WX9731)
--	WX9734 = DFF(WX9733)
--	WX9736 = DFF(WX9735)
--	WX9738 = DFF(WX9737)
--	WX9740 = DFF(WX9739)
--	WX9742 = DFF(WX9741)
--	WX9744 = DFF(WX9743)
--	WX9746 = DFF(WX9745)
--	WX9748 = DFF(WX9747)
--	WX9750 = DFF(WX9749)
--	WX9752 = DFF(WX9751)
--	WX9754 = DFF(WX9753)
--	WX9756 = DFF(WX9755)
--	WX9758 = DFF(WX9757)
--	WX9760 = DFF(WX9759)
--	WX9762 = DFF(WX9761)
--	WX9764 = DFF(WX9763)
--	WX9766 = DFF(WX9765)
--	WX9768 = DFF(WX9767)
--	WX9770 = DFF(WX9769)
--	WX9772 = DFF(WX9771)
--	WX9774 = DFF(WX9773)
--	WX9776 = DFF(WX9775)
--	WX9778 = DFF(WX9777)
--	WX9780 = DFF(WX9779)
--	WX9782 = DFF(WX9781)
--	WX9784 = DFF(WX9783)
--	WX9786 = DFF(WX9785)
--	WX9788 = DFF(WX9787)
--	WX9790 = DFF(WX9789)
--	WX9792 = DFF(WX9791)
--	WX9794 = DFF(WX9793)
--	WX9796 = DFF(WX9795)
--	WX9798 = DFF(WX9797)
--	WX9800 = DFF(WX9799)
--	WX9802 = DFF(WX9801)
--	WX9804 = DFF(WX9803)
--	WX9806 = DFF(WX9805)
--	WX9808 = DFF(WX9807)
--	WX9810 = DFF(WX9809)
--	WX9812 = DFF(WX9811)
--	WX9814 = DFF(WX9813)
--	WX9816 = DFF(WX9815)
--	WX9818 = DFF(WX9817)
--	WX9820 = DFF(WX9819)
--	WX9822 = DFF(WX9821)
--	WX9824 = DFF(WX9823)
--	WX9826 = DFF(WX9825)
--	WX9828 = DFF(WX9827)
--	WX9830 = DFF(WX9829)
--	WX9832 = DFF(WX9831)
--	WX9834 = DFF(WX9833)
--	WX9836 = DFF(WX9835)
--	WX9838 = DFF(WX9837)
--	WX9840 = DFF(WX9839)
--	WX9842 = DFF(WX9841)
--	WX9844 = DFF(WX9843)
--	WX9846 = DFF(WX9845)
--	WX9848 = DFF(WX9847)
--	WX9850 = DFF(WX9849)
--	WX9852 = DFF(WX9851)
--	WX9854 = DFF(WX9853)
--	WX9856 = DFF(WX9855)
--	WX9858 = DFF(WX9857)
--	WX9860 = DFF(WX9859)
--	WX9862 = DFF(WX9861)
--	WX9864 = DFF(WX9863)
--	WX9866 = DFF(WX9865)
--	WX9868 = DFF(WX9867)
--	WX9870 = DFF(WX9869)
--	WX9872 = DFF(WX9871)
--	WX9874 = DFF(WX9873)
--	WX9876 = DFF(WX9875)
--	WX9878 = DFF(WX9877)
--	WX9880 = DFF(WX9879)
--	WX9882 = DFF(WX9881)
--	WX9884 = DFF(WX9883)
--	WX9886 = DFF(WX9885)
--	WX9888 = DFF(WX9887)
--	WX9890 = DFF(WX9889)
--	WX9892 = DFF(WX9891)
--	WX9894 = DFF(WX9893)
--	WX9896 = DFF(WX9895)
--	WX9898 = DFF(WX9897)
--	WX9900 = DFF(WX9899)
--	WX9902 = DFF(WX9901)
--	WX9904 = DFF(WX9903)
--	WX9906 = DFF(WX9905)
--	WX9908 = DFF(WX9907)
--	WX9910 = DFF(WX9909)
--	WX9912 = DFF(WX9911)
--	WX9914 = DFF(WX9913)
--	WX9916 = DFF(WX9915)
--	WX9918 = DFF(WX9917)
--	WX9920 = DFF(WX9919)
--	WX9922 = DFF(WX9921)
--	WX9924 = DFF(WX9923)
--	WX9926 = DFF(WX9925)
--	WX9928 = DFF(WX9927)
--	WX9930 = DFF(WX9929)
--	WX9932 = DFF(WX9931)
--	WX9934 = DFF(WX9933)
--	WX9936 = DFF(WX9935)
--	WX9938 = DFF(WX9937)
--	WX9940 = DFF(WX9939)
--	WX9942 = DFF(WX9941)
--	WX9944 = DFF(WX9943)
--	WX9946 = DFF(WX9945)
--	WX9948 = DFF(WX9947)
--	WX9950 = DFF(WX9949)
--	CRC_OUT_2_0 = DFF(WX10315)
--	CRC_OUT_2_1 = DFF(WX10317)
--	CRC_OUT_2_2 = DFF(WX10319)
--	CRC_OUT_2_3 = DFF(WX10321)
--	CRC_OUT_2_4 = DFF(WX10323)
--	CRC_OUT_2_5 = DFF(WX10325)
--	CRC_OUT_2_6 = DFF(WX10327)
--	CRC_OUT_2_7 = DFF(WX10329)
--	CRC_OUT_2_8 = DFF(WX10331)
--	CRC_OUT_2_9 = DFF(WX10333)
--	CRC_OUT_2_10 = DFF(WX10335)
--	CRC_OUT_2_11 = DFF(WX10337)
--	CRC_OUT_2_12 = DFF(WX10339)
--	CRC_OUT_2_13 = DFF(WX10341)
--	CRC_OUT_2_14 = DFF(WX10343)
--	CRC_OUT_2_15 = DFF(WX10345)
--	CRC_OUT_2_16 = DFF(WX10347)
--	CRC_OUT_2_17 = DFF(WX10349)
--	CRC_OUT_2_18 = DFF(WX10351)
--	CRC_OUT_2_19 = DFF(WX10353)
--	CRC_OUT_2_20 = DFF(WX10355)
--	CRC_OUT_2_21 = DFF(WX10357)
--	CRC_OUT_2_22 = DFF(WX10359)
--	CRC_OUT_2_23 = DFF(WX10361)
--	CRC_OUT_2_24 = DFF(WX10363)
--	CRC_OUT_2_25 = DFF(WX10365)
--	CRC_OUT_2_26 = DFF(WX10367)
--	CRC_OUT_2_27 = DFF(WX10369)
--	CRC_OUT_2_28 = DFF(WX10371)
--	CRC_OUT_2_29 = DFF(WX10373)
--	CRC_OUT_2_30 = DFF(WX10375)
--	CRC_OUT_2_31 = DFF(WX10377)
--	WX10829 = DFF(WX10828)
--	WX10831 = DFF(WX10830)
--	WX10833 = DFF(WX10832)
--	WX10835 = DFF(WX10834)
--	WX10837 = DFF(WX10836)
--	WX10839 = DFF(WX10838)
--	WX10841 = DFF(WX10840)
--	WX10843 = DFF(WX10842)
--	WX10845 = DFF(WX10844)
--	WX10847 = DFF(WX10846)
--	WX10849 = DFF(WX10848)
--	WX10851 = DFF(WX10850)
--	WX10853 = DFF(WX10852)
--	WX10855 = DFF(WX10854)
--	WX10857 = DFF(WX10856)
--	WX10859 = DFF(WX10858)
--	WX10861 = DFF(WX10860)
--	WX10863 = DFF(WX10862)
--	WX10865 = DFF(WX10864)
--	WX10867 = DFF(WX10866)
--	WX10869 = DFF(WX10868)
--	WX10871 = DFF(WX10870)
--	WX10873 = DFF(WX10872)
--	WX10875 = DFF(WX10874)
--	WX10877 = DFF(WX10876)
--	WX10879 = DFF(WX10878)
--	WX10881 = DFF(WX10880)
--	WX10883 = DFF(WX10882)
--	WX10885 = DFF(WX10884)
--	WX10887 = DFF(WX10886)
--	WX10889 = DFF(WX10888)
--	WX10891 = DFF(WX10890)
--	WX10989 = DFF(WX10988)
--	WX10991 = DFF(WX10990)
--	WX10993 = DFF(WX10992)
--	WX10995 = DFF(WX10994)
--	WX10997 = DFF(WX10996)
--	WX10999 = DFF(WX10998)
--	WX11001 = DFF(WX11000)
--	WX11003 = DFF(WX11002)
--	WX11005 = DFF(WX11004)
--	WX11007 = DFF(WX11006)
--	WX11009 = DFF(WX11008)
--	WX11011 = DFF(WX11010)
--	WX11013 = DFF(WX11012)
--	WX11015 = DFF(WX11014)
--	WX11017 = DFF(WX11016)
--	WX11019 = DFF(WX11018)
--	WX11021 = DFF(WX11020)
--	WX11023 = DFF(WX11022)
--	WX11025 = DFF(WX11024)
--	WX11027 = DFF(WX11026)
--	WX11029 = DFF(WX11028)
--	WX11031 = DFF(WX11030)
--	WX11033 = DFF(WX11032)
--	WX11035 = DFF(WX11034)
--	WX11037 = DFF(WX11036)
--	WX11039 = DFF(WX11038)
--	WX11041 = DFF(WX11040)
--	WX11043 = DFF(WX11042)
--	WX11045 = DFF(WX11044)
--	WX11047 = DFF(WX11046)
--	WX11049 = DFF(WX11048)
--	WX11051 = DFF(WX11050)
--	WX11053 = DFF(WX11052)
--	WX11055 = DFF(WX11054)
--	WX11057 = DFF(WX11056)
--	WX11059 = DFF(WX11058)
--	WX11061 = DFF(WX11060)
--	WX11063 = DFF(WX11062)
--	WX11065 = DFF(WX11064)
--	WX11067 = DFF(WX11066)
--	WX11069 = DFF(WX11068)
--	WX11071 = DFF(WX11070)
--	WX11073 = DFF(WX11072)
--	WX11075 = DFF(WX11074)
--	WX11077 = DFF(WX11076)
--	WX11079 = DFF(WX11078)
--	WX11081 = DFF(WX11080)
--	WX11083 = DFF(WX11082)
--	WX11085 = DFF(WX11084)
--	WX11087 = DFF(WX11086)
--	WX11089 = DFF(WX11088)
--	WX11091 = DFF(WX11090)
--	WX11093 = DFF(WX11092)
--	WX11095 = DFF(WX11094)
--	WX11097 = DFF(WX11096)
--	WX11099 = DFF(WX11098)
--	WX11101 = DFF(WX11100)
--	WX11103 = DFF(WX11102)
--	WX11105 = DFF(WX11104)
--	WX11107 = DFF(WX11106)
--	WX11109 = DFF(WX11108)
--	WX11111 = DFF(WX11110)
--	WX11113 = DFF(WX11112)
--	WX11115 = DFF(WX11114)
--	WX11117 = DFF(WX11116)
--	WX11119 = DFF(WX11118)
--	WX11121 = DFF(WX11120)
--	WX11123 = DFF(WX11122)
--	WX11125 = DFF(WX11124)
--	WX11127 = DFF(WX11126)
--	WX11129 = DFF(WX11128)
--	WX11131 = DFF(WX11130)
--	WX11133 = DFF(WX11132)
--	WX11135 = DFF(WX11134)
--	WX11137 = DFF(WX11136)
--	WX11139 = DFF(WX11138)
--	WX11141 = DFF(WX11140)
--	WX11143 = DFF(WX11142)
--	WX11145 = DFF(WX11144)
--	WX11147 = DFF(WX11146)
--	WX11149 = DFF(WX11148)
--	WX11151 = DFF(WX11150)
--	WX11153 = DFF(WX11152)
--	WX11155 = DFF(WX11154)
--	WX11157 = DFF(WX11156)
--	WX11159 = DFF(WX11158)
--	WX11161 = DFF(WX11160)
--	WX11163 = DFF(WX11162)
--	WX11165 = DFF(WX11164)
--	WX11167 = DFF(WX11166)
--	WX11169 = DFF(WX11168)
--	WX11171 = DFF(WX11170)
--	WX11173 = DFF(WX11172)
--	WX11175 = DFF(WX11174)
--	WX11177 = DFF(WX11176)
--	WX11179 = DFF(WX11178)
--	WX11181 = DFF(WX11180)
--	WX11183 = DFF(WX11182)
--	WX11185 = DFF(WX11184)
--	WX11187 = DFF(WX11186)
--	WX11189 = DFF(WX11188)
--	WX11191 = DFF(WX11190)
--	WX11193 = DFF(WX11192)
--	WX11195 = DFF(WX11194)
--	WX11197 = DFF(WX11196)
--	WX11199 = DFF(WX11198)
--	WX11201 = DFF(WX11200)
--	WX11203 = DFF(WX11202)
--	WX11205 = DFF(WX11204)
--	WX11207 = DFF(WX11206)
--	WX11209 = DFF(WX11208)
--	WX11211 = DFF(WX11210)
--	WX11213 = DFF(WX11212)
--	WX11215 = DFF(WX11214)
--	WX11217 = DFF(WX11216)
--	WX11219 = DFF(WX11218)
--	WX11221 = DFF(WX11220)
--	WX11223 = DFF(WX11222)
--	WX11225 = DFF(WX11224)
--	WX11227 = DFF(WX11226)
--	WX11229 = DFF(WX11228)
--	WX11231 = DFF(WX11230)
--	WX11233 = DFF(WX11232)
--	WX11235 = DFF(WX11234)
--	WX11237 = DFF(WX11236)
--	WX11239 = DFF(WX11238)
--	WX11241 = DFF(WX11240)
--	WX11243 = DFF(WX11242)
--	CRC_OUT_1_0 = DFF(WX11608)
--	CRC_OUT_1_1 = DFF(WX11610)
--	CRC_OUT_1_2 = DFF(WX11612)
--	CRC_OUT_1_3 = DFF(WX11614)
--	CRC_OUT_1_4 = DFF(WX11616)
--	CRC_OUT_1_5 = DFF(WX11618)
--	CRC_OUT_1_6 = DFF(WX11620)
--	CRC_OUT_1_7 = DFF(WX11622)
--	CRC_OUT_1_8 = DFF(WX11624)
--	CRC_OUT_1_9 = DFF(WX11626)
--	CRC_OUT_1_10 = DFF(WX11628)
--	CRC_OUT_1_11 = DFF(WX11630)
--	CRC_OUT_1_12 = DFF(WX11632)
--	CRC_OUT_1_13 = DFF(WX11634)
--	CRC_OUT_1_14 = DFF(WX11636)
--	CRC_OUT_1_15 = DFF(WX11638)
--	CRC_OUT_1_16 = DFF(WX11640)
--	CRC_OUT_1_17 = DFF(WX11642)
--	CRC_OUT_1_18 = DFF(WX11644)
--	CRC_OUT_1_19 = DFF(WX11646)
--	CRC_OUT_1_20 = DFF(WX11648)
--	CRC_OUT_1_21 = DFF(WX11650)
--	CRC_OUT_1_22 = DFF(WX11652)
--	CRC_OUT_1_23 = DFF(WX11654)
--	CRC_OUT_1_24 = DFF(WX11656)
--	CRC_OUT_1_25 = DFF(WX11658)
--	CRC_OUT_1_26 = DFF(WX11660)
--	CRC_OUT_1_27 = DFF(WX11662)
--	CRC_OUT_1_28 = DFF(WX11664)
--	CRC_OUT_1_29 = DFF(WX11666)
--	CRC_OUT_1_30 = DFF(WX11668)
--	CRC_OUT_1_31 = DFF(WX11670)
--	
--	WX37 = NOT(WX1003)
--	WX41 = NOT(WX1004)
--	WX45 = NOT(WX1004)
--	WX47 = NOT(WX38)
--	WX48 = NOT(WX47)
--	WX51 = NOT(WX1003)
--	WX55 = NOT(WX1004)
--	WX59 = NOT(WX1004)
--	WX61 = NOT(WX52)
--	WX62 = NOT(WX61)
--	WX65 = NOT(WX1003)
--	WX69 = NOT(WX1004)
--	WX73 = NOT(WX1004)
--	WX75 = NOT(WX66)
--	WX76 = NOT(WX75)
--	WX79 = NOT(WX1003)
--	WX83 = NOT(WX1004)
--	WX87 = NOT(WX1004)
--	WX89 = NOT(WX80)
--	WX90 = NOT(WX89)
--	WX93 = NOT(WX1003)
--	WX97 = NOT(WX1004)
--	WX101 = NOT(WX1004)
--	WX103 = NOT(WX94)
--	WX104 = NOT(WX103)
--	WX107 = NOT(WX1003)
--	WX111 = NOT(WX1004)
--	WX115 = NOT(WX1004)
--	WX117 = NOT(WX108)
--	WX118 = NOT(WX117)
--	WX121 = NOT(WX1003)
--	WX125 = NOT(WX1004)
--	WX129 = NOT(WX1004)
--	WX131 = NOT(WX122)
--	WX132 = NOT(WX131)
--	WX135 = NOT(WX1003)
--	WX139 = NOT(WX1004)
--	WX143 = NOT(WX1004)
--	WX145 = NOT(WX136)
--	WX146 = NOT(WX145)
--	WX149 = NOT(WX1003)
--	WX153 = NOT(WX1004)
--	WX157 = NOT(WX1004)
--	WX159 = NOT(WX150)
--	WX160 = NOT(WX159)
--	WX163 = NOT(WX1003)
--	WX167 = NOT(WX1004)
--	WX171 = NOT(WX1004)
--	WX173 = NOT(WX164)
--	WX174 = NOT(WX173)
--	WX177 = NOT(WX1003)
--	WX181 = NOT(WX1004)
--	WX185 = NOT(WX1004)
--	WX187 = NOT(WX178)
--	WX188 = NOT(WX187)
--	WX191 = NOT(WX1003)
--	WX195 = NOT(WX1004)
--	WX199 = NOT(WX1004)
--	WX201 = NOT(WX192)
--	WX202 = NOT(WX201)
--	WX205 = NOT(WX1003)
--	WX209 = NOT(WX1004)
--	WX213 = NOT(WX1004)
--	WX215 = NOT(WX206)
--	WX216 = NOT(WX215)
--	WX219 = NOT(WX1003)
--	WX223 = NOT(WX1004)
--	WX227 = NOT(WX1004)
--	WX229 = NOT(WX220)
--	WX230 = NOT(WX229)
--	WX233 = NOT(WX1003)
--	WX237 = NOT(WX1004)
--	WX241 = NOT(WX1004)
--	WX243 = NOT(WX234)
--	WX244 = NOT(WX243)
--	WX247 = NOT(WX1003)
--	WX251 = NOT(WX1004)
--	WX255 = NOT(WX1004)
--	WX257 = NOT(WX248)
--	WX258 = NOT(WX257)
--	WX261 = NOT(WX1003)
--	WX265 = NOT(WX1004)
--	WX269 = NOT(WX1004)
--	WX271 = NOT(WX262)
--	WX272 = NOT(WX271)
--	WX275 = NOT(WX1003)
--	WX279 = NOT(WX1004)
--	WX283 = NOT(WX1004)
--	WX285 = NOT(WX276)
--	WX286 = NOT(WX285)
--	WX289 = NOT(WX1003)
--	WX293 = NOT(WX1004)
--	WX297 = NOT(WX1004)
--	WX299 = NOT(WX290)
--	WX300 = NOT(WX299)
--	WX303 = NOT(WX1003)
--	WX307 = NOT(WX1004)
--	WX311 = NOT(WX1004)
--	WX313 = NOT(WX304)
--	WX314 = NOT(WX313)
--	WX317 = NOT(WX1003)
--	WX321 = NOT(WX1004)
--	WX325 = NOT(WX1004)
--	WX327 = NOT(WX318)
--	WX328 = NOT(WX327)
--	WX331 = NOT(WX1003)
--	WX335 = NOT(WX1004)
--	WX339 = NOT(WX1004)
--	WX341 = NOT(WX332)
--	WX342 = NOT(WX341)
--	WX345 = NOT(WX1003)
--	WX349 = NOT(WX1004)
--	WX353 = NOT(WX1004)
--	WX355 = NOT(WX346)
--	WX356 = NOT(WX355)
--	WX359 = NOT(WX1003)
--	WX363 = NOT(WX1004)
--	WX367 = NOT(WX1004)
--	WX369 = NOT(WX360)
--	WX370 = NOT(WX369)
--	WX373 = NOT(WX1003)
--	WX377 = NOT(WX1004)
--	WX381 = NOT(WX1004)
--	WX383 = NOT(WX374)
--	WX384 = NOT(WX383)
--	WX387 = NOT(WX1003)
--	WX391 = NOT(WX1004)
--	WX395 = NOT(WX1004)
--	WX397 = NOT(WX388)
--	WX398 = NOT(WX397)
--	WX401 = NOT(WX1003)
--	WX405 = NOT(WX1004)
--	WX409 = NOT(WX1004)
--	WX411 = NOT(WX402)
--	WX412 = NOT(WX411)
--	WX415 = NOT(WX1003)
--	WX419 = NOT(WX1004)
--	WX423 = NOT(WX1004)
--	WX425 = NOT(WX416)
--	WX426 = NOT(WX425)
--	WX429 = NOT(WX1003)
--	WX433 = NOT(WX1004)
--	WX437 = NOT(WX1004)
--	WX439 = NOT(WX430)
--	WX440 = NOT(WX439)
--	WX443 = NOT(WX1003)
--	WX447 = NOT(WX1004)
--	WX451 = NOT(WX1004)
--	WX453 = NOT(WX444)
--	WX454 = NOT(WX453)
--	WX457 = NOT(WX1003)
--	WX461 = NOT(WX1004)
--	WX465 = NOT(WX1004)
--	WX467 = NOT(WX458)
--	WX468 = NOT(WX467)
--	WX471 = NOT(WX1003)
--	WX475 = NOT(WX1004)
--	WX479 = NOT(WX1004)
--	WX481 = NOT(WX472)
--	WX482 = NOT(WX481)
--	WX483 = NOT(WX485)
--	WX548 = NOT(WX965)
--	WX549 = NOT(WX967)
--	WX550 = NOT(WX969)
--	WX551 = NOT(WX971)
--	WX552 = NOT(WX973)
--	WX553 = NOT(WX975)
--	WX554 = NOT(WX977)
--	WX555 = NOT(WX979)
--	WX556 = NOT(WX981)
--	WX557 = NOT(WX983)
--	WX558 = NOT(WX985)
--	WX559 = NOT(WX987)
--	WX560 = NOT(WX989)
--	WX561 = NOT(WX991)
--	WX562 = NOT(WX993)
--	WX563 = NOT(WX995)
--	WX564 = NOT(WX933)
--	WX565 = NOT(WX935)
--	WX566 = NOT(WX937)
--	WX567 = NOT(WX939)
--	WX568 = NOT(WX941)
--	WX569 = NOT(WX943)
--	WX570 = NOT(WX945)
--	WX571 = NOT(WX947)
--	WX572 = NOT(WX949)
--	WX573 = NOT(WX951)
--	WX574 = NOT(WX953)
--	WX575 = NOT(WX955)
--	WX576 = NOT(WX957)
--	WX577 = NOT(WX959)
--	WX578 = NOT(WX961)
--	WX579 = NOT(WX963)
--	WX580 = NOT(WX548)
--	WX581 = NOT(WX549)
--	WX582 = NOT(WX550)
--	WX583 = NOT(WX551)
--	WX584 = NOT(WX552)
--	WX585 = NOT(WX553)
--	WX586 = NOT(WX554)
--	WX587 = NOT(WX555)
--	WX588 = NOT(WX556)
--	WX589 = NOT(WX557)
--	WX590 = NOT(WX558)
--	WX591 = NOT(WX559)
--	WX592 = NOT(WX560)
--	WX593 = NOT(WX561)
--	WX594 = NOT(WX562)
--	WX595 = NOT(WX563)
--	WX596 = NOT(WX564)
--	WX597 = NOT(WX565)
--	WX598 = NOT(WX566)
--	WX599 = NOT(WX567)
--	WX600 = NOT(WX568)
--	WX601 = NOT(WX569)
--	WX602 = NOT(WX570)
--	WX603 = NOT(WX571)
--	WX604 = NOT(WX572)
--	WX605 = NOT(WX573)
--	WX606 = NOT(WX574)
--	WX607 = NOT(WX575)
--	WX608 = NOT(WX576)
--	WX609 = NOT(WX577)
--	WX610 = NOT(WX578)
--	WX611 = NOT(WX579)
--	WX612 = NOT(WX837)
--	WX613 = NOT(WX839)
--	WX614 = NOT(WX841)
--	WX615 = NOT(WX843)
--	WX616 = NOT(WX845)
--	WX617 = NOT(WX847)
--	WX618 = NOT(WX849)
--	WX619 = NOT(WX851)
--	WX620 = NOT(WX853)
--	WX621 = NOT(WX855)
--	WX622 = NOT(WX857)
--	WX623 = NOT(WX859)
--	WX624 = NOT(WX861)
--	WX625 = NOT(WX863)
--	WX626 = NOT(WX865)
--	WX627 = NOT(WX867)
--	WX628 = NOT(WX869)
--	WX629 = NOT(WX871)
--	WX630 = NOT(WX873)
--	WX631 = NOT(WX875)
--	WX632 = NOT(WX877)
--	WX633 = NOT(WX879)
--	WX634 = NOT(WX881)
--	WX635 = NOT(WX883)
--	WX636 = NOT(WX885)
--	WX637 = NOT(WX887)
--	WX638 = NOT(WX889)
--	WX639 = NOT(WX891)
--	WX640 = NOT(WX893)
--	WX641 = NOT(WX895)
--	WX642 = NOT(WX897)
--	WX643 = NOT(WX899)
--	WX932 = NOT(WX916)
--	WX933 = NOT(WX932)
--	WX934 = NOT(WX917)
--	WX935 = NOT(WX934)
--	WX936 = NOT(WX918)
--	WX937 = NOT(WX936)
--	WX938 = NOT(WX919)
--	WX939 = NOT(WX938)
--	WX940 = NOT(WX920)
--	WX941 = NOT(WX940)
--	WX942 = NOT(WX921)
--	WX943 = NOT(WX942)
--	WX944 = NOT(WX922)
--	WX945 = NOT(WX944)
--	WX946 = NOT(WX923)
--	WX947 = NOT(WX946)
--	WX948 = NOT(WX924)
--	WX949 = NOT(WX948)
--	WX950 = NOT(WX925)
--	WX951 = NOT(WX950)
--	WX952 = NOT(WX926)
--	WX953 = NOT(WX952)
--	WX954 = NOT(WX927)
--	WX955 = NOT(WX954)
--	WX956 = NOT(WX928)
--	WX957 = NOT(WX956)
--	WX958 = NOT(WX929)
--	WX959 = NOT(WX958)
--	WX960 = NOT(WX930)
--	WX961 = NOT(WX960)
--	WX962 = NOT(WX931)
--	WX963 = NOT(WX962)
--	WX964 = NOT(WX900)
--	WX965 = NOT(WX964)
--	WX966 = NOT(WX901)
--	WX967 = NOT(WX966)
--	WX968 = NOT(WX902)
--	WX969 = NOT(WX968)
--	WX970 = NOT(WX903)
--	WX971 = NOT(WX970)
--	WX972 = NOT(WX904)
--	WX973 = NOT(WX972)
--	WX974 = NOT(WX905)
--	WX975 = NOT(WX974)
--	WX976 = NOT(WX906)
--	WX977 = NOT(WX976)
--	WX978 = NOT(WX907)
--	WX979 = NOT(WX978)
--	WX980 = NOT(WX908)
--	WX981 = NOT(WX980)
--	WX982 = NOT(WX909)
--	WX983 = NOT(WX982)
--	WX984 = NOT(WX910)
--	WX985 = NOT(WX984)
--	WX986 = NOT(WX911)
--	WX987 = NOT(WX986)
--	WX988 = NOT(WX912)
--	WX989 = NOT(WX988)
--	WX990 = NOT(WX913)
--	WX991 = NOT(WX990)
--	WX992 = NOT(WX914)
--	WX993 = NOT(WX992)
--	WX994 = NOT(WX915)
--	WX995 = NOT(WX994)
--	WX996 = NOT(TM0)
--	WX997 = NOT(TM0)
--	WX998 = NOT(TM0)
--	WX999 = NOT(TM1)
--	WX1000 = NOT(TM1)
--	WX1001 = NOT(WX1000)
--	WX1002 = NOT(WX998)
--	WX1003 = NOT(WX999)
--	WX1004 = NOT(WX997)
--	WX1005 = NOT(WX996)
--	WX1009 = NOT(WX1005)
--	WX1011 = NOT(WX1010)
--	DATA_9_31 = NOT(WX1011)
--	WX1016 = NOT(WX1005)
--	WX1018 = NOT(WX1017)
--	DATA_9_30 = NOT(WX1018)
--	WX1023 = NOT(WX1005)
--	WX1025 = NOT(WX1024)
--	DATA_9_29 = NOT(WX1025)
--	WX1030 = NOT(WX1005)
--	WX1032 = NOT(WX1031)
--	DATA_9_28 = NOT(WX1032)
--	WX1037 = NOT(WX1005)
--	WX1039 = NOT(WX1038)
--	DATA_9_27 = NOT(WX1039)
--	WX1044 = NOT(WX1005)
--	WX1046 = NOT(WX1045)
--	DATA_9_26 = NOT(WX1046)
--	WX1051 = NOT(WX1005)
--	WX1053 = NOT(WX1052)
--	DATA_9_25 = NOT(WX1053)
--	WX1058 = NOT(WX1005)
--	WX1060 = NOT(WX1059)
--	DATA_9_24 = NOT(WX1060)
--	WX1065 = NOT(WX1005)
--	WX1067 = NOT(WX1066)
--	DATA_9_23 = NOT(WX1067)
--	WX1072 = NOT(WX1005)
--	WX1074 = NOT(WX1073)
--	DATA_9_22 = NOT(WX1074)
--	WX1079 = NOT(WX1005)
--	WX1081 = NOT(WX1080)
--	DATA_9_21 = NOT(WX1081)
--	WX1086 = NOT(WX1005)
--	WX1088 = NOT(WX1087)
--	DATA_9_20 = NOT(WX1088)
--	WX1093 = NOT(WX1005)
--	WX1095 = NOT(WX1094)
--	DATA_9_19 = NOT(WX1095)
--	WX1100 = NOT(WX1005)
--	WX1102 = NOT(WX1101)
--	DATA_9_18 = NOT(WX1102)
--	WX1107 = NOT(WX1005)
--	WX1109 = NOT(WX1108)
--	DATA_9_17 = NOT(WX1109)
--	WX1114 = NOT(WX1005)
--	WX1116 = NOT(WX1115)
--	DATA_9_16 = NOT(WX1116)
--	WX1121 = NOT(WX1005)
--	WX1123 = NOT(WX1122)
--	DATA_9_15 = NOT(WX1123)
--	WX1128 = NOT(WX1005)
--	WX1130 = NOT(WX1129)
--	DATA_9_14 = NOT(WX1130)
--	WX1135 = NOT(WX1005)
--	WX1137 = NOT(WX1136)
--	DATA_9_13 = NOT(WX1137)
--	WX1142 = NOT(WX1005)
--	WX1144 = NOT(WX1143)
--	DATA_9_12 = NOT(WX1144)
--	WX1149 = NOT(WX1005)
--	WX1151 = NOT(WX1150)
--	DATA_9_11 = NOT(WX1151)
--	WX1156 = NOT(WX1005)
--	WX1158 = NOT(WX1157)
--	DATA_9_10 = NOT(WX1158)
--	WX1163 = NOT(WX1005)
--	WX1165 = NOT(WX1164)
--	DATA_9_9 = NOT(WX1165)
--	WX1170 = NOT(WX1005)
--	WX1172 = NOT(WX1171)
--	DATA_9_8 = NOT(WX1172)
--	WX1177 = NOT(WX1005)
--	WX1179 = NOT(WX1178)
--	DATA_9_7 = NOT(WX1179)
--	WX1184 = NOT(WX1005)
--	WX1186 = NOT(WX1185)
--	DATA_9_6 = NOT(WX1186)
--	WX1191 = NOT(WX1005)
--	WX1193 = NOT(WX1192)
--	DATA_9_5 = NOT(WX1193)
--	WX1198 = NOT(WX1005)
--	WX1200 = NOT(WX1199)
--	DATA_9_4 = NOT(WX1200)
--	WX1205 = NOT(WX1005)
--	WX1207 = NOT(WX1206)
--	DATA_9_3 = NOT(WX1207)
--	WX1212 = NOT(WX1005)
--	WX1214 = NOT(WX1213)
--	DATA_9_2 = NOT(WX1214)
--	WX1219 = NOT(WX1005)
--	WX1221 = NOT(WX1220)
--	DATA_9_1 = NOT(WX1221)
--	WX1226 = NOT(WX1005)
--	WX1228 = NOT(WX1227)
--	DATA_9_0 = NOT(WX1228)
--	WX1230 = NOT(RESET)
--	WX1263 = NOT(WX1230)
--	WX1330 = NOT(WX2296)
--	WX1334 = NOT(WX2297)
--	WX1338 = NOT(WX2297)
--	WX1340 = NOT(WX1331)
--	WX1341 = NOT(WX1340)
--	WX1344 = NOT(WX2296)
--	WX1348 = NOT(WX2297)
--	WX1352 = NOT(WX2297)
--	WX1354 = NOT(WX1345)
--	WX1355 = NOT(WX1354)
--	WX1358 = NOT(WX2296)
--	WX1362 = NOT(WX2297)
--	WX1366 = NOT(WX2297)
--	WX1368 = NOT(WX1359)
--	WX1369 = NOT(WX1368)
--	WX1372 = NOT(WX2296)
--	WX1376 = NOT(WX2297)
--	WX1380 = NOT(WX2297)
--	WX1382 = NOT(WX1373)
--	WX1383 = NOT(WX1382)
--	WX1386 = NOT(WX2296)
--	WX1390 = NOT(WX2297)
--	WX1394 = NOT(WX2297)
--	WX1396 = NOT(WX1387)
--	WX1397 = NOT(WX1396)
--	WX1400 = NOT(WX2296)
--	WX1404 = NOT(WX2297)
--	WX1408 = NOT(WX2297)
--	WX1410 = NOT(WX1401)
--	WX1411 = NOT(WX1410)
--	WX1414 = NOT(WX2296)
--	WX1418 = NOT(WX2297)
--	WX1422 = NOT(WX2297)
--	WX1424 = NOT(WX1415)
--	WX1425 = NOT(WX1424)
--	WX1428 = NOT(WX2296)
--	WX1432 = NOT(WX2297)
--	WX1436 = NOT(WX2297)
--	WX1438 = NOT(WX1429)
--	WX1439 = NOT(WX1438)
--	WX1442 = NOT(WX2296)
--	WX1446 = NOT(WX2297)
--	WX1450 = NOT(WX2297)
--	WX1452 = NOT(WX1443)
--	WX1453 = NOT(WX1452)
--	WX1456 = NOT(WX2296)
--	WX1460 = NOT(WX2297)
--	WX1464 = NOT(WX2297)
--	WX1466 = NOT(WX1457)
--	WX1467 = NOT(WX1466)
--	WX1470 = NOT(WX2296)
--	WX1474 = NOT(WX2297)
--	WX1478 = NOT(WX2297)
--	WX1480 = NOT(WX1471)
--	WX1481 = NOT(WX1480)
--	WX1484 = NOT(WX2296)
--	WX1488 = NOT(WX2297)
--	WX1492 = NOT(WX2297)
--	WX1494 = NOT(WX1485)
--	WX1495 = NOT(WX1494)
--	WX1498 = NOT(WX2296)
--	WX1502 = NOT(WX2297)
--	WX1506 = NOT(WX2297)
--	WX1508 = NOT(WX1499)
--	WX1509 = NOT(WX1508)
--	WX1512 = NOT(WX2296)
--	WX1516 = NOT(WX2297)
--	WX1520 = NOT(WX2297)
--	WX1522 = NOT(WX1513)
--	WX1523 = NOT(WX1522)
--	WX1526 = NOT(WX2296)
--	WX1530 = NOT(WX2297)
--	WX1534 = NOT(WX2297)
--	WX1536 = NOT(WX1527)
--	WX1537 = NOT(WX1536)
--	WX1540 = NOT(WX2296)
--	WX1544 = NOT(WX2297)
--	WX1548 = NOT(WX2297)
--	WX1550 = NOT(WX1541)
--	WX1551 = NOT(WX1550)
--	WX1554 = NOT(WX2296)
--	WX1558 = NOT(WX2297)
--	WX1562 = NOT(WX2297)
--	WX1564 = NOT(WX1555)
--	WX1565 = NOT(WX1564)
--	WX1568 = NOT(WX2296)
--	WX1572 = NOT(WX2297)
--	WX1576 = NOT(WX2297)
--	WX1578 = NOT(WX1569)
--	WX1579 = NOT(WX1578)
--	WX1582 = NOT(WX2296)
--	WX1586 = NOT(WX2297)
--	WX1590 = NOT(WX2297)
--	WX1592 = NOT(WX1583)
--	WX1593 = NOT(WX1592)
--	WX1596 = NOT(WX2296)
--	WX1600 = NOT(WX2297)
--	WX1604 = NOT(WX2297)
--	WX1606 = NOT(WX1597)
--	WX1607 = NOT(WX1606)
--	WX1610 = NOT(WX2296)
--	WX1614 = NOT(WX2297)
--	WX1618 = NOT(WX2297)
--	WX1620 = NOT(WX1611)
--	WX1621 = NOT(WX1620)
--	WX1624 = NOT(WX2296)
--	WX1628 = NOT(WX2297)
--	WX1632 = NOT(WX2297)
--	WX1634 = NOT(WX1625)
--	WX1635 = NOT(WX1634)
--	WX1638 = NOT(WX2296)
--	WX1642 = NOT(WX2297)
--	WX1646 = NOT(WX2297)
--	WX1648 = NOT(WX1639)
--	WX1649 = NOT(WX1648)
--	WX1652 = NOT(WX2296)
--	WX1656 = NOT(WX2297)
--	WX1660 = NOT(WX2297)
--	WX1662 = NOT(WX1653)
--	WX1663 = NOT(WX1662)
--	WX1666 = NOT(WX2296)
--	WX1670 = NOT(WX2297)
--	WX1674 = NOT(WX2297)
--	WX1676 = NOT(WX1667)
--	WX1677 = NOT(WX1676)
--	WX1680 = NOT(WX2296)
--	WX1684 = NOT(WX2297)
--	WX1688 = NOT(WX2297)
--	WX1690 = NOT(WX1681)
--	WX1691 = NOT(WX1690)
--	WX1694 = NOT(WX2296)
--	WX1698 = NOT(WX2297)
--	WX1702 = NOT(WX2297)
--	WX1704 = NOT(WX1695)
--	WX1705 = NOT(WX1704)
--	WX1708 = NOT(WX2296)
--	WX1712 = NOT(WX2297)
--	WX1716 = NOT(WX2297)
--	WX1718 = NOT(WX1709)
--	WX1719 = NOT(WX1718)
--	WX1722 = NOT(WX2296)
--	WX1726 = NOT(WX2297)
--	WX1730 = NOT(WX2297)
--	WX1732 = NOT(WX1723)
--	WX1733 = NOT(WX1732)
--	WX1736 = NOT(WX2296)
--	WX1740 = NOT(WX2297)
--	WX1744 = NOT(WX2297)
--	WX1746 = NOT(WX1737)
--	WX1747 = NOT(WX1746)
--	WX1750 = NOT(WX2296)
--	WX1754 = NOT(WX2297)
--	WX1758 = NOT(WX2297)
--	WX1760 = NOT(WX1751)
--	WX1761 = NOT(WX1760)
--	WX1764 = NOT(WX2296)
--	WX1768 = NOT(WX2297)
--	WX1772 = NOT(WX2297)
--	WX1774 = NOT(WX1765)
--	WX1775 = NOT(WX1774)
--	WX1776 = NOT(WX1778)
--	WX1841 = NOT(WX2258)
--	WX1842 = NOT(WX2260)
--	WX1843 = NOT(WX2262)
--	WX1844 = NOT(WX2264)
--	WX1845 = NOT(WX2266)
--	WX1846 = NOT(WX2268)
--	WX1847 = NOT(WX2270)
--	WX1848 = NOT(WX2272)
--	WX1849 = NOT(WX2274)
--	WX1850 = NOT(WX2276)
--	WX1851 = NOT(WX2278)
--	WX1852 = NOT(WX2280)
--	WX1853 = NOT(WX2282)
--	WX1854 = NOT(WX2284)
--	WX1855 = NOT(WX2286)
--	WX1856 = NOT(WX2288)
--	WX1857 = NOT(WX2226)
--	WX1858 = NOT(WX2228)
--	WX1859 = NOT(WX2230)
--	WX1860 = NOT(WX2232)
--	WX1861 = NOT(WX2234)
--	WX1862 = NOT(WX2236)
--	WX1863 = NOT(WX2238)
--	WX1864 = NOT(WX2240)
--	WX1865 = NOT(WX2242)
--	WX1866 = NOT(WX2244)
--	WX1867 = NOT(WX2246)
--	WX1868 = NOT(WX2248)
--	WX1869 = NOT(WX2250)
--	WX1870 = NOT(WX2252)
--	WX1871 = NOT(WX2254)
--	WX1872 = NOT(WX2256)
--	WX1873 = NOT(WX1841)
--	WX1874 = NOT(WX1842)
--	WX1875 = NOT(WX1843)
--	WX1876 = NOT(WX1844)
--	WX1877 = NOT(WX1845)
--	WX1878 = NOT(WX1846)
--	WX1879 = NOT(WX1847)
--	WX1880 = NOT(WX1848)
--	WX1881 = NOT(WX1849)
--	WX1882 = NOT(WX1850)
--	WX1883 = NOT(WX1851)
--	WX1884 = NOT(WX1852)
--	WX1885 = NOT(WX1853)
--	WX1886 = NOT(WX1854)
--	WX1887 = NOT(WX1855)
--	WX1888 = NOT(WX1856)
--	WX1889 = NOT(WX1857)
--	WX1890 = NOT(WX1858)
--	WX1891 = NOT(WX1859)
--	WX1892 = NOT(WX1860)
--	WX1893 = NOT(WX1861)
--	WX1894 = NOT(WX1862)
--	WX1895 = NOT(WX1863)
--	WX1896 = NOT(WX1864)
--	WX1897 = NOT(WX1865)
--	WX1898 = NOT(WX1866)
--	WX1899 = NOT(WX1867)
--	WX1900 = NOT(WX1868)
--	WX1901 = NOT(WX1869)
--	WX1902 = NOT(WX1870)
--	WX1903 = NOT(WX1871)
--	WX1904 = NOT(WX1872)
--	WX1905 = NOT(WX2130)
--	WX1906 = NOT(WX2132)
--	WX1907 = NOT(WX2134)
--	WX1908 = NOT(WX2136)
--	WX1909 = NOT(WX2138)
--	WX1910 = NOT(WX2140)
--	WX1911 = NOT(WX2142)
--	WX1912 = NOT(WX2144)
--	WX1913 = NOT(WX2146)
--	WX1914 = NOT(WX2148)
--	WX1915 = NOT(WX2150)
--	WX1916 = NOT(WX2152)
--	WX1917 = NOT(WX2154)
--	WX1918 = NOT(WX2156)
--	WX1919 = NOT(WX2158)
--	WX1920 = NOT(WX2160)
--	WX1921 = NOT(WX2162)
--	WX1922 = NOT(WX2164)
--	WX1923 = NOT(WX2166)
--	WX1924 = NOT(WX2168)
--	WX1925 = NOT(WX2170)
--	WX1926 = NOT(WX2172)
--	WX1927 = NOT(WX2174)
--	WX1928 = NOT(WX2176)
--	WX1929 = NOT(WX2178)
--	WX1930 = NOT(WX2180)
--	WX1931 = NOT(WX2182)
--	WX1932 = NOT(WX2184)
--	WX1933 = NOT(WX2186)
--	WX1934 = NOT(WX2188)
--	WX1935 = NOT(WX2190)
--	WX1936 = NOT(WX2192)
--	WX2225 = NOT(WX2209)
--	WX2226 = NOT(WX2225)
--	WX2227 = NOT(WX2210)
--	WX2228 = NOT(WX2227)
--	WX2229 = NOT(WX2211)
--	WX2230 = NOT(WX2229)
--	WX2231 = NOT(WX2212)
--	WX2232 = NOT(WX2231)
--	WX2233 = NOT(WX2213)
--	WX2234 = NOT(WX2233)
--	WX2235 = NOT(WX2214)
--	WX2236 = NOT(WX2235)
--	WX2237 = NOT(WX2215)
--	WX2238 = NOT(WX2237)
--	WX2239 = NOT(WX2216)
--	WX2240 = NOT(WX2239)
--	WX2241 = NOT(WX2217)
--	WX2242 = NOT(WX2241)
--	WX2243 = NOT(WX2218)
--	WX2244 = NOT(WX2243)
--	WX2245 = NOT(WX2219)
--	WX2246 = NOT(WX2245)
--	WX2247 = NOT(WX2220)
--	WX2248 = NOT(WX2247)
--	WX2249 = NOT(WX2221)
--	WX2250 = NOT(WX2249)
--	WX2251 = NOT(WX2222)
--	WX2252 = NOT(WX2251)
--	WX2253 = NOT(WX2223)
--	WX2254 = NOT(WX2253)
--	WX2255 = NOT(WX2224)
--	WX2256 = NOT(WX2255)
--	WX2257 = NOT(WX2193)
--	WX2258 = NOT(WX2257)
--	WX2259 = NOT(WX2194)
--	WX2260 = NOT(WX2259)
--	WX2261 = NOT(WX2195)
--	WX2262 = NOT(WX2261)
--	WX2263 = NOT(WX2196)
--	WX2264 = NOT(WX2263)
--	WX2265 = NOT(WX2197)
--	WX2266 = NOT(WX2265)
--	WX2267 = NOT(WX2198)
--	WX2268 = NOT(WX2267)
--	WX2269 = NOT(WX2199)
--	WX2270 = NOT(WX2269)
--	WX2271 = NOT(WX2200)
--	WX2272 = NOT(WX2271)
--	WX2273 = NOT(WX2201)
--	WX2274 = NOT(WX2273)
--	WX2275 = NOT(WX2202)
--	WX2276 = NOT(WX2275)
--	WX2277 = NOT(WX2203)
--	WX2278 = NOT(WX2277)
--	WX2279 = NOT(WX2204)
--	WX2280 = NOT(WX2279)
--	WX2281 = NOT(WX2205)
--	WX2282 = NOT(WX2281)
--	WX2283 = NOT(WX2206)
--	WX2284 = NOT(WX2283)
--	WX2285 = NOT(WX2207)
--	WX2286 = NOT(WX2285)
--	WX2287 = NOT(WX2208)
--	WX2288 = NOT(WX2287)
--	WX2289 = NOT(TM0)
--	WX2290 = NOT(TM0)
--	WX2291 = NOT(TM0)
--	WX2292 = NOT(TM1)
--	WX2293 = NOT(TM1)
--	WX2294 = NOT(WX2293)
--	WX2295 = NOT(WX2291)
--	WX2296 = NOT(WX2292)
--	WX2297 = NOT(WX2290)
--	WX2298 = NOT(WX2289)
--	WX2302 = NOT(WX2298)
--	WX2304 = NOT(WX2303)
--	WX2305 = NOT(WX2304)
--	WX2309 = NOT(WX2298)
--	WX2311 = NOT(WX2310)
--	WX2312 = NOT(WX2311)
--	WX2316 = NOT(WX2298)
--	WX2318 = NOT(WX2317)
--	WX2319 = NOT(WX2318)
--	WX2323 = NOT(WX2298)
--	WX2325 = NOT(WX2324)
--	WX2326 = NOT(WX2325)
--	WX2330 = NOT(WX2298)
--	WX2332 = NOT(WX2331)
--	WX2333 = NOT(WX2332)
--	WX2337 = NOT(WX2298)
--	WX2339 = NOT(WX2338)
--	WX2340 = NOT(WX2339)
--	WX2344 = NOT(WX2298)
--	WX2346 = NOT(WX2345)
--	WX2347 = NOT(WX2346)
--	WX2351 = NOT(WX2298)
--	WX2353 = NOT(WX2352)
--	WX2354 = NOT(WX2353)
--	WX2358 = NOT(WX2298)
--	WX2360 = NOT(WX2359)
--	WX2361 = NOT(WX2360)
--	WX2365 = NOT(WX2298)
--	WX2367 = NOT(WX2366)
--	WX2368 = NOT(WX2367)
--	WX2372 = NOT(WX2298)
--	WX2374 = NOT(WX2373)
--	WX2375 = NOT(WX2374)
--	WX2379 = NOT(WX2298)
--	WX2381 = NOT(WX2380)
--	WX2382 = NOT(WX2381)
--	WX2386 = NOT(WX2298)
--	WX2388 = NOT(WX2387)
--	WX2389 = NOT(WX2388)
--	WX2393 = NOT(WX2298)
--	WX2395 = NOT(WX2394)
--	WX2396 = NOT(WX2395)
--	WX2400 = NOT(WX2298)
--	WX2402 = NOT(WX2401)
--	WX2403 = NOT(WX2402)
--	WX2407 = NOT(WX2298)
--	WX2409 = NOT(WX2408)
--	WX2410 = NOT(WX2409)
--	WX2414 = NOT(WX2298)
--	WX2416 = NOT(WX2415)
--	WX2417 = NOT(WX2416)
--	WX2421 = NOT(WX2298)
--	WX2423 = NOT(WX2422)
--	WX2424 = NOT(WX2423)
--	WX2428 = NOT(WX2298)
--	WX2430 = NOT(WX2429)
--	WX2431 = NOT(WX2430)
--	WX2435 = NOT(WX2298)
--	WX2437 = NOT(WX2436)
--	WX2438 = NOT(WX2437)
--	WX2442 = NOT(WX2298)
--	WX2444 = NOT(WX2443)
--	WX2445 = NOT(WX2444)
--	WX2449 = NOT(WX2298)
--	WX2451 = NOT(WX2450)
--	WX2452 = NOT(WX2451)
--	WX2456 = NOT(WX2298)
--	WX2458 = NOT(WX2457)
--	WX2459 = NOT(WX2458)
--	WX2463 = NOT(WX2298)
--	WX2465 = NOT(WX2464)
--	WX2466 = NOT(WX2465)
--	WX2470 = NOT(WX2298)
--	WX2472 = NOT(WX2471)
--	WX2473 = NOT(WX2472)
--	WX2477 = NOT(WX2298)
--	WX2479 = NOT(WX2478)
--	WX2480 = NOT(WX2479)
--	WX2484 = NOT(WX2298)
--	WX2486 = NOT(WX2485)
--	WX2487 = NOT(WX2486)
--	WX2491 = NOT(WX2298)
--	WX2493 = NOT(WX2492)
--	WX2494 = NOT(WX2493)
--	WX2498 = NOT(WX2298)
--	WX2500 = NOT(WX2499)
--	WX2501 = NOT(WX2500)
--	WX2505 = NOT(WX2298)
--	WX2507 = NOT(WX2506)
--	WX2508 = NOT(WX2507)
--	WX2512 = NOT(WX2298)
--	WX2514 = NOT(WX2513)
--	WX2515 = NOT(WX2514)
--	WX2519 = NOT(WX2298)
--	WX2521 = NOT(WX2520)
--	WX2522 = NOT(WX2521)
--	WX2523 = NOT(RESET)
--	WX2556 = NOT(WX2523)
--	WX2623 = NOT(WX3589)
--	WX2627 = NOT(WX3590)
--	WX2631 = NOT(WX3590)
--	WX2633 = NOT(WX2624)
--	WX2634 = NOT(WX2633)
--	WX2637 = NOT(WX3589)
--	WX2641 = NOT(WX3590)
--	WX2645 = NOT(WX3590)
--	WX2647 = NOT(WX2638)
--	WX2648 = NOT(WX2647)
--	WX2651 = NOT(WX3589)
--	WX2655 = NOT(WX3590)
--	WX2659 = NOT(WX3590)
--	WX2661 = NOT(WX2652)
--	WX2662 = NOT(WX2661)
--	WX2665 = NOT(WX3589)
--	WX2669 = NOT(WX3590)
--	WX2673 = NOT(WX3590)
--	WX2675 = NOT(WX2666)
--	WX2676 = NOT(WX2675)
--	WX2679 = NOT(WX3589)
--	WX2683 = NOT(WX3590)
--	WX2687 = NOT(WX3590)
--	WX2689 = NOT(WX2680)
--	WX2690 = NOT(WX2689)
--	WX2693 = NOT(WX3589)
--	WX2697 = NOT(WX3590)
--	WX2701 = NOT(WX3590)
--	WX2703 = NOT(WX2694)
--	WX2704 = NOT(WX2703)
--	WX2707 = NOT(WX3589)
--	WX2711 = NOT(WX3590)
--	WX2715 = NOT(WX3590)
--	WX2717 = NOT(WX2708)
--	WX2718 = NOT(WX2717)
--	WX2721 = NOT(WX3589)
--	WX2725 = NOT(WX3590)
--	WX2729 = NOT(WX3590)
--	WX2731 = NOT(WX2722)
--	WX2732 = NOT(WX2731)
--	WX2735 = NOT(WX3589)
--	WX2739 = NOT(WX3590)
--	WX2743 = NOT(WX3590)
--	WX2745 = NOT(WX2736)
--	WX2746 = NOT(WX2745)
--	WX2749 = NOT(WX3589)
--	WX2753 = NOT(WX3590)
--	WX2757 = NOT(WX3590)
--	WX2759 = NOT(WX2750)
--	WX2760 = NOT(WX2759)
--	WX2763 = NOT(WX3589)
--	WX2767 = NOT(WX3590)
--	WX2771 = NOT(WX3590)
--	WX2773 = NOT(WX2764)
--	WX2774 = NOT(WX2773)
--	WX2777 = NOT(WX3589)
--	WX2781 = NOT(WX3590)
--	WX2785 = NOT(WX3590)
--	WX2787 = NOT(WX2778)
--	WX2788 = NOT(WX2787)
--	WX2791 = NOT(WX3589)
--	WX2795 = NOT(WX3590)
--	WX2799 = NOT(WX3590)
--	WX2801 = NOT(WX2792)
--	WX2802 = NOT(WX2801)
--	WX2805 = NOT(WX3589)
--	WX2809 = NOT(WX3590)
--	WX2813 = NOT(WX3590)
--	WX2815 = NOT(WX2806)
--	WX2816 = NOT(WX2815)
--	WX2819 = NOT(WX3589)
--	WX2823 = NOT(WX3590)
--	WX2827 = NOT(WX3590)
--	WX2829 = NOT(WX2820)
--	WX2830 = NOT(WX2829)
--	WX2833 = NOT(WX3589)
--	WX2837 = NOT(WX3590)
--	WX2841 = NOT(WX3590)
--	WX2843 = NOT(WX2834)
--	WX2844 = NOT(WX2843)
--	WX2847 = NOT(WX3589)
--	WX2851 = NOT(WX3590)
--	WX2855 = NOT(WX3590)
--	WX2857 = NOT(WX2848)
--	WX2858 = NOT(WX2857)
--	WX2861 = NOT(WX3589)
--	WX2865 = NOT(WX3590)
--	WX2869 = NOT(WX3590)
--	WX2871 = NOT(WX2862)
--	WX2872 = NOT(WX2871)
--	WX2875 = NOT(WX3589)
--	WX2879 = NOT(WX3590)
--	WX2883 = NOT(WX3590)
--	WX2885 = NOT(WX2876)
--	WX2886 = NOT(WX2885)
--	WX2889 = NOT(WX3589)
--	WX2893 = NOT(WX3590)
--	WX2897 = NOT(WX3590)
--	WX2899 = NOT(WX2890)
--	WX2900 = NOT(WX2899)
--	WX2903 = NOT(WX3589)
--	WX2907 = NOT(WX3590)
--	WX2911 = NOT(WX3590)
--	WX2913 = NOT(WX2904)
--	WX2914 = NOT(WX2913)
--	WX2917 = NOT(WX3589)
--	WX2921 = NOT(WX3590)
--	WX2925 = NOT(WX3590)
--	WX2927 = NOT(WX2918)
--	WX2928 = NOT(WX2927)
--	WX2931 = NOT(WX3589)
--	WX2935 = NOT(WX3590)
--	WX2939 = NOT(WX3590)
--	WX2941 = NOT(WX2932)
--	WX2942 = NOT(WX2941)
--	WX2945 = NOT(WX3589)
--	WX2949 = NOT(WX3590)
--	WX2953 = NOT(WX3590)
--	WX2955 = NOT(WX2946)
--	WX2956 = NOT(WX2955)
--	WX2959 = NOT(WX3589)
--	WX2963 = NOT(WX3590)
--	WX2967 = NOT(WX3590)
--	WX2969 = NOT(WX2960)
--	WX2970 = NOT(WX2969)
--	WX2973 = NOT(WX3589)
--	WX2977 = NOT(WX3590)
--	WX2981 = NOT(WX3590)
--	WX2983 = NOT(WX2974)
--	WX2984 = NOT(WX2983)
--	WX2987 = NOT(WX3589)
--	WX2991 = NOT(WX3590)
--	WX2995 = NOT(WX3590)
--	WX2997 = NOT(WX2988)
--	WX2998 = NOT(WX2997)
--	WX3001 = NOT(WX3589)
--	WX3005 = NOT(WX3590)
--	WX3009 = NOT(WX3590)
--	WX3011 = NOT(WX3002)
--	WX3012 = NOT(WX3011)
--	WX3015 = NOT(WX3589)
--	WX3019 = NOT(WX3590)
--	WX3023 = NOT(WX3590)
--	WX3025 = NOT(WX3016)
--	WX3026 = NOT(WX3025)
--	WX3029 = NOT(WX3589)
--	WX3033 = NOT(WX3590)
--	WX3037 = NOT(WX3590)
--	WX3039 = NOT(WX3030)
--	WX3040 = NOT(WX3039)
--	WX3043 = NOT(WX3589)
--	WX3047 = NOT(WX3590)
--	WX3051 = NOT(WX3590)
--	WX3053 = NOT(WX3044)
--	WX3054 = NOT(WX3053)
--	WX3057 = NOT(WX3589)
--	WX3061 = NOT(WX3590)
--	WX3065 = NOT(WX3590)
--	WX3067 = NOT(WX3058)
--	WX3068 = NOT(WX3067)
--	WX3069 = NOT(WX3071)
--	WX3134 = NOT(WX3551)
--	WX3135 = NOT(WX3553)
--	WX3136 = NOT(WX3555)
--	WX3137 = NOT(WX3557)
--	WX3138 = NOT(WX3559)
--	WX3139 = NOT(WX3561)
--	WX3140 = NOT(WX3563)
--	WX3141 = NOT(WX3565)
--	WX3142 = NOT(WX3567)
--	WX3143 = NOT(WX3569)
--	WX3144 = NOT(WX3571)
--	WX3145 = NOT(WX3573)
--	WX3146 = NOT(WX3575)
--	WX3147 = NOT(WX3577)
--	WX3148 = NOT(WX3579)
--	WX3149 = NOT(WX3581)
--	WX3150 = NOT(WX3519)
--	WX3151 = NOT(WX3521)
--	WX3152 = NOT(WX3523)
--	WX3153 = NOT(WX3525)
--	WX3154 = NOT(WX3527)
--	WX3155 = NOT(WX3529)
--	WX3156 = NOT(WX3531)
--	WX3157 = NOT(WX3533)
--	WX3158 = NOT(WX3535)
--	WX3159 = NOT(WX3537)
--	WX3160 = NOT(WX3539)
--	WX3161 = NOT(WX3541)
--	WX3162 = NOT(WX3543)
--	WX3163 = NOT(WX3545)
--	WX3164 = NOT(WX3547)
--	WX3165 = NOT(WX3549)
--	WX3166 = NOT(WX3134)
--	WX3167 = NOT(WX3135)
--	WX3168 = NOT(WX3136)
--	WX3169 = NOT(WX3137)
--	WX3170 = NOT(WX3138)
--	WX3171 = NOT(WX3139)
--	WX3172 = NOT(WX3140)
--	WX3173 = NOT(WX3141)
--	WX3174 = NOT(WX3142)
--	WX3175 = NOT(WX3143)
--	WX3176 = NOT(WX3144)
--	WX3177 = NOT(WX3145)
--	WX3178 = NOT(WX3146)
--	WX3179 = NOT(WX3147)
--	WX3180 = NOT(WX3148)
--	WX3181 = NOT(WX3149)
--	WX3182 = NOT(WX3150)
--	WX3183 = NOT(WX3151)
--	WX3184 = NOT(WX3152)
--	WX3185 = NOT(WX3153)
--	WX3186 = NOT(WX3154)
--	WX3187 = NOT(WX3155)
--	WX3188 = NOT(WX3156)
--	WX3189 = NOT(WX3157)
--	WX3190 = NOT(WX3158)
--	WX3191 = NOT(WX3159)
--	WX3192 = NOT(WX3160)
--	WX3193 = NOT(WX3161)
--	WX3194 = NOT(WX3162)
--	WX3195 = NOT(WX3163)
--	WX3196 = NOT(WX3164)
--	WX3197 = NOT(WX3165)
--	WX3198 = NOT(WX3423)
--	WX3199 = NOT(WX3425)
--	WX3200 = NOT(WX3427)
--	WX3201 = NOT(WX3429)
--	WX3202 = NOT(WX3431)
--	WX3203 = NOT(WX3433)
--	WX3204 = NOT(WX3435)
--	WX3205 = NOT(WX3437)
--	WX3206 = NOT(WX3439)
--	WX3207 = NOT(WX3441)
--	WX3208 = NOT(WX3443)
--	WX3209 = NOT(WX3445)
--	WX3210 = NOT(WX3447)
--	WX3211 = NOT(WX3449)
--	WX3212 = NOT(WX3451)
--	WX3213 = NOT(WX3453)
--	WX3214 = NOT(WX3455)
--	WX3215 = NOT(WX3457)
--	WX3216 = NOT(WX3459)
--	WX3217 = NOT(WX3461)
--	WX3218 = NOT(WX3463)
--	WX3219 = NOT(WX3465)
--	WX3220 = NOT(WX3467)
--	WX3221 = NOT(WX3469)
--	WX3222 = NOT(WX3471)
--	WX3223 = NOT(WX3473)
--	WX3224 = NOT(WX3475)
--	WX3225 = NOT(WX3477)
--	WX3226 = NOT(WX3479)
--	WX3227 = NOT(WX3481)
--	WX3228 = NOT(WX3483)
--	WX3229 = NOT(WX3485)
--	WX3518 = NOT(WX3502)
--	WX3519 = NOT(WX3518)
--	WX3520 = NOT(WX3503)
--	WX3521 = NOT(WX3520)
--	WX3522 = NOT(WX3504)
--	WX3523 = NOT(WX3522)
--	WX3524 = NOT(WX3505)
--	WX3525 = NOT(WX3524)
--	WX3526 = NOT(WX3506)
--	WX3527 = NOT(WX3526)
--	WX3528 = NOT(WX3507)
--	WX3529 = NOT(WX3528)
--	WX3530 = NOT(WX3508)
--	WX3531 = NOT(WX3530)
--	WX3532 = NOT(WX3509)
--	WX3533 = NOT(WX3532)
--	WX3534 = NOT(WX3510)
--	WX3535 = NOT(WX3534)
--	WX3536 = NOT(WX3511)
--	WX3537 = NOT(WX3536)
--	WX3538 = NOT(WX3512)
--	WX3539 = NOT(WX3538)
--	WX3540 = NOT(WX3513)
--	WX3541 = NOT(WX3540)
--	WX3542 = NOT(WX3514)
--	WX3543 = NOT(WX3542)
--	WX3544 = NOT(WX3515)
--	WX3545 = NOT(WX3544)
--	WX3546 = NOT(WX3516)
--	WX3547 = NOT(WX3546)
--	WX3548 = NOT(WX3517)
--	WX3549 = NOT(WX3548)
--	WX3550 = NOT(WX3486)
--	WX3551 = NOT(WX3550)
--	WX3552 = NOT(WX3487)
--	WX3553 = NOT(WX3552)
--	WX3554 = NOT(WX3488)
--	WX3555 = NOT(WX3554)
--	WX3556 = NOT(WX3489)
--	WX3557 = NOT(WX3556)
--	WX3558 = NOT(WX3490)
--	WX3559 = NOT(WX3558)
--	WX3560 = NOT(WX3491)
--	WX3561 = NOT(WX3560)
--	WX3562 = NOT(WX3492)
--	WX3563 = NOT(WX3562)
--	WX3564 = NOT(WX3493)
--	WX3565 = NOT(WX3564)
--	WX3566 = NOT(WX3494)
--	WX3567 = NOT(WX3566)
--	WX3568 = NOT(WX3495)
--	WX3569 = NOT(WX3568)
--	WX3570 = NOT(WX3496)
--	WX3571 = NOT(WX3570)
--	WX3572 = NOT(WX3497)
--	WX3573 = NOT(WX3572)
--	WX3574 = NOT(WX3498)
--	WX3575 = NOT(WX3574)
--	WX3576 = NOT(WX3499)
--	WX3577 = NOT(WX3576)
--	WX3578 = NOT(WX3500)
--	WX3579 = NOT(WX3578)
--	WX3580 = NOT(WX3501)
--	WX3581 = NOT(WX3580)
--	WX3582 = NOT(TM0)
--	WX3583 = NOT(TM0)
--	WX3584 = NOT(TM0)
--	WX3585 = NOT(TM1)
--	WX3586 = NOT(TM1)
--	WX3587 = NOT(WX3586)
--	WX3588 = NOT(WX3584)
--	WX3589 = NOT(WX3585)
--	WX3590 = NOT(WX3583)
--	WX3591 = NOT(WX3582)
--	WX3595 = NOT(WX3591)
--	WX3597 = NOT(WX3596)
--	WX3598 = NOT(WX3597)
--	WX3602 = NOT(WX3591)
--	WX3604 = NOT(WX3603)
--	WX3605 = NOT(WX3604)
--	WX3609 = NOT(WX3591)
--	WX3611 = NOT(WX3610)
--	WX3612 = NOT(WX3611)
--	WX3616 = NOT(WX3591)
--	WX3618 = NOT(WX3617)
--	WX3619 = NOT(WX3618)
--	WX3623 = NOT(WX3591)
--	WX3625 = NOT(WX3624)
--	WX3626 = NOT(WX3625)
--	WX3630 = NOT(WX3591)
--	WX3632 = NOT(WX3631)
--	WX3633 = NOT(WX3632)
--	WX3637 = NOT(WX3591)
--	WX3639 = NOT(WX3638)
--	WX3640 = NOT(WX3639)
--	WX3644 = NOT(WX3591)
--	WX3646 = NOT(WX3645)
--	WX3647 = NOT(WX3646)
--	WX3651 = NOT(WX3591)
--	WX3653 = NOT(WX3652)
--	WX3654 = NOT(WX3653)
--	WX3658 = NOT(WX3591)
--	WX3660 = NOT(WX3659)
--	WX3661 = NOT(WX3660)
--	WX3665 = NOT(WX3591)
--	WX3667 = NOT(WX3666)
--	WX3668 = NOT(WX3667)
--	WX3672 = NOT(WX3591)
--	WX3674 = NOT(WX3673)
--	WX3675 = NOT(WX3674)
--	WX3679 = NOT(WX3591)
--	WX3681 = NOT(WX3680)
--	WX3682 = NOT(WX3681)
--	WX3686 = NOT(WX3591)
--	WX3688 = NOT(WX3687)
--	WX3689 = NOT(WX3688)
--	WX3693 = NOT(WX3591)
--	WX3695 = NOT(WX3694)
--	WX3696 = NOT(WX3695)
--	WX3700 = NOT(WX3591)
--	WX3702 = NOT(WX3701)
--	WX3703 = NOT(WX3702)
--	WX3707 = NOT(WX3591)
--	WX3709 = NOT(WX3708)
--	WX3710 = NOT(WX3709)
--	WX3714 = NOT(WX3591)
--	WX3716 = NOT(WX3715)
--	WX3717 = NOT(WX3716)
--	WX3721 = NOT(WX3591)
--	WX3723 = NOT(WX3722)
--	WX3724 = NOT(WX3723)
--	WX3728 = NOT(WX3591)
--	WX3730 = NOT(WX3729)
--	WX3731 = NOT(WX3730)
--	WX3735 = NOT(WX3591)
--	WX3737 = NOT(WX3736)
--	WX3738 = NOT(WX3737)
--	WX3742 = NOT(WX3591)
--	WX3744 = NOT(WX3743)
--	WX3745 = NOT(WX3744)
--	WX3749 = NOT(WX3591)
--	WX3751 = NOT(WX3750)
--	WX3752 = NOT(WX3751)
--	WX3756 = NOT(WX3591)
--	WX3758 = NOT(WX3757)
--	WX3759 = NOT(WX3758)
--	WX3763 = NOT(WX3591)
--	WX3765 = NOT(WX3764)
--	WX3766 = NOT(WX3765)
--	WX3770 = NOT(WX3591)
--	WX3772 = NOT(WX3771)
--	WX3773 = NOT(WX3772)
--	WX3777 = NOT(WX3591)
--	WX3779 = NOT(WX3778)
--	WX3780 = NOT(WX3779)
--	WX3784 = NOT(WX3591)
--	WX3786 = NOT(WX3785)
--	WX3787 = NOT(WX3786)
--	WX3791 = NOT(WX3591)
--	WX3793 = NOT(WX3792)
--	WX3794 = NOT(WX3793)
--	WX3798 = NOT(WX3591)
--	WX3800 = NOT(WX3799)
--	WX3801 = NOT(WX3800)
--	WX3805 = NOT(WX3591)
--	WX3807 = NOT(WX3806)
--	WX3808 = NOT(WX3807)
--	WX3812 = NOT(WX3591)
--	WX3814 = NOT(WX3813)
--	WX3815 = NOT(WX3814)
--	WX3816 = NOT(RESET)
--	WX3849 = NOT(WX3816)
--	WX3916 = NOT(WX4882)
--	WX3920 = NOT(WX4883)
--	WX3924 = NOT(WX4883)
--	WX3926 = NOT(WX3917)
--	WX3927 = NOT(WX3926)
--	WX3930 = NOT(WX4882)
--	WX3934 = NOT(WX4883)
--	WX3938 = NOT(WX4883)
--	WX3940 = NOT(WX3931)
--	WX3941 = NOT(WX3940)
--	WX3944 = NOT(WX4882)
--	WX3948 = NOT(WX4883)
--	WX3952 = NOT(WX4883)
--	WX3954 = NOT(WX3945)
--	WX3955 = NOT(WX3954)
--	WX3958 = NOT(WX4882)
--	WX3962 = NOT(WX4883)
--	WX3966 = NOT(WX4883)
--	WX3968 = NOT(WX3959)
--	WX3969 = NOT(WX3968)
--	WX3972 = NOT(WX4882)
--	WX3976 = NOT(WX4883)
--	WX3980 = NOT(WX4883)
--	WX3982 = NOT(WX3973)
--	WX3983 = NOT(WX3982)
--	WX3986 = NOT(WX4882)
--	WX3990 = NOT(WX4883)
--	WX3994 = NOT(WX4883)
--	WX3996 = NOT(WX3987)
--	WX3997 = NOT(WX3996)
--	WX4000 = NOT(WX4882)
--	WX4004 = NOT(WX4883)
--	WX4008 = NOT(WX4883)
--	WX4010 = NOT(WX4001)
--	WX4011 = NOT(WX4010)
--	WX4014 = NOT(WX4882)
--	WX4018 = NOT(WX4883)
--	WX4022 = NOT(WX4883)
--	WX4024 = NOT(WX4015)
--	WX4025 = NOT(WX4024)
--	WX4028 = NOT(WX4882)
--	WX4032 = NOT(WX4883)
--	WX4036 = NOT(WX4883)
--	WX4038 = NOT(WX4029)
--	WX4039 = NOT(WX4038)
--	WX4042 = NOT(WX4882)
--	WX4046 = NOT(WX4883)
--	WX4050 = NOT(WX4883)
--	WX4052 = NOT(WX4043)
--	WX4053 = NOT(WX4052)
--	WX4056 = NOT(WX4882)
--	WX4060 = NOT(WX4883)
--	WX4064 = NOT(WX4883)
--	WX4066 = NOT(WX4057)
--	WX4067 = NOT(WX4066)
--	WX4070 = NOT(WX4882)
--	WX4074 = NOT(WX4883)
--	WX4078 = NOT(WX4883)
--	WX4080 = NOT(WX4071)
--	WX4081 = NOT(WX4080)
--	WX4084 = NOT(WX4882)
--	WX4088 = NOT(WX4883)
--	WX4092 = NOT(WX4883)
--	WX4094 = NOT(WX4085)
--	WX4095 = NOT(WX4094)
--	WX4098 = NOT(WX4882)
--	WX4102 = NOT(WX4883)
--	WX4106 = NOT(WX4883)
--	WX4108 = NOT(WX4099)
--	WX4109 = NOT(WX4108)
--	WX4112 = NOT(WX4882)
--	WX4116 = NOT(WX4883)
--	WX4120 = NOT(WX4883)
--	WX4122 = NOT(WX4113)
--	WX4123 = NOT(WX4122)
--	WX4126 = NOT(WX4882)
--	WX4130 = NOT(WX4883)
--	WX4134 = NOT(WX4883)
--	WX4136 = NOT(WX4127)
--	WX4137 = NOT(WX4136)
--	WX4140 = NOT(WX4882)
--	WX4144 = NOT(WX4883)
--	WX4148 = NOT(WX4883)
--	WX4150 = NOT(WX4141)
--	WX4151 = NOT(WX4150)
--	WX4154 = NOT(WX4882)
--	WX4158 = NOT(WX4883)
--	WX4162 = NOT(WX4883)
--	WX4164 = NOT(WX4155)
--	WX4165 = NOT(WX4164)
--	WX4168 = NOT(WX4882)
--	WX4172 = NOT(WX4883)
--	WX4176 = NOT(WX4883)
--	WX4178 = NOT(WX4169)
--	WX4179 = NOT(WX4178)
--	WX4182 = NOT(WX4882)
--	WX4186 = NOT(WX4883)
--	WX4190 = NOT(WX4883)
--	WX4192 = NOT(WX4183)
--	WX4193 = NOT(WX4192)
--	WX4196 = NOT(WX4882)
--	WX4200 = NOT(WX4883)
--	WX4204 = NOT(WX4883)
--	WX4206 = NOT(WX4197)
--	WX4207 = NOT(WX4206)
--	WX4210 = NOT(WX4882)
--	WX4214 = NOT(WX4883)
--	WX4218 = NOT(WX4883)
--	WX4220 = NOT(WX4211)
--	WX4221 = NOT(WX4220)
--	WX4224 = NOT(WX4882)
--	WX4228 = NOT(WX4883)
--	WX4232 = NOT(WX4883)
--	WX4234 = NOT(WX4225)
--	WX4235 = NOT(WX4234)
--	WX4238 = NOT(WX4882)
--	WX4242 = NOT(WX4883)
--	WX4246 = NOT(WX4883)
--	WX4248 = NOT(WX4239)
--	WX4249 = NOT(WX4248)
--	WX4252 = NOT(WX4882)
--	WX4256 = NOT(WX4883)
--	WX4260 = NOT(WX4883)
--	WX4262 = NOT(WX4253)
--	WX4263 = NOT(WX4262)
--	WX4266 = NOT(WX4882)
--	WX4270 = NOT(WX4883)
--	WX4274 = NOT(WX4883)
--	WX4276 = NOT(WX4267)
--	WX4277 = NOT(WX4276)
--	WX4280 = NOT(WX4882)
--	WX4284 = NOT(WX4883)
--	WX4288 = NOT(WX4883)
--	WX4290 = NOT(WX4281)
--	WX4291 = NOT(WX4290)
--	WX4294 = NOT(WX4882)
--	WX4298 = NOT(WX4883)
--	WX4302 = NOT(WX4883)
--	WX4304 = NOT(WX4295)
--	WX4305 = NOT(WX4304)
--	WX4308 = NOT(WX4882)
--	WX4312 = NOT(WX4883)
--	WX4316 = NOT(WX4883)
--	WX4318 = NOT(WX4309)
--	WX4319 = NOT(WX4318)
--	WX4322 = NOT(WX4882)
--	WX4326 = NOT(WX4883)
--	WX4330 = NOT(WX4883)
--	WX4332 = NOT(WX4323)
--	WX4333 = NOT(WX4332)
--	WX4336 = NOT(WX4882)
--	WX4340 = NOT(WX4883)
--	WX4344 = NOT(WX4883)
--	WX4346 = NOT(WX4337)
--	WX4347 = NOT(WX4346)
--	WX4350 = NOT(WX4882)
--	WX4354 = NOT(WX4883)
--	WX4358 = NOT(WX4883)
--	WX4360 = NOT(WX4351)
--	WX4361 = NOT(WX4360)
--	WX4362 = NOT(WX4364)
--	WX4427 = NOT(WX4844)
--	WX4428 = NOT(WX4846)
--	WX4429 = NOT(WX4848)
--	WX4430 = NOT(WX4850)
--	WX4431 = NOT(WX4852)
--	WX4432 = NOT(WX4854)
--	WX4433 = NOT(WX4856)
--	WX4434 = NOT(WX4858)
--	WX4435 = NOT(WX4860)
--	WX4436 = NOT(WX4862)
--	WX4437 = NOT(WX4864)
--	WX4438 = NOT(WX4866)
--	WX4439 = NOT(WX4868)
--	WX4440 = NOT(WX4870)
--	WX4441 = NOT(WX4872)
--	WX4442 = NOT(WX4874)
--	WX4443 = NOT(WX4812)
--	WX4444 = NOT(WX4814)
--	WX4445 = NOT(WX4816)
--	WX4446 = NOT(WX4818)
--	WX4447 = NOT(WX4820)
--	WX4448 = NOT(WX4822)
--	WX4449 = NOT(WX4824)
--	WX4450 = NOT(WX4826)
--	WX4451 = NOT(WX4828)
--	WX4452 = NOT(WX4830)
--	WX4453 = NOT(WX4832)
--	WX4454 = NOT(WX4834)
--	WX4455 = NOT(WX4836)
--	WX4456 = NOT(WX4838)
--	WX4457 = NOT(WX4840)
--	WX4458 = NOT(WX4842)
--	WX4459 = NOT(WX4427)
--	WX4460 = NOT(WX4428)
--	WX4461 = NOT(WX4429)
--	WX4462 = NOT(WX4430)
--	WX4463 = NOT(WX4431)
--	WX4464 = NOT(WX4432)
--	WX4465 = NOT(WX4433)
--	WX4466 = NOT(WX4434)
--	WX4467 = NOT(WX4435)
--	WX4468 = NOT(WX4436)
--	WX4469 = NOT(WX4437)
--	WX4470 = NOT(WX4438)
--	WX4471 = NOT(WX4439)
--	WX4472 = NOT(WX4440)
--	WX4473 = NOT(WX4441)
--	WX4474 = NOT(WX4442)
--	WX4475 = NOT(WX4443)
--	WX4476 = NOT(WX4444)
--	WX4477 = NOT(WX4445)
--	WX4478 = NOT(WX4446)
--	WX4479 = NOT(WX4447)
--	WX4480 = NOT(WX4448)
--	WX4481 = NOT(WX4449)
--	WX4482 = NOT(WX4450)
--	WX4483 = NOT(WX4451)
--	WX4484 = NOT(WX4452)
--	WX4485 = NOT(WX4453)
--	WX4486 = NOT(WX4454)
--	WX4487 = NOT(WX4455)
--	WX4488 = NOT(WX4456)
--	WX4489 = NOT(WX4457)
--	WX4490 = NOT(WX4458)
--	WX4491 = NOT(WX4716)
--	WX4492 = NOT(WX4718)
--	WX4493 = NOT(WX4720)
--	WX4494 = NOT(WX4722)
--	WX4495 = NOT(WX4724)
--	WX4496 = NOT(WX4726)
--	WX4497 = NOT(WX4728)
--	WX4498 = NOT(WX4730)
--	WX4499 = NOT(WX4732)
--	WX4500 = NOT(WX4734)
--	WX4501 = NOT(WX4736)
--	WX4502 = NOT(WX4738)
--	WX4503 = NOT(WX4740)
--	WX4504 = NOT(WX4742)
--	WX4505 = NOT(WX4744)
--	WX4506 = NOT(WX4746)
--	WX4507 = NOT(WX4748)
--	WX4508 = NOT(WX4750)
--	WX4509 = NOT(WX4752)
--	WX4510 = NOT(WX4754)
--	WX4511 = NOT(WX4756)
--	WX4512 = NOT(WX4758)
--	WX4513 = NOT(WX4760)
--	WX4514 = NOT(WX4762)
--	WX4515 = NOT(WX4764)
--	WX4516 = NOT(WX4766)
--	WX4517 = NOT(WX4768)
--	WX4518 = NOT(WX4770)
--	WX4519 = NOT(WX4772)
--	WX4520 = NOT(WX4774)
--	WX4521 = NOT(WX4776)
--	WX4522 = NOT(WX4778)
--	WX4811 = NOT(WX4795)
--	WX4812 = NOT(WX4811)
--	WX4813 = NOT(WX4796)
--	WX4814 = NOT(WX4813)
--	WX4815 = NOT(WX4797)
--	WX4816 = NOT(WX4815)
--	WX4817 = NOT(WX4798)
--	WX4818 = NOT(WX4817)
--	WX4819 = NOT(WX4799)
--	WX4820 = NOT(WX4819)
--	WX4821 = NOT(WX4800)
--	WX4822 = NOT(WX4821)
--	WX4823 = NOT(WX4801)
--	WX4824 = NOT(WX4823)
--	WX4825 = NOT(WX4802)
--	WX4826 = NOT(WX4825)
--	WX4827 = NOT(WX4803)
--	WX4828 = NOT(WX4827)
--	WX4829 = NOT(WX4804)
--	WX4830 = NOT(WX4829)
--	WX4831 = NOT(WX4805)
--	WX4832 = NOT(WX4831)
--	WX4833 = NOT(WX4806)
--	WX4834 = NOT(WX4833)
--	WX4835 = NOT(WX4807)
--	WX4836 = NOT(WX4835)
--	WX4837 = NOT(WX4808)
--	WX4838 = NOT(WX4837)
--	WX4839 = NOT(WX4809)
--	WX4840 = NOT(WX4839)
--	WX4841 = NOT(WX4810)
--	WX4842 = NOT(WX4841)
--	WX4843 = NOT(WX4779)
--	WX4844 = NOT(WX4843)
--	WX4845 = NOT(WX4780)
--	WX4846 = NOT(WX4845)
--	WX4847 = NOT(WX4781)
--	WX4848 = NOT(WX4847)
--	WX4849 = NOT(WX4782)
--	WX4850 = NOT(WX4849)
--	WX4851 = NOT(WX4783)
--	WX4852 = NOT(WX4851)
--	WX4853 = NOT(WX4784)
--	WX4854 = NOT(WX4853)
--	WX4855 = NOT(WX4785)
--	WX4856 = NOT(WX4855)
--	WX4857 = NOT(WX4786)
--	WX4858 = NOT(WX4857)
--	WX4859 = NOT(WX4787)
--	WX4860 = NOT(WX4859)
--	WX4861 = NOT(WX4788)
--	WX4862 = NOT(WX4861)
--	WX4863 = NOT(WX4789)
--	WX4864 = NOT(WX4863)
--	WX4865 = NOT(WX4790)
--	WX4866 = NOT(WX4865)
--	WX4867 = NOT(WX4791)
--	WX4868 = NOT(WX4867)
--	WX4869 = NOT(WX4792)
--	WX4870 = NOT(WX4869)
--	WX4871 = NOT(WX4793)
--	WX4872 = NOT(WX4871)
--	WX4873 = NOT(WX4794)
--	WX4874 = NOT(WX4873)
--	WX4875 = NOT(TM0)
--	WX4876 = NOT(TM0)
--	WX4877 = NOT(TM0)
--	WX4878 = NOT(TM1)
--	WX4879 = NOT(TM1)
--	WX4880 = NOT(WX4879)
--	WX4881 = NOT(WX4877)
--	WX4882 = NOT(WX4878)
--	WX4883 = NOT(WX4876)
--	WX4884 = NOT(WX4875)
--	WX4888 = NOT(WX4884)
--	WX4890 = NOT(WX4889)
--	WX4891 = NOT(WX4890)
--	WX4895 = NOT(WX4884)
--	WX4897 = NOT(WX4896)
--	WX4898 = NOT(WX4897)
--	WX4902 = NOT(WX4884)
--	WX4904 = NOT(WX4903)
--	WX4905 = NOT(WX4904)
--	WX4909 = NOT(WX4884)
--	WX4911 = NOT(WX4910)
--	WX4912 = NOT(WX4911)
--	WX4916 = NOT(WX4884)
--	WX4918 = NOT(WX4917)
--	WX4919 = NOT(WX4918)
--	WX4923 = NOT(WX4884)
--	WX4925 = NOT(WX4924)
--	WX4926 = NOT(WX4925)
--	WX4930 = NOT(WX4884)
--	WX4932 = NOT(WX4931)
--	WX4933 = NOT(WX4932)
--	WX4937 = NOT(WX4884)
--	WX4939 = NOT(WX4938)
--	WX4940 = NOT(WX4939)
--	WX4944 = NOT(WX4884)
--	WX4946 = NOT(WX4945)
--	WX4947 = NOT(WX4946)
--	WX4951 = NOT(WX4884)
--	WX4953 = NOT(WX4952)
--	WX4954 = NOT(WX4953)
--	WX4958 = NOT(WX4884)
--	WX4960 = NOT(WX4959)
--	WX4961 = NOT(WX4960)
--	WX4965 = NOT(WX4884)
--	WX4967 = NOT(WX4966)
--	WX4968 = NOT(WX4967)
--	WX4972 = NOT(WX4884)
--	WX4974 = NOT(WX4973)
--	WX4975 = NOT(WX4974)
--	WX4979 = NOT(WX4884)
--	WX4981 = NOT(WX4980)
--	WX4982 = NOT(WX4981)
--	WX4986 = NOT(WX4884)
--	WX4988 = NOT(WX4987)
--	WX4989 = NOT(WX4988)
--	WX4993 = NOT(WX4884)
--	WX4995 = NOT(WX4994)
--	WX4996 = NOT(WX4995)
--	WX5000 = NOT(WX4884)
--	WX5002 = NOT(WX5001)
--	WX5003 = NOT(WX5002)
--	WX5007 = NOT(WX4884)
--	WX5009 = NOT(WX5008)
--	WX5010 = NOT(WX5009)
--	WX5014 = NOT(WX4884)
--	WX5016 = NOT(WX5015)
--	WX5017 = NOT(WX5016)
--	WX5021 = NOT(WX4884)
--	WX5023 = NOT(WX5022)
--	WX5024 = NOT(WX5023)
--	WX5028 = NOT(WX4884)
--	WX5030 = NOT(WX5029)
--	WX5031 = NOT(WX5030)
--	WX5035 = NOT(WX4884)
--	WX5037 = NOT(WX5036)
--	WX5038 = NOT(WX5037)
--	WX5042 = NOT(WX4884)
--	WX5044 = NOT(WX5043)
--	WX5045 = NOT(WX5044)
--	WX5049 = NOT(WX4884)
--	WX5051 = NOT(WX5050)
--	WX5052 = NOT(WX5051)
--	WX5056 = NOT(WX4884)
--	WX5058 = NOT(WX5057)
--	WX5059 = NOT(WX5058)
--	WX5063 = NOT(WX4884)
--	WX5065 = NOT(WX5064)
--	WX5066 = NOT(WX5065)
--	WX5070 = NOT(WX4884)
--	WX5072 = NOT(WX5071)
--	WX5073 = NOT(WX5072)
--	WX5077 = NOT(WX4884)
--	WX5079 = NOT(WX5078)
--	WX5080 = NOT(WX5079)
--	WX5084 = NOT(WX4884)
--	WX5086 = NOT(WX5085)
--	WX5087 = NOT(WX5086)
--	WX5091 = NOT(WX4884)
--	WX5093 = NOT(WX5092)
--	WX5094 = NOT(WX5093)
--	WX5098 = NOT(WX4884)
--	WX5100 = NOT(WX5099)
--	WX5101 = NOT(WX5100)
--	WX5105 = NOT(WX4884)
--	WX5107 = NOT(WX5106)
--	WX5108 = NOT(WX5107)
--	WX5109 = NOT(RESET)
--	WX5142 = NOT(WX5109)
--	WX5209 = NOT(WX6175)
--	WX5213 = NOT(WX6176)
--	WX5217 = NOT(WX6176)
--	WX5219 = NOT(WX5210)
--	WX5220 = NOT(WX5219)
--	WX5223 = NOT(WX6175)
--	WX5227 = NOT(WX6176)
--	WX5231 = NOT(WX6176)
--	WX5233 = NOT(WX5224)
--	WX5234 = NOT(WX5233)
--	WX5237 = NOT(WX6175)
--	WX5241 = NOT(WX6176)
--	WX5245 = NOT(WX6176)
--	WX5247 = NOT(WX5238)
--	WX5248 = NOT(WX5247)
--	WX5251 = NOT(WX6175)
--	WX5255 = NOT(WX6176)
--	WX5259 = NOT(WX6176)
--	WX5261 = NOT(WX5252)
--	WX5262 = NOT(WX5261)
--	WX5265 = NOT(WX6175)
--	WX5269 = NOT(WX6176)
--	WX5273 = NOT(WX6176)
--	WX5275 = NOT(WX5266)
--	WX5276 = NOT(WX5275)
--	WX5279 = NOT(WX6175)
--	WX5283 = NOT(WX6176)
--	WX5287 = NOT(WX6176)
--	WX5289 = NOT(WX5280)
--	WX5290 = NOT(WX5289)
--	WX5293 = NOT(WX6175)
--	WX5297 = NOT(WX6176)
--	WX5301 = NOT(WX6176)
--	WX5303 = NOT(WX5294)
--	WX5304 = NOT(WX5303)
--	WX5307 = NOT(WX6175)
--	WX5311 = NOT(WX6176)
--	WX5315 = NOT(WX6176)
--	WX5317 = NOT(WX5308)
--	WX5318 = NOT(WX5317)
--	WX5321 = NOT(WX6175)
--	WX5325 = NOT(WX6176)
--	WX5329 = NOT(WX6176)
--	WX5331 = NOT(WX5322)
--	WX5332 = NOT(WX5331)
--	WX5335 = NOT(WX6175)
--	WX5339 = NOT(WX6176)
--	WX5343 = NOT(WX6176)
--	WX5345 = NOT(WX5336)
--	WX5346 = NOT(WX5345)
--	WX5349 = NOT(WX6175)
--	WX5353 = NOT(WX6176)
--	WX5357 = NOT(WX6176)
--	WX5359 = NOT(WX5350)
--	WX5360 = NOT(WX5359)
--	WX5363 = NOT(WX6175)
--	WX5367 = NOT(WX6176)
--	WX5371 = NOT(WX6176)
--	WX5373 = NOT(WX5364)
--	WX5374 = NOT(WX5373)
--	WX5377 = NOT(WX6175)
--	WX5381 = NOT(WX6176)
--	WX5385 = NOT(WX6176)
--	WX5387 = NOT(WX5378)
--	WX5388 = NOT(WX5387)
--	WX5391 = NOT(WX6175)
--	WX5395 = NOT(WX6176)
--	WX5399 = NOT(WX6176)
--	WX5401 = NOT(WX5392)
--	WX5402 = NOT(WX5401)
--	WX5405 = NOT(WX6175)
--	WX5409 = NOT(WX6176)
--	WX5413 = NOT(WX6176)
--	WX5415 = NOT(WX5406)
--	WX5416 = NOT(WX5415)
--	WX5419 = NOT(WX6175)
--	WX5423 = NOT(WX6176)
--	WX5427 = NOT(WX6176)
--	WX5429 = NOT(WX5420)
--	WX5430 = NOT(WX5429)
--	WX5433 = NOT(WX6175)
--	WX5437 = NOT(WX6176)
--	WX5441 = NOT(WX6176)
--	WX5443 = NOT(WX5434)
--	WX5444 = NOT(WX5443)
--	WX5447 = NOT(WX6175)
--	WX5451 = NOT(WX6176)
--	WX5455 = NOT(WX6176)
--	WX5457 = NOT(WX5448)
--	WX5458 = NOT(WX5457)
--	WX5461 = NOT(WX6175)
--	WX5465 = NOT(WX6176)
--	WX5469 = NOT(WX6176)
--	WX5471 = NOT(WX5462)
--	WX5472 = NOT(WX5471)
--	WX5475 = NOT(WX6175)
--	WX5479 = NOT(WX6176)
--	WX5483 = NOT(WX6176)
--	WX5485 = NOT(WX5476)
--	WX5486 = NOT(WX5485)
--	WX5489 = NOT(WX6175)
--	WX5493 = NOT(WX6176)
--	WX5497 = NOT(WX6176)
--	WX5499 = NOT(WX5490)
--	WX5500 = NOT(WX5499)
--	WX5503 = NOT(WX6175)
--	WX5507 = NOT(WX6176)
--	WX5511 = NOT(WX6176)
--	WX5513 = NOT(WX5504)
--	WX5514 = NOT(WX5513)
--	WX5517 = NOT(WX6175)
--	WX5521 = NOT(WX6176)
--	WX5525 = NOT(WX6176)
--	WX5527 = NOT(WX5518)
--	WX5528 = NOT(WX5527)
--	WX5531 = NOT(WX6175)
--	WX5535 = NOT(WX6176)
--	WX5539 = NOT(WX6176)
--	WX5541 = NOT(WX5532)
--	WX5542 = NOT(WX5541)
--	WX5545 = NOT(WX6175)
--	WX5549 = NOT(WX6176)
--	WX5553 = NOT(WX6176)
--	WX5555 = NOT(WX5546)
--	WX5556 = NOT(WX5555)
--	WX5559 = NOT(WX6175)
--	WX5563 = NOT(WX6176)
--	WX5567 = NOT(WX6176)
--	WX5569 = NOT(WX5560)
--	WX5570 = NOT(WX5569)
--	WX5573 = NOT(WX6175)
--	WX5577 = NOT(WX6176)
--	WX5581 = NOT(WX6176)
--	WX5583 = NOT(WX5574)
--	WX5584 = NOT(WX5583)
--	WX5587 = NOT(WX6175)
--	WX5591 = NOT(WX6176)
--	WX5595 = NOT(WX6176)
--	WX5597 = NOT(WX5588)
--	WX5598 = NOT(WX5597)
--	WX5601 = NOT(WX6175)
--	WX5605 = NOT(WX6176)
--	WX5609 = NOT(WX6176)
--	WX5611 = NOT(WX5602)
--	WX5612 = NOT(WX5611)
--	WX5615 = NOT(WX6175)
--	WX5619 = NOT(WX6176)
--	WX5623 = NOT(WX6176)
--	WX5625 = NOT(WX5616)
--	WX5626 = NOT(WX5625)
--	WX5629 = NOT(WX6175)
--	WX5633 = NOT(WX6176)
--	WX5637 = NOT(WX6176)
--	WX5639 = NOT(WX5630)
--	WX5640 = NOT(WX5639)
--	WX5643 = NOT(WX6175)
--	WX5647 = NOT(WX6176)
--	WX5651 = NOT(WX6176)
--	WX5653 = NOT(WX5644)
--	WX5654 = NOT(WX5653)
--	WX5655 = NOT(WX5657)
--	WX5720 = NOT(WX6137)
--	WX5721 = NOT(WX6139)
--	WX5722 = NOT(WX6141)
--	WX5723 = NOT(WX6143)
--	WX5724 = NOT(WX6145)
--	WX5725 = NOT(WX6147)
--	WX5726 = NOT(WX6149)
--	WX5727 = NOT(WX6151)
--	WX5728 = NOT(WX6153)
--	WX5729 = NOT(WX6155)
--	WX5730 = NOT(WX6157)
--	WX5731 = NOT(WX6159)
--	WX5732 = NOT(WX6161)
--	WX5733 = NOT(WX6163)
--	WX5734 = NOT(WX6165)
--	WX5735 = NOT(WX6167)
--	WX5736 = NOT(WX6105)
--	WX5737 = NOT(WX6107)
--	WX5738 = NOT(WX6109)
--	WX5739 = NOT(WX6111)
--	WX5740 = NOT(WX6113)
--	WX5741 = NOT(WX6115)
--	WX5742 = NOT(WX6117)
--	WX5743 = NOT(WX6119)
--	WX5744 = NOT(WX6121)
--	WX5745 = NOT(WX6123)
--	WX5746 = NOT(WX6125)
--	WX5747 = NOT(WX6127)
--	WX5748 = NOT(WX6129)
--	WX5749 = NOT(WX6131)
--	WX5750 = NOT(WX6133)
--	WX5751 = NOT(WX6135)
--	WX5752 = NOT(WX5720)
--	WX5753 = NOT(WX5721)
--	WX5754 = NOT(WX5722)
--	WX5755 = NOT(WX5723)
--	WX5756 = NOT(WX5724)
--	WX5757 = NOT(WX5725)
--	WX5758 = NOT(WX5726)
--	WX5759 = NOT(WX5727)
--	WX5760 = NOT(WX5728)
--	WX5761 = NOT(WX5729)
--	WX5762 = NOT(WX5730)
--	WX5763 = NOT(WX5731)
--	WX5764 = NOT(WX5732)
--	WX5765 = NOT(WX5733)
--	WX5766 = NOT(WX5734)
--	WX5767 = NOT(WX5735)
--	WX5768 = NOT(WX5736)
--	WX5769 = NOT(WX5737)
--	WX5770 = NOT(WX5738)
--	WX5771 = NOT(WX5739)
--	WX5772 = NOT(WX5740)
--	WX5773 = NOT(WX5741)
--	WX5774 = NOT(WX5742)
--	WX5775 = NOT(WX5743)
--	WX5776 = NOT(WX5744)
--	WX5777 = NOT(WX5745)
--	WX5778 = NOT(WX5746)
--	WX5779 = NOT(WX5747)
--	WX5780 = NOT(WX5748)
--	WX5781 = NOT(WX5749)
--	WX5782 = NOT(WX5750)
--	WX5783 = NOT(WX5751)
--	WX5784 = NOT(WX6009)
--	WX5785 = NOT(WX6011)
--	WX5786 = NOT(WX6013)
--	WX5787 = NOT(WX6015)
--	WX5788 = NOT(WX6017)
--	WX5789 = NOT(WX6019)
--	WX5790 = NOT(WX6021)
--	WX5791 = NOT(WX6023)
--	WX5792 = NOT(WX6025)
--	WX5793 = NOT(WX6027)
--	WX5794 = NOT(WX6029)
--	WX5795 = NOT(WX6031)
--	WX5796 = NOT(WX6033)
--	WX5797 = NOT(WX6035)
--	WX5798 = NOT(WX6037)
--	WX5799 = NOT(WX6039)
--	WX5800 = NOT(WX6041)
--	WX5801 = NOT(WX6043)
--	WX5802 = NOT(WX6045)
--	WX5803 = NOT(WX6047)
--	WX5804 = NOT(WX6049)
--	WX5805 = NOT(WX6051)
--	WX5806 = NOT(WX6053)
--	WX5807 = NOT(WX6055)
--	WX5808 = NOT(WX6057)
--	WX5809 = NOT(WX6059)
--	WX5810 = NOT(WX6061)
--	WX5811 = NOT(WX6063)
--	WX5812 = NOT(WX6065)
--	WX5813 = NOT(WX6067)
--	WX5814 = NOT(WX6069)
--	WX5815 = NOT(WX6071)
--	WX6104 = NOT(WX6088)
--	WX6105 = NOT(WX6104)
--	WX6106 = NOT(WX6089)
--	WX6107 = NOT(WX6106)
--	WX6108 = NOT(WX6090)
--	WX6109 = NOT(WX6108)
--	WX6110 = NOT(WX6091)
--	WX6111 = NOT(WX6110)
--	WX6112 = NOT(WX6092)
--	WX6113 = NOT(WX6112)
--	WX6114 = NOT(WX6093)
--	WX6115 = NOT(WX6114)
--	WX6116 = NOT(WX6094)
--	WX6117 = NOT(WX6116)
--	WX6118 = NOT(WX6095)
--	WX6119 = NOT(WX6118)
--	WX6120 = NOT(WX6096)
--	WX6121 = NOT(WX6120)
--	WX6122 = NOT(WX6097)
--	WX6123 = NOT(WX6122)
--	WX6124 = NOT(WX6098)
--	WX6125 = NOT(WX6124)
--	WX6126 = NOT(WX6099)
--	WX6127 = NOT(WX6126)
--	WX6128 = NOT(WX6100)
--	WX6129 = NOT(WX6128)
--	WX6130 = NOT(WX6101)
--	WX6131 = NOT(WX6130)
--	WX6132 = NOT(WX6102)
--	WX6133 = NOT(WX6132)
--	WX6134 = NOT(WX6103)
--	WX6135 = NOT(WX6134)
--	WX6136 = NOT(WX6072)
--	WX6137 = NOT(WX6136)
--	WX6138 = NOT(WX6073)
--	WX6139 = NOT(WX6138)
--	WX6140 = NOT(WX6074)
--	WX6141 = NOT(WX6140)
--	WX6142 = NOT(WX6075)
--	WX6143 = NOT(WX6142)
--	WX6144 = NOT(WX6076)
--	WX6145 = NOT(WX6144)
--	WX6146 = NOT(WX6077)
--	WX6147 = NOT(WX6146)
--	WX6148 = NOT(WX6078)
--	WX6149 = NOT(WX6148)
--	WX6150 = NOT(WX6079)
--	WX6151 = NOT(WX6150)
--	WX6152 = NOT(WX6080)
--	WX6153 = NOT(WX6152)
--	WX6154 = NOT(WX6081)
--	WX6155 = NOT(WX6154)
--	WX6156 = NOT(WX6082)
--	WX6157 = NOT(WX6156)
--	WX6158 = NOT(WX6083)
--	WX6159 = NOT(WX6158)
--	WX6160 = NOT(WX6084)
--	WX6161 = NOT(WX6160)
--	WX6162 = NOT(WX6085)
--	WX6163 = NOT(WX6162)
--	WX6164 = NOT(WX6086)
--	WX6165 = NOT(WX6164)
--	WX6166 = NOT(WX6087)
--	WX6167 = NOT(WX6166)
--	WX6168 = NOT(TM0)
--	WX6169 = NOT(TM0)
--	WX6170 = NOT(TM0)
--	WX6171 = NOT(TM1)
--	WX6172 = NOT(TM1)
--	WX6173 = NOT(WX6172)
--	WX6174 = NOT(WX6170)
--	WX6175 = NOT(WX6171)
--	WX6176 = NOT(WX6169)
--	WX6177 = NOT(WX6168)
--	WX6181 = NOT(WX6177)
--	WX6183 = NOT(WX6182)
--	WX6184 = NOT(WX6183)
--	WX6188 = NOT(WX6177)
--	WX6190 = NOT(WX6189)
--	WX6191 = NOT(WX6190)
--	WX6195 = NOT(WX6177)
--	WX6197 = NOT(WX6196)
--	WX6198 = NOT(WX6197)
--	WX6202 = NOT(WX6177)
--	WX6204 = NOT(WX6203)
--	WX6205 = NOT(WX6204)
--	WX6209 = NOT(WX6177)
--	WX6211 = NOT(WX6210)
--	WX6212 = NOT(WX6211)
--	WX6216 = NOT(WX6177)
--	WX6218 = NOT(WX6217)
--	WX6219 = NOT(WX6218)
--	WX6223 = NOT(WX6177)
--	WX6225 = NOT(WX6224)
--	WX6226 = NOT(WX6225)
--	WX6230 = NOT(WX6177)
--	WX6232 = NOT(WX6231)
--	WX6233 = NOT(WX6232)
--	WX6237 = NOT(WX6177)
--	WX6239 = NOT(WX6238)
--	WX6240 = NOT(WX6239)
--	WX6244 = NOT(WX6177)
--	WX6246 = NOT(WX6245)
--	WX6247 = NOT(WX6246)
--	WX6251 = NOT(WX6177)
--	WX6253 = NOT(WX6252)
--	WX6254 = NOT(WX6253)
--	WX6258 = NOT(WX6177)
--	WX6260 = NOT(WX6259)
--	WX6261 = NOT(WX6260)
--	WX6265 = NOT(WX6177)
--	WX6267 = NOT(WX6266)
--	WX6268 = NOT(WX6267)
--	WX6272 = NOT(WX6177)
--	WX6274 = NOT(WX6273)
--	WX6275 = NOT(WX6274)
--	WX6279 = NOT(WX6177)
--	WX6281 = NOT(WX6280)
--	WX6282 = NOT(WX6281)
--	WX6286 = NOT(WX6177)
--	WX6288 = NOT(WX6287)
--	WX6289 = NOT(WX6288)
--	WX6293 = NOT(WX6177)
--	WX6295 = NOT(WX6294)
--	WX6296 = NOT(WX6295)
--	WX6300 = NOT(WX6177)
--	WX6302 = NOT(WX6301)
--	WX6303 = NOT(WX6302)
--	WX6307 = NOT(WX6177)
--	WX6309 = NOT(WX6308)
--	WX6310 = NOT(WX6309)
--	WX6314 = NOT(WX6177)
--	WX6316 = NOT(WX6315)
--	WX6317 = NOT(WX6316)
--	WX6321 = NOT(WX6177)
--	WX6323 = NOT(WX6322)
--	WX6324 = NOT(WX6323)
--	WX6328 = NOT(WX6177)
--	WX6330 = NOT(WX6329)
--	WX6331 = NOT(WX6330)
--	WX6335 = NOT(WX6177)
--	WX6337 = NOT(WX6336)
--	WX6338 = NOT(WX6337)
--	WX6342 = NOT(WX6177)
--	WX6344 = NOT(WX6343)
--	WX6345 = NOT(WX6344)
--	WX6349 = NOT(WX6177)
--	WX6351 = NOT(WX6350)
--	WX6352 = NOT(WX6351)
--	WX6356 = NOT(WX6177)
--	WX6358 = NOT(WX6357)
--	WX6359 = NOT(WX6358)
--	WX6363 = NOT(WX6177)
--	WX6365 = NOT(WX6364)
--	WX6366 = NOT(WX6365)
--	WX6370 = NOT(WX6177)
--	WX6372 = NOT(WX6371)
--	WX6373 = NOT(WX6372)
--	WX6377 = NOT(WX6177)
--	WX6379 = NOT(WX6378)
--	WX6380 = NOT(WX6379)
--	WX6384 = NOT(WX6177)
--	WX6386 = NOT(WX6385)
--	WX6387 = NOT(WX6386)
--	WX6391 = NOT(WX6177)
--	WX6393 = NOT(WX6392)
--	WX6394 = NOT(WX6393)
--	WX6398 = NOT(WX6177)
--	WX6400 = NOT(WX6399)
--	WX6401 = NOT(WX6400)
--	WX6402 = NOT(RESET)
--	WX6435 = NOT(WX6402)
--	WX6502 = NOT(WX7468)
--	WX6506 = NOT(WX7469)
--	WX6510 = NOT(WX7469)
--	WX6512 = NOT(WX6503)
--	WX6513 = NOT(WX6512)
--	WX6516 = NOT(WX7468)
--	WX6520 = NOT(WX7469)
--	WX6524 = NOT(WX7469)
--	WX6526 = NOT(WX6517)
--	WX6527 = NOT(WX6526)
--	WX6530 = NOT(WX7468)
--	WX6534 = NOT(WX7469)
--	WX6538 = NOT(WX7469)
--	WX6540 = NOT(WX6531)
--	WX6541 = NOT(WX6540)
--	WX6544 = NOT(WX7468)
--	WX6548 = NOT(WX7469)
--	WX6552 = NOT(WX7469)
--	WX6554 = NOT(WX6545)
--	WX6555 = NOT(WX6554)
--	WX6558 = NOT(WX7468)
--	WX6562 = NOT(WX7469)
--	WX6566 = NOT(WX7469)
--	WX6568 = NOT(WX6559)
--	WX6569 = NOT(WX6568)
--	WX6572 = NOT(WX7468)
--	WX6576 = NOT(WX7469)
--	WX6580 = NOT(WX7469)
--	WX6582 = NOT(WX6573)
--	WX6583 = NOT(WX6582)
--	WX6586 = NOT(WX7468)
--	WX6590 = NOT(WX7469)
--	WX6594 = NOT(WX7469)
--	WX6596 = NOT(WX6587)
--	WX6597 = NOT(WX6596)
--	WX6600 = NOT(WX7468)
--	WX6604 = NOT(WX7469)
--	WX6608 = NOT(WX7469)
--	WX6610 = NOT(WX6601)
--	WX6611 = NOT(WX6610)
--	WX6614 = NOT(WX7468)
--	WX6618 = NOT(WX7469)
--	WX6622 = NOT(WX7469)
--	WX6624 = NOT(WX6615)
--	WX6625 = NOT(WX6624)
--	WX6628 = NOT(WX7468)
--	WX6632 = NOT(WX7469)
--	WX6636 = NOT(WX7469)
--	WX6638 = NOT(WX6629)
--	WX6639 = NOT(WX6638)
--	WX6642 = NOT(WX7468)
--	WX6646 = NOT(WX7469)
--	WX6650 = NOT(WX7469)
--	WX6652 = NOT(WX6643)
--	WX6653 = NOT(WX6652)
--	WX6656 = NOT(WX7468)
--	WX6660 = NOT(WX7469)
--	WX6664 = NOT(WX7469)
--	WX6666 = NOT(WX6657)
--	WX6667 = NOT(WX6666)
--	WX6670 = NOT(WX7468)
--	WX6674 = NOT(WX7469)
--	WX6678 = NOT(WX7469)
--	WX6680 = NOT(WX6671)
--	WX6681 = NOT(WX6680)
--	WX6684 = NOT(WX7468)
--	WX6688 = NOT(WX7469)
--	WX6692 = NOT(WX7469)
--	WX6694 = NOT(WX6685)
--	WX6695 = NOT(WX6694)
--	WX6698 = NOT(WX7468)
--	WX6702 = NOT(WX7469)
--	WX6706 = NOT(WX7469)
--	WX6708 = NOT(WX6699)
--	WX6709 = NOT(WX6708)
--	WX6712 = NOT(WX7468)
--	WX6716 = NOT(WX7469)
--	WX6720 = NOT(WX7469)
--	WX6722 = NOT(WX6713)
--	WX6723 = NOT(WX6722)
--	WX6726 = NOT(WX7468)
--	WX6730 = NOT(WX7469)
--	WX6734 = NOT(WX7469)
--	WX6736 = NOT(WX6727)
--	WX6737 = NOT(WX6736)
--	WX6740 = NOT(WX7468)
--	WX6744 = NOT(WX7469)
--	WX6748 = NOT(WX7469)
--	WX6750 = NOT(WX6741)
--	WX6751 = NOT(WX6750)
--	WX6754 = NOT(WX7468)
--	WX6758 = NOT(WX7469)
--	WX6762 = NOT(WX7469)
--	WX6764 = NOT(WX6755)
--	WX6765 = NOT(WX6764)
--	WX6768 = NOT(WX7468)
--	WX6772 = NOT(WX7469)
--	WX6776 = NOT(WX7469)
--	WX6778 = NOT(WX6769)
--	WX6779 = NOT(WX6778)
--	WX6782 = NOT(WX7468)
--	WX6786 = NOT(WX7469)
--	WX6790 = NOT(WX7469)
--	WX6792 = NOT(WX6783)
--	WX6793 = NOT(WX6792)
--	WX6796 = NOT(WX7468)
--	WX6800 = NOT(WX7469)
--	WX6804 = NOT(WX7469)
--	WX6806 = NOT(WX6797)
--	WX6807 = NOT(WX6806)
--	WX6810 = NOT(WX7468)
--	WX6814 = NOT(WX7469)
--	WX6818 = NOT(WX7469)
--	WX6820 = NOT(WX6811)
--	WX6821 = NOT(WX6820)
--	WX6824 = NOT(WX7468)
--	WX6828 = NOT(WX7469)
--	WX6832 = NOT(WX7469)
--	WX6834 = NOT(WX6825)
--	WX6835 = NOT(WX6834)
--	WX6838 = NOT(WX7468)
--	WX6842 = NOT(WX7469)
--	WX6846 = NOT(WX7469)
--	WX6848 = NOT(WX6839)
--	WX6849 = NOT(WX6848)
--	WX6852 = NOT(WX7468)
--	WX6856 = NOT(WX7469)
--	WX6860 = NOT(WX7469)
--	WX6862 = NOT(WX6853)
--	WX6863 = NOT(WX6862)
--	WX6866 = NOT(WX7468)
--	WX6870 = NOT(WX7469)
--	WX6874 = NOT(WX7469)
--	WX6876 = NOT(WX6867)
--	WX6877 = NOT(WX6876)
--	WX6880 = NOT(WX7468)
--	WX6884 = NOT(WX7469)
--	WX6888 = NOT(WX7469)
--	WX6890 = NOT(WX6881)
--	WX6891 = NOT(WX6890)
--	WX6894 = NOT(WX7468)
--	WX6898 = NOT(WX7469)
--	WX6902 = NOT(WX7469)
--	WX6904 = NOT(WX6895)
--	WX6905 = NOT(WX6904)
--	WX6908 = NOT(WX7468)
--	WX6912 = NOT(WX7469)
--	WX6916 = NOT(WX7469)
--	WX6918 = NOT(WX6909)
--	WX6919 = NOT(WX6918)
--	WX6922 = NOT(WX7468)
--	WX6926 = NOT(WX7469)
--	WX6930 = NOT(WX7469)
--	WX6932 = NOT(WX6923)
--	WX6933 = NOT(WX6932)
--	WX6936 = NOT(WX7468)
--	WX6940 = NOT(WX7469)
--	WX6944 = NOT(WX7469)
--	WX6946 = NOT(WX6937)
--	WX6947 = NOT(WX6946)
--	WX6948 = NOT(WX6950)
--	WX7013 = NOT(WX7430)
--	WX7014 = NOT(WX7432)
--	WX7015 = NOT(WX7434)
--	WX7016 = NOT(WX7436)
--	WX7017 = NOT(WX7438)
--	WX7018 = NOT(WX7440)
--	WX7019 = NOT(WX7442)
--	WX7020 = NOT(WX7444)
--	WX7021 = NOT(WX7446)
--	WX7022 = NOT(WX7448)
--	WX7023 = NOT(WX7450)
--	WX7024 = NOT(WX7452)
--	WX7025 = NOT(WX7454)
--	WX7026 = NOT(WX7456)
--	WX7027 = NOT(WX7458)
--	WX7028 = NOT(WX7460)
--	WX7029 = NOT(WX7398)
--	WX7030 = NOT(WX7400)
--	WX7031 = NOT(WX7402)
--	WX7032 = NOT(WX7404)
--	WX7033 = NOT(WX7406)
--	WX7034 = NOT(WX7408)
--	WX7035 = NOT(WX7410)
--	WX7036 = NOT(WX7412)
--	WX7037 = NOT(WX7414)
--	WX7038 = NOT(WX7416)
--	WX7039 = NOT(WX7418)
--	WX7040 = NOT(WX7420)
--	WX7041 = NOT(WX7422)
--	WX7042 = NOT(WX7424)
--	WX7043 = NOT(WX7426)
--	WX7044 = NOT(WX7428)
--	WX7045 = NOT(WX7013)
--	WX7046 = NOT(WX7014)
--	WX7047 = NOT(WX7015)
--	WX7048 = NOT(WX7016)
--	WX7049 = NOT(WX7017)
--	WX7050 = NOT(WX7018)
--	WX7051 = NOT(WX7019)
--	WX7052 = NOT(WX7020)
--	WX7053 = NOT(WX7021)
--	WX7054 = NOT(WX7022)
--	WX7055 = NOT(WX7023)
--	WX7056 = NOT(WX7024)
--	WX7057 = NOT(WX7025)
--	WX7058 = NOT(WX7026)
--	WX7059 = NOT(WX7027)
--	WX7060 = NOT(WX7028)
--	WX7061 = NOT(WX7029)
--	WX7062 = NOT(WX7030)
--	WX7063 = NOT(WX7031)
--	WX7064 = NOT(WX7032)
--	WX7065 = NOT(WX7033)
--	WX7066 = NOT(WX7034)
--	WX7067 = NOT(WX7035)
--	WX7068 = NOT(WX7036)
--	WX7069 = NOT(WX7037)
--	WX7070 = NOT(WX7038)
--	WX7071 = NOT(WX7039)
--	WX7072 = NOT(WX7040)
--	WX7073 = NOT(WX7041)
--	WX7074 = NOT(WX7042)
--	WX7075 = NOT(WX7043)
--	WX7076 = NOT(WX7044)
--	WX7077 = NOT(WX7302)
--	WX7078 = NOT(WX7304)
--	WX7079 = NOT(WX7306)
--	WX7080 = NOT(WX7308)
--	WX7081 = NOT(WX7310)
--	WX7082 = NOT(WX7312)
--	WX7083 = NOT(WX7314)
--	WX7084 = NOT(WX7316)
--	WX7085 = NOT(WX7318)
--	WX7086 = NOT(WX7320)
--	WX7087 = NOT(WX7322)
--	WX7088 = NOT(WX7324)
--	WX7089 = NOT(WX7326)
--	WX7090 = NOT(WX7328)
--	WX7091 = NOT(WX7330)
--	WX7092 = NOT(WX7332)
--	WX7093 = NOT(WX7334)
--	WX7094 = NOT(WX7336)
--	WX7095 = NOT(WX7338)
--	WX7096 = NOT(WX7340)
--	WX7097 = NOT(WX7342)
--	WX7098 = NOT(WX7344)
--	WX7099 = NOT(WX7346)
--	WX7100 = NOT(WX7348)
--	WX7101 = NOT(WX7350)
--	WX7102 = NOT(WX7352)
--	WX7103 = NOT(WX7354)
--	WX7104 = NOT(WX7356)
--	WX7105 = NOT(WX7358)
--	WX7106 = NOT(WX7360)
--	WX7107 = NOT(WX7362)
--	WX7108 = NOT(WX7364)
--	WX7397 = NOT(WX7381)
--	WX7398 = NOT(WX7397)
--	WX7399 = NOT(WX7382)
--	WX7400 = NOT(WX7399)
--	WX7401 = NOT(WX7383)
--	WX7402 = NOT(WX7401)
--	WX7403 = NOT(WX7384)
--	WX7404 = NOT(WX7403)
--	WX7405 = NOT(WX7385)
--	WX7406 = NOT(WX7405)
--	WX7407 = NOT(WX7386)
--	WX7408 = NOT(WX7407)
--	WX7409 = NOT(WX7387)
--	WX7410 = NOT(WX7409)
--	WX7411 = NOT(WX7388)
--	WX7412 = NOT(WX7411)
--	WX7413 = NOT(WX7389)
--	WX7414 = NOT(WX7413)
--	WX7415 = NOT(WX7390)
--	WX7416 = NOT(WX7415)
--	WX7417 = NOT(WX7391)
--	WX7418 = NOT(WX7417)
--	WX7419 = NOT(WX7392)
--	WX7420 = NOT(WX7419)
--	WX7421 = NOT(WX7393)
--	WX7422 = NOT(WX7421)
--	WX7423 = NOT(WX7394)
--	WX7424 = NOT(WX7423)
--	WX7425 = NOT(WX7395)
--	WX7426 = NOT(WX7425)
--	WX7427 = NOT(WX7396)
--	WX7428 = NOT(WX7427)
--	WX7429 = NOT(WX7365)
--	WX7430 = NOT(WX7429)
--	WX7431 = NOT(WX7366)
--	WX7432 = NOT(WX7431)
--	WX7433 = NOT(WX7367)
--	WX7434 = NOT(WX7433)
--	WX7435 = NOT(WX7368)
--	WX7436 = NOT(WX7435)
--	WX7437 = NOT(WX7369)
--	WX7438 = NOT(WX7437)
--	WX7439 = NOT(WX7370)
--	WX7440 = NOT(WX7439)
--	WX7441 = NOT(WX7371)
--	WX7442 = NOT(WX7441)
--	WX7443 = NOT(WX7372)
--	WX7444 = NOT(WX7443)
--	WX7445 = NOT(WX7373)
--	WX7446 = NOT(WX7445)
--	WX7447 = NOT(WX7374)
--	WX7448 = NOT(WX7447)
--	WX7449 = NOT(WX7375)
--	WX7450 = NOT(WX7449)
--	WX7451 = NOT(WX7376)
--	WX7452 = NOT(WX7451)
--	WX7453 = NOT(WX7377)
--	WX7454 = NOT(WX7453)
--	WX7455 = NOT(WX7378)
--	WX7456 = NOT(WX7455)
--	WX7457 = NOT(WX7379)
--	WX7458 = NOT(WX7457)
--	WX7459 = NOT(WX7380)
--	WX7460 = NOT(WX7459)
--	WX7461 = NOT(TM0)
--	WX7462 = NOT(TM0)
--	WX7463 = NOT(TM0)
--	WX7464 = NOT(TM1)
--	WX7465 = NOT(TM1)
--	WX7466 = NOT(WX7465)
--	WX7467 = NOT(WX7463)
--	WX7468 = NOT(WX7464)
--	WX7469 = NOT(WX7462)
--	WX7470 = NOT(WX7461)
--	WX7474 = NOT(WX7470)
--	WX7476 = NOT(WX7475)
--	WX7477 = NOT(WX7476)
--	WX7481 = NOT(WX7470)
--	WX7483 = NOT(WX7482)
--	WX7484 = NOT(WX7483)
--	WX7488 = NOT(WX7470)
--	WX7490 = NOT(WX7489)
--	WX7491 = NOT(WX7490)
--	WX7495 = NOT(WX7470)
--	WX7497 = NOT(WX7496)
--	WX7498 = NOT(WX7497)
--	WX7502 = NOT(WX7470)
--	WX7504 = NOT(WX7503)
--	WX7505 = NOT(WX7504)
--	WX7509 = NOT(WX7470)
--	WX7511 = NOT(WX7510)
--	WX7512 = NOT(WX7511)
--	WX7516 = NOT(WX7470)
--	WX7518 = NOT(WX7517)
--	WX7519 = NOT(WX7518)
--	WX7523 = NOT(WX7470)
--	WX7525 = NOT(WX7524)
--	WX7526 = NOT(WX7525)
--	WX7530 = NOT(WX7470)
--	WX7532 = NOT(WX7531)
--	WX7533 = NOT(WX7532)
--	WX7537 = NOT(WX7470)
--	WX7539 = NOT(WX7538)
--	WX7540 = NOT(WX7539)
--	WX7544 = NOT(WX7470)
--	WX7546 = NOT(WX7545)
--	WX7547 = NOT(WX7546)
--	WX7551 = NOT(WX7470)
--	WX7553 = NOT(WX7552)
--	WX7554 = NOT(WX7553)
--	WX7558 = NOT(WX7470)
--	WX7560 = NOT(WX7559)
--	WX7561 = NOT(WX7560)
--	WX7565 = NOT(WX7470)
--	WX7567 = NOT(WX7566)
--	WX7568 = NOT(WX7567)
--	WX7572 = NOT(WX7470)
--	WX7574 = NOT(WX7573)
--	WX7575 = NOT(WX7574)
--	WX7579 = NOT(WX7470)
--	WX7581 = NOT(WX7580)
--	WX7582 = NOT(WX7581)
--	WX7586 = NOT(WX7470)
--	WX7588 = NOT(WX7587)
--	WX7589 = NOT(WX7588)
--	WX7593 = NOT(WX7470)
--	WX7595 = NOT(WX7594)
--	WX7596 = NOT(WX7595)
--	WX7600 = NOT(WX7470)
--	WX7602 = NOT(WX7601)
--	WX7603 = NOT(WX7602)
--	WX7607 = NOT(WX7470)
--	WX7609 = NOT(WX7608)
--	WX7610 = NOT(WX7609)
--	WX7614 = NOT(WX7470)
--	WX7616 = NOT(WX7615)
--	WX7617 = NOT(WX7616)
--	WX7621 = NOT(WX7470)
--	WX7623 = NOT(WX7622)
--	WX7624 = NOT(WX7623)
--	WX7628 = NOT(WX7470)
--	WX7630 = NOT(WX7629)
--	WX7631 = NOT(WX7630)
--	WX7635 = NOT(WX7470)
--	WX7637 = NOT(WX7636)
--	WX7638 = NOT(WX7637)
--	WX7642 = NOT(WX7470)
--	WX7644 = NOT(WX7643)
--	WX7645 = NOT(WX7644)
--	WX7649 = NOT(WX7470)
--	WX7651 = NOT(WX7650)
--	WX7652 = NOT(WX7651)
--	WX7656 = NOT(WX7470)
--	WX7658 = NOT(WX7657)
--	WX7659 = NOT(WX7658)
--	WX7663 = NOT(WX7470)
--	WX7665 = NOT(WX7664)
--	WX7666 = NOT(WX7665)
--	WX7670 = NOT(WX7470)
--	WX7672 = NOT(WX7671)
--	WX7673 = NOT(WX7672)
--	WX7677 = NOT(WX7470)
--	WX7679 = NOT(WX7678)
--	WX7680 = NOT(WX7679)
--	WX7684 = NOT(WX7470)
--	WX7686 = NOT(WX7685)
--	WX7687 = NOT(WX7686)
--	WX7691 = NOT(WX7470)
--	WX7693 = NOT(WX7692)
--	WX7694 = NOT(WX7693)
--	WX7695 = NOT(RESET)
--	WX7728 = NOT(WX7695)
--	WX7795 = NOT(WX8761)
--	WX7799 = NOT(WX8762)
--	WX7803 = NOT(WX8762)
--	WX7805 = NOT(WX7796)
--	WX7806 = NOT(WX7805)
--	WX7809 = NOT(WX8761)
--	WX7813 = NOT(WX8762)
--	WX7817 = NOT(WX8762)
--	WX7819 = NOT(WX7810)
--	WX7820 = NOT(WX7819)
--	WX7823 = NOT(WX8761)
--	WX7827 = NOT(WX8762)
--	WX7831 = NOT(WX8762)
--	WX7833 = NOT(WX7824)
--	WX7834 = NOT(WX7833)
--	WX7837 = NOT(WX8761)
--	WX7841 = NOT(WX8762)
--	WX7845 = NOT(WX8762)
--	WX7847 = NOT(WX7838)
--	WX7848 = NOT(WX7847)
--	WX7851 = NOT(WX8761)
--	WX7855 = NOT(WX8762)
--	WX7859 = NOT(WX8762)
--	WX7861 = NOT(WX7852)
--	WX7862 = NOT(WX7861)
--	WX7865 = NOT(WX8761)
--	WX7869 = NOT(WX8762)
--	WX7873 = NOT(WX8762)
--	WX7875 = NOT(WX7866)
--	WX7876 = NOT(WX7875)
--	WX7879 = NOT(WX8761)
--	WX7883 = NOT(WX8762)
--	WX7887 = NOT(WX8762)
--	WX7889 = NOT(WX7880)
--	WX7890 = NOT(WX7889)
--	WX7893 = NOT(WX8761)
--	WX7897 = NOT(WX8762)
--	WX7901 = NOT(WX8762)
--	WX7903 = NOT(WX7894)
--	WX7904 = NOT(WX7903)
--	WX7907 = NOT(WX8761)
--	WX7911 = NOT(WX8762)
--	WX7915 = NOT(WX8762)
--	WX7917 = NOT(WX7908)
--	WX7918 = NOT(WX7917)
--	WX7921 = NOT(WX8761)
--	WX7925 = NOT(WX8762)
--	WX7929 = NOT(WX8762)
--	WX7931 = NOT(WX7922)
--	WX7932 = NOT(WX7931)
--	WX7935 = NOT(WX8761)
--	WX7939 = NOT(WX8762)
--	WX7943 = NOT(WX8762)
--	WX7945 = NOT(WX7936)
--	WX7946 = NOT(WX7945)
--	WX7949 = NOT(WX8761)
--	WX7953 = NOT(WX8762)
--	WX7957 = NOT(WX8762)
--	WX7959 = NOT(WX7950)
--	WX7960 = NOT(WX7959)
--	WX7963 = NOT(WX8761)
--	WX7967 = NOT(WX8762)
--	WX7971 = NOT(WX8762)
--	WX7973 = NOT(WX7964)
--	WX7974 = NOT(WX7973)
--	WX7977 = NOT(WX8761)
--	WX7981 = NOT(WX8762)
--	WX7985 = NOT(WX8762)
--	WX7987 = NOT(WX7978)
--	WX7988 = NOT(WX7987)
--	WX7991 = NOT(WX8761)
--	WX7995 = NOT(WX8762)
--	WX7999 = NOT(WX8762)
--	WX8001 = NOT(WX7992)
--	WX8002 = NOT(WX8001)
--	WX8005 = NOT(WX8761)
--	WX8009 = NOT(WX8762)
--	WX8013 = NOT(WX8762)
--	WX8015 = NOT(WX8006)
--	WX8016 = NOT(WX8015)
--	WX8019 = NOT(WX8761)
--	WX8023 = NOT(WX8762)
--	WX8027 = NOT(WX8762)
--	WX8029 = NOT(WX8020)
--	WX8030 = NOT(WX8029)
--	WX8033 = NOT(WX8761)
--	WX8037 = NOT(WX8762)
--	WX8041 = NOT(WX8762)
--	WX8043 = NOT(WX8034)
--	WX8044 = NOT(WX8043)
--	WX8047 = NOT(WX8761)
--	WX8051 = NOT(WX8762)
--	WX8055 = NOT(WX8762)
--	WX8057 = NOT(WX8048)
--	WX8058 = NOT(WX8057)
--	WX8061 = NOT(WX8761)
--	WX8065 = NOT(WX8762)
--	WX8069 = NOT(WX8762)
--	WX8071 = NOT(WX8062)
--	WX8072 = NOT(WX8071)
--	WX8075 = NOT(WX8761)
--	WX8079 = NOT(WX8762)
--	WX8083 = NOT(WX8762)
--	WX8085 = NOT(WX8076)
--	WX8086 = NOT(WX8085)
--	WX8089 = NOT(WX8761)
--	WX8093 = NOT(WX8762)
--	WX8097 = NOT(WX8762)
--	WX8099 = NOT(WX8090)
--	WX8100 = NOT(WX8099)
--	WX8103 = NOT(WX8761)
--	WX8107 = NOT(WX8762)
--	WX8111 = NOT(WX8762)
--	WX8113 = NOT(WX8104)
--	WX8114 = NOT(WX8113)
--	WX8117 = NOT(WX8761)
--	WX8121 = NOT(WX8762)
--	WX8125 = NOT(WX8762)
--	WX8127 = NOT(WX8118)
--	WX8128 = NOT(WX8127)
--	WX8131 = NOT(WX8761)
--	WX8135 = NOT(WX8762)
--	WX8139 = NOT(WX8762)
--	WX8141 = NOT(WX8132)
--	WX8142 = NOT(WX8141)
--	WX8145 = NOT(WX8761)
--	WX8149 = NOT(WX8762)
--	WX8153 = NOT(WX8762)
--	WX8155 = NOT(WX8146)
--	WX8156 = NOT(WX8155)
--	WX8159 = NOT(WX8761)
--	WX8163 = NOT(WX8762)
--	WX8167 = NOT(WX8762)
--	WX8169 = NOT(WX8160)
--	WX8170 = NOT(WX8169)
--	WX8173 = NOT(WX8761)
--	WX8177 = NOT(WX8762)
--	WX8181 = NOT(WX8762)
--	WX8183 = NOT(WX8174)
--	WX8184 = NOT(WX8183)
--	WX8187 = NOT(WX8761)
--	WX8191 = NOT(WX8762)
--	WX8195 = NOT(WX8762)
--	WX8197 = NOT(WX8188)
--	WX8198 = NOT(WX8197)
--	WX8201 = NOT(WX8761)
--	WX8205 = NOT(WX8762)
--	WX8209 = NOT(WX8762)
--	WX8211 = NOT(WX8202)
--	WX8212 = NOT(WX8211)
--	WX8215 = NOT(WX8761)
--	WX8219 = NOT(WX8762)
--	WX8223 = NOT(WX8762)
--	WX8225 = NOT(WX8216)
--	WX8226 = NOT(WX8225)
--	WX8229 = NOT(WX8761)
--	WX8233 = NOT(WX8762)
--	WX8237 = NOT(WX8762)
--	WX8239 = NOT(WX8230)
--	WX8240 = NOT(WX8239)
--	WX8241 = NOT(WX8243)
--	WX8306 = NOT(WX8723)
--	WX8307 = NOT(WX8725)
--	WX8308 = NOT(WX8727)
--	WX8309 = NOT(WX8729)
--	WX8310 = NOT(WX8731)
--	WX8311 = NOT(WX8733)
--	WX8312 = NOT(WX8735)
--	WX8313 = NOT(WX8737)
--	WX8314 = NOT(WX8739)
--	WX8315 = NOT(WX8741)
--	WX8316 = NOT(WX8743)
--	WX8317 = NOT(WX8745)
--	WX8318 = NOT(WX8747)
--	WX8319 = NOT(WX8749)
--	WX8320 = NOT(WX8751)
--	WX8321 = NOT(WX8753)
--	WX8322 = NOT(WX8691)
--	WX8323 = NOT(WX8693)
--	WX8324 = NOT(WX8695)
--	WX8325 = NOT(WX8697)
--	WX8326 = NOT(WX8699)
--	WX8327 = NOT(WX8701)
--	WX8328 = NOT(WX8703)
--	WX8329 = NOT(WX8705)
--	WX8330 = NOT(WX8707)
--	WX8331 = NOT(WX8709)
--	WX8332 = NOT(WX8711)
--	WX8333 = NOT(WX8713)
--	WX8334 = NOT(WX8715)
--	WX8335 = NOT(WX8717)
--	WX8336 = NOT(WX8719)
--	WX8337 = NOT(WX8721)
--	WX8338 = NOT(WX8306)
--	WX8339 = NOT(WX8307)
--	WX8340 = NOT(WX8308)
--	WX8341 = NOT(WX8309)
--	WX8342 = NOT(WX8310)
--	WX8343 = NOT(WX8311)
--	WX8344 = NOT(WX8312)
--	WX8345 = NOT(WX8313)
--	WX8346 = NOT(WX8314)
--	WX8347 = NOT(WX8315)
--	WX8348 = NOT(WX8316)
--	WX8349 = NOT(WX8317)
--	WX8350 = NOT(WX8318)
--	WX8351 = NOT(WX8319)
--	WX8352 = NOT(WX8320)
--	WX8353 = NOT(WX8321)
--	WX8354 = NOT(WX8322)
--	WX8355 = NOT(WX8323)
--	WX8356 = NOT(WX8324)
--	WX8357 = NOT(WX8325)
--	WX8358 = NOT(WX8326)
--	WX8359 = NOT(WX8327)
--	WX8360 = NOT(WX8328)
--	WX8361 = NOT(WX8329)
--	WX8362 = NOT(WX8330)
--	WX8363 = NOT(WX8331)
--	WX8364 = NOT(WX8332)
--	WX8365 = NOT(WX8333)
--	WX8366 = NOT(WX8334)
--	WX8367 = NOT(WX8335)
--	WX8368 = NOT(WX8336)
--	WX8369 = NOT(WX8337)
--	WX8370 = NOT(WX8595)
--	WX8371 = NOT(WX8597)
--	WX8372 = NOT(WX8599)
--	WX8373 = NOT(WX8601)
--	WX8374 = NOT(WX8603)
--	WX8375 = NOT(WX8605)
--	WX8376 = NOT(WX8607)
--	WX8377 = NOT(WX8609)
--	WX8378 = NOT(WX8611)
--	WX8379 = NOT(WX8613)
--	WX8380 = NOT(WX8615)
--	WX8381 = NOT(WX8617)
--	WX8382 = NOT(WX8619)
--	WX8383 = NOT(WX8621)
--	WX8384 = NOT(WX8623)
--	WX8385 = NOT(WX8625)
--	WX8386 = NOT(WX8627)
--	WX8387 = NOT(WX8629)
--	WX8388 = NOT(WX8631)
--	WX8389 = NOT(WX8633)
--	WX8390 = NOT(WX8635)
--	WX8391 = NOT(WX8637)
--	WX8392 = NOT(WX8639)
--	WX8393 = NOT(WX8641)
--	WX8394 = NOT(WX8643)
--	WX8395 = NOT(WX8645)
--	WX8396 = NOT(WX8647)
--	WX8397 = NOT(WX8649)
--	WX8398 = NOT(WX8651)
--	WX8399 = NOT(WX8653)
--	WX8400 = NOT(WX8655)
--	WX8401 = NOT(WX8657)
--	WX8690 = NOT(WX8674)
--	WX8691 = NOT(WX8690)
--	WX8692 = NOT(WX8675)
--	WX8693 = NOT(WX8692)
--	WX8694 = NOT(WX8676)
--	WX8695 = NOT(WX8694)
--	WX8696 = NOT(WX8677)
--	WX8697 = NOT(WX8696)
--	WX8698 = NOT(WX8678)
--	WX8699 = NOT(WX8698)
--	WX8700 = NOT(WX8679)
--	WX8701 = NOT(WX8700)
--	WX8702 = NOT(WX8680)
--	WX8703 = NOT(WX8702)
--	WX8704 = NOT(WX8681)
--	WX8705 = NOT(WX8704)
--	WX8706 = NOT(WX8682)
--	WX8707 = NOT(WX8706)
--	WX8708 = NOT(WX8683)
--	WX8709 = NOT(WX8708)
--	WX8710 = NOT(WX8684)
--	WX8711 = NOT(WX8710)
--	WX8712 = NOT(WX8685)
--	WX8713 = NOT(WX8712)
--	WX8714 = NOT(WX8686)
--	WX8715 = NOT(WX8714)
--	WX8716 = NOT(WX8687)
--	WX8717 = NOT(WX8716)
--	WX8718 = NOT(WX8688)
--	WX8719 = NOT(WX8718)
--	WX8720 = NOT(WX8689)
--	WX8721 = NOT(WX8720)
--	WX8722 = NOT(WX8658)
--	WX8723 = NOT(WX8722)
--	WX8724 = NOT(WX8659)
--	WX8725 = NOT(WX8724)
--	WX8726 = NOT(WX8660)
--	WX8727 = NOT(WX8726)
--	WX8728 = NOT(WX8661)
--	WX8729 = NOT(WX8728)
--	WX8730 = NOT(WX8662)
--	WX8731 = NOT(WX8730)
--	WX8732 = NOT(WX8663)
--	WX8733 = NOT(WX8732)
--	WX8734 = NOT(WX8664)
--	WX8735 = NOT(WX8734)
--	WX8736 = NOT(WX8665)
--	WX8737 = NOT(WX8736)
--	WX8738 = NOT(WX8666)
--	WX8739 = NOT(WX8738)
--	WX8740 = NOT(WX8667)
--	WX8741 = NOT(WX8740)
--	WX8742 = NOT(WX8668)
--	WX8743 = NOT(WX8742)
--	WX8744 = NOT(WX8669)
--	WX8745 = NOT(WX8744)
--	WX8746 = NOT(WX8670)
--	WX8747 = NOT(WX8746)
--	WX8748 = NOT(WX8671)
--	WX8749 = NOT(WX8748)
--	WX8750 = NOT(WX8672)
--	WX8751 = NOT(WX8750)
--	WX8752 = NOT(WX8673)
--	WX8753 = NOT(WX8752)
--	WX8754 = NOT(TM0)
--	WX8755 = NOT(TM0)
--	WX8756 = NOT(TM0)
--	WX8757 = NOT(TM1)
--	WX8758 = NOT(TM1)
--	WX8759 = NOT(WX8758)
--	WX8760 = NOT(WX8756)
--	WX8761 = NOT(WX8757)
--	WX8762 = NOT(WX8755)
--	WX8763 = NOT(WX8754)
--	WX8767 = NOT(WX8763)
--	WX8769 = NOT(WX8768)
--	WX8770 = NOT(WX8769)
--	WX8774 = NOT(WX8763)
--	WX8776 = NOT(WX8775)
--	WX8777 = NOT(WX8776)
--	WX8781 = NOT(WX8763)
--	WX8783 = NOT(WX8782)
--	WX8784 = NOT(WX8783)
--	WX8788 = NOT(WX8763)
--	WX8790 = NOT(WX8789)
--	WX8791 = NOT(WX8790)
--	WX8795 = NOT(WX8763)
--	WX8797 = NOT(WX8796)
--	WX8798 = NOT(WX8797)
--	WX8802 = NOT(WX8763)
--	WX8804 = NOT(WX8803)
--	WX8805 = NOT(WX8804)
--	WX8809 = NOT(WX8763)
--	WX8811 = NOT(WX8810)
--	WX8812 = NOT(WX8811)
--	WX8816 = NOT(WX8763)
--	WX8818 = NOT(WX8817)
--	WX8819 = NOT(WX8818)
--	WX8823 = NOT(WX8763)
--	WX8825 = NOT(WX8824)
--	WX8826 = NOT(WX8825)
--	WX8830 = NOT(WX8763)
--	WX8832 = NOT(WX8831)
--	WX8833 = NOT(WX8832)
--	WX8837 = NOT(WX8763)
--	WX8839 = NOT(WX8838)
--	WX8840 = NOT(WX8839)
--	WX8844 = NOT(WX8763)
--	WX8846 = NOT(WX8845)
--	WX8847 = NOT(WX8846)
--	WX8851 = NOT(WX8763)
--	WX8853 = NOT(WX8852)
--	WX8854 = NOT(WX8853)
--	WX8858 = NOT(WX8763)
--	WX8860 = NOT(WX8859)
--	WX8861 = NOT(WX8860)
--	WX8865 = NOT(WX8763)
--	WX8867 = NOT(WX8866)
--	WX8868 = NOT(WX8867)
--	WX8872 = NOT(WX8763)
--	WX8874 = NOT(WX8873)
--	WX8875 = NOT(WX8874)
--	WX8879 = NOT(WX8763)
--	WX8881 = NOT(WX8880)
--	WX8882 = NOT(WX8881)
--	WX8886 = NOT(WX8763)
--	WX8888 = NOT(WX8887)
--	WX8889 = NOT(WX8888)
--	WX8893 = NOT(WX8763)
--	WX8895 = NOT(WX8894)
--	WX8896 = NOT(WX8895)
--	WX8900 = NOT(WX8763)
--	WX8902 = NOT(WX8901)
--	WX8903 = NOT(WX8902)
--	WX8907 = NOT(WX8763)
--	WX8909 = NOT(WX8908)
--	WX8910 = NOT(WX8909)
--	WX8914 = NOT(WX8763)
--	WX8916 = NOT(WX8915)
--	WX8917 = NOT(WX8916)
--	WX8921 = NOT(WX8763)
--	WX8923 = NOT(WX8922)
--	WX8924 = NOT(WX8923)
--	WX8928 = NOT(WX8763)
--	WX8930 = NOT(WX8929)
--	WX8931 = NOT(WX8930)
--	WX8935 = NOT(WX8763)
--	WX8937 = NOT(WX8936)
--	WX8938 = NOT(WX8937)
--	WX8942 = NOT(WX8763)
--	WX8944 = NOT(WX8943)
--	WX8945 = NOT(WX8944)
--	WX8949 = NOT(WX8763)
--	WX8951 = NOT(WX8950)
--	WX8952 = NOT(WX8951)
--	WX8956 = NOT(WX8763)
--	WX8958 = NOT(WX8957)
--	WX8959 = NOT(WX8958)
--	WX8963 = NOT(WX8763)
--	WX8965 = NOT(WX8964)
--	WX8966 = NOT(WX8965)
--	WX8970 = NOT(WX8763)
--	WX8972 = NOT(WX8971)
--	WX8973 = NOT(WX8972)
--	WX8977 = NOT(WX8763)
--	WX8979 = NOT(WX8978)
--	WX8980 = NOT(WX8979)
--	WX8984 = NOT(WX8763)
--	WX8986 = NOT(WX8985)
--	WX8987 = NOT(WX8986)
--	WX8988 = NOT(RESET)
--	WX9021 = NOT(WX8988)
--	WX9088 = NOT(WX10054)
--	WX9092 = NOT(WX10055)
--	WX9096 = NOT(WX10055)
--	WX9098 = NOT(WX9089)
--	WX9099 = NOT(WX9098)
--	WX9102 = NOT(WX10054)
--	WX9106 = NOT(WX10055)
--	WX9110 = NOT(WX10055)
--	WX9112 = NOT(WX9103)
--	WX9113 = NOT(WX9112)
--	WX9116 = NOT(WX10054)
--	WX9120 = NOT(WX10055)
--	WX9124 = NOT(WX10055)
--	WX9126 = NOT(WX9117)
--	WX9127 = NOT(WX9126)
--	WX9130 = NOT(WX10054)
--	WX9134 = NOT(WX10055)
--	WX9138 = NOT(WX10055)
--	WX9140 = NOT(WX9131)
--	WX9141 = NOT(WX9140)
--	WX9144 = NOT(WX10054)
--	WX9148 = NOT(WX10055)
--	WX9152 = NOT(WX10055)
--	WX9154 = NOT(WX9145)
--	WX9155 = NOT(WX9154)
--	WX9158 = NOT(WX10054)
--	WX9162 = NOT(WX10055)
--	WX9166 = NOT(WX10055)
--	WX9168 = NOT(WX9159)
--	WX9169 = NOT(WX9168)
--	WX9172 = NOT(WX10054)
--	WX9176 = NOT(WX10055)
--	WX9180 = NOT(WX10055)
--	WX9182 = NOT(WX9173)
--	WX9183 = NOT(WX9182)
--	WX9186 = NOT(WX10054)
--	WX9190 = NOT(WX10055)
--	WX9194 = NOT(WX10055)
--	WX9196 = NOT(WX9187)
--	WX9197 = NOT(WX9196)
--	WX9200 = NOT(WX10054)
--	WX9204 = NOT(WX10055)
--	WX9208 = NOT(WX10055)
--	WX9210 = NOT(WX9201)
--	WX9211 = NOT(WX9210)
--	WX9214 = NOT(WX10054)
--	WX9218 = NOT(WX10055)
--	WX9222 = NOT(WX10055)
--	WX9224 = NOT(WX9215)
--	WX9225 = NOT(WX9224)
--	WX9228 = NOT(WX10054)
--	WX9232 = NOT(WX10055)
--	WX9236 = NOT(WX10055)
--	WX9238 = NOT(WX9229)
--	WX9239 = NOT(WX9238)
--	WX9242 = NOT(WX10054)
--	WX9246 = NOT(WX10055)
--	WX9250 = NOT(WX10055)
--	WX9252 = NOT(WX9243)
--	WX9253 = NOT(WX9252)
--	WX9256 = NOT(WX10054)
--	WX9260 = NOT(WX10055)
--	WX9264 = NOT(WX10055)
--	WX9266 = NOT(WX9257)
--	WX9267 = NOT(WX9266)
--	WX9270 = NOT(WX10054)
--	WX9274 = NOT(WX10055)
--	WX9278 = NOT(WX10055)
--	WX9280 = NOT(WX9271)
--	WX9281 = NOT(WX9280)
--	WX9284 = NOT(WX10054)
--	WX9288 = NOT(WX10055)
--	WX9292 = NOT(WX10055)
--	WX9294 = NOT(WX9285)
--	WX9295 = NOT(WX9294)
--	WX9298 = NOT(WX10054)
--	WX9302 = NOT(WX10055)
--	WX9306 = NOT(WX10055)
--	WX9308 = NOT(WX9299)
--	WX9309 = NOT(WX9308)
--	WX9312 = NOT(WX10054)
--	WX9316 = NOT(WX10055)
--	WX9320 = NOT(WX10055)
--	WX9322 = NOT(WX9313)
--	WX9323 = NOT(WX9322)
--	WX9326 = NOT(WX10054)
--	WX9330 = NOT(WX10055)
--	WX9334 = NOT(WX10055)
--	WX9336 = NOT(WX9327)
--	WX9337 = NOT(WX9336)
--	WX9340 = NOT(WX10054)
--	WX9344 = NOT(WX10055)
--	WX9348 = NOT(WX10055)
--	WX9350 = NOT(WX9341)
--	WX9351 = NOT(WX9350)
--	WX9354 = NOT(WX10054)
--	WX9358 = NOT(WX10055)
--	WX9362 = NOT(WX10055)
--	WX9364 = NOT(WX9355)
--	WX9365 = NOT(WX9364)
--	WX9368 = NOT(WX10054)
--	WX9372 = NOT(WX10055)
--	WX9376 = NOT(WX10055)
--	WX9378 = NOT(WX9369)
--	WX9379 = NOT(WX9378)
--	WX9382 = NOT(WX10054)
--	WX9386 = NOT(WX10055)
--	WX9390 = NOT(WX10055)
--	WX9392 = NOT(WX9383)
--	WX9393 = NOT(WX9392)
--	WX9396 = NOT(WX10054)
--	WX9400 = NOT(WX10055)
--	WX9404 = NOT(WX10055)
--	WX9406 = NOT(WX9397)
--	WX9407 = NOT(WX9406)
--	WX9410 = NOT(WX10054)
--	WX9414 = NOT(WX10055)
--	WX9418 = NOT(WX10055)
--	WX9420 = NOT(WX9411)
--	WX9421 = NOT(WX9420)
--	WX9424 = NOT(WX10054)
--	WX9428 = NOT(WX10055)
--	WX9432 = NOT(WX10055)
--	WX9434 = NOT(WX9425)
--	WX9435 = NOT(WX9434)
--	WX9438 = NOT(WX10054)
--	WX9442 = NOT(WX10055)
--	WX9446 = NOT(WX10055)
--	WX9448 = NOT(WX9439)
--	WX9449 = NOT(WX9448)
--	WX9452 = NOT(WX10054)
--	WX9456 = NOT(WX10055)
--	WX9460 = NOT(WX10055)
--	WX9462 = NOT(WX9453)
--	WX9463 = NOT(WX9462)
--	WX9466 = NOT(WX10054)
--	WX9470 = NOT(WX10055)
--	WX9474 = NOT(WX10055)
--	WX9476 = NOT(WX9467)
--	WX9477 = NOT(WX9476)
--	WX9480 = NOT(WX10054)
--	WX9484 = NOT(WX10055)
--	WX9488 = NOT(WX10055)
--	WX9490 = NOT(WX9481)
--	WX9491 = NOT(WX9490)
--	WX9494 = NOT(WX10054)
--	WX9498 = NOT(WX10055)
--	WX9502 = NOT(WX10055)
--	WX9504 = NOT(WX9495)
--	WX9505 = NOT(WX9504)
--	WX9508 = NOT(WX10054)
--	WX9512 = NOT(WX10055)
--	WX9516 = NOT(WX10055)
--	WX9518 = NOT(WX9509)
--	WX9519 = NOT(WX9518)
--	WX9522 = NOT(WX10054)
--	WX9526 = NOT(WX10055)
--	WX9530 = NOT(WX10055)
--	WX9532 = NOT(WX9523)
--	WX9533 = NOT(WX9532)
--	WX9534 = NOT(WX9536)
--	WX9599 = NOT(WX10016)
--	WX9600 = NOT(WX10018)
--	WX9601 = NOT(WX10020)
--	WX9602 = NOT(WX10022)
--	WX9603 = NOT(WX10024)
--	WX9604 = NOT(WX10026)
--	WX9605 = NOT(WX10028)
--	WX9606 = NOT(WX10030)
--	WX9607 = NOT(WX10032)
--	WX9608 = NOT(WX10034)
--	WX9609 = NOT(WX10036)
--	WX9610 = NOT(WX10038)
--	WX9611 = NOT(WX10040)
--	WX9612 = NOT(WX10042)
--	WX9613 = NOT(WX10044)
--	WX9614 = NOT(WX10046)
--	WX9615 = NOT(WX9984)
--	WX9616 = NOT(WX9986)
--	WX9617 = NOT(WX9988)
--	WX9618 = NOT(WX9990)
--	WX9619 = NOT(WX9992)
--	WX9620 = NOT(WX9994)
--	WX9621 = NOT(WX9996)
--	WX9622 = NOT(WX9998)
--	WX9623 = NOT(WX10000)
--	WX9624 = NOT(WX10002)
--	WX9625 = NOT(WX10004)
--	WX9626 = NOT(WX10006)
--	WX9627 = NOT(WX10008)
--	WX9628 = NOT(WX10010)
--	WX9629 = NOT(WX10012)
--	WX9630 = NOT(WX10014)
--	WX9631 = NOT(WX9599)
--	WX9632 = NOT(WX9600)
--	WX9633 = NOT(WX9601)
--	WX9634 = NOT(WX9602)
--	WX9635 = NOT(WX9603)
--	WX9636 = NOT(WX9604)
--	WX9637 = NOT(WX9605)
--	WX9638 = NOT(WX9606)
--	WX9639 = NOT(WX9607)
--	WX9640 = NOT(WX9608)
--	WX9641 = NOT(WX9609)
--	WX9642 = NOT(WX9610)
--	WX9643 = NOT(WX9611)
--	WX9644 = NOT(WX9612)
--	WX9645 = NOT(WX9613)
--	WX9646 = NOT(WX9614)
--	WX9647 = NOT(WX9615)
--	WX9648 = NOT(WX9616)
--	WX9649 = NOT(WX9617)
--	WX9650 = NOT(WX9618)
--	WX9651 = NOT(WX9619)
--	WX9652 = NOT(WX9620)
--	WX9653 = NOT(WX9621)
--	WX9654 = NOT(WX9622)
--	WX9655 = NOT(WX9623)
--	WX9656 = NOT(WX9624)
--	WX9657 = NOT(WX9625)
--	WX9658 = NOT(WX9626)
--	WX9659 = NOT(WX9627)
--	WX9660 = NOT(WX9628)
--	WX9661 = NOT(WX9629)
--	WX9662 = NOT(WX9630)
--	WX9663 = NOT(WX9888)
--	WX9664 = NOT(WX9890)
--	WX9665 = NOT(WX9892)
--	WX9666 = NOT(WX9894)
--	WX9667 = NOT(WX9896)
--	WX9668 = NOT(WX9898)
--	WX9669 = NOT(WX9900)
--	WX9670 = NOT(WX9902)
--	WX9671 = NOT(WX9904)
--	WX9672 = NOT(WX9906)
--	WX9673 = NOT(WX9908)
--	WX9674 = NOT(WX9910)
--	WX9675 = NOT(WX9912)
--	WX9676 = NOT(WX9914)
--	WX9677 = NOT(WX9916)
--	WX9678 = NOT(WX9918)
--	WX9679 = NOT(WX9920)
--	WX9680 = NOT(WX9922)
--	WX9681 = NOT(WX9924)
--	WX9682 = NOT(WX9926)
--	WX9683 = NOT(WX9928)
--	WX9684 = NOT(WX9930)
--	WX9685 = NOT(WX9932)
--	WX9686 = NOT(WX9934)
--	WX9687 = NOT(WX9936)
--	WX9688 = NOT(WX9938)
--	WX9689 = NOT(WX9940)
--	WX9690 = NOT(WX9942)
--	WX9691 = NOT(WX9944)
--	WX9692 = NOT(WX9946)
--	WX9693 = NOT(WX9948)
--	WX9694 = NOT(WX9950)
--	WX9983 = NOT(WX9967)
--	WX9984 = NOT(WX9983)
--	WX9985 = NOT(WX9968)
--	WX9986 = NOT(WX9985)
--	WX9987 = NOT(WX9969)
--	WX9988 = NOT(WX9987)
--	WX9989 = NOT(WX9970)
--	WX9990 = NOT(WX9989)
--	WX9991 = NOT(WX9971)
--	WX9992 = NOT(WX9991)
--	WX9993 = NOT(WX9972)
--	WX9994 = NOT(WX9993)
--	WX9995 = NOT(WX9973)
--	WX9996 = NOT(WX9995)
--	WX9997 = NOT(WX9974)
--	WX9998 = NOT(WX9997)
--	WX9999 = NOT(WX9975)
--	WX10000 = NOT(WX9999)
--	WX10001 = NOT(WX9976)
--	WX10002 = NOT(WX10001)
--	WX10003 = NOT(WX9977)
--	WX10004 = NOT(WX10003)
--	WX10005 = NOT(WX9978)
--	WX10006 = NOT(WX10005)
--	WX10007 = NOT(WX9979)
--	WX10008 = NOT(WX10007)
--	WX10009 = NOT(WX9980)
--	WX10010 = NOT(WX10009)
--	WX10011 = NOT(WX9981)
--	WX10012 = NOT(WX10011)
--	WX10013 = NOT(WX9982)
--	WX10014 = NOT(WX10013)
--	WX10015 = NOT(WX9951)
--	WX10016 = NOT(WX10015)
--	WX10017 = NOT(WX9952)
--	WX10018 = NOT(WX10017)
--	WX10019 = NOT(WX9953)
--	WX10020 = NOT(WX10019)
--	WX10021 = NOT(WX9954)
--	WX10022 = NOT(WX10021)
--	WX10023 = NOT(WX9955)
--	WX10024 = NOT(WX10023)
--	WX10025 = NOT(WX9956)
--	WX10026 = NOT(WX10025)
--	WX10027 = NOT(WX9957)
--	WX10028 = NOT(WX10027)
--	WX10029 = NOT(WX9958)
--	WX10030 = NOT(WX10029)
--	WX10031 = NOT(WX9959)
--	WX10032 = NOT(WX10031)
--	WX10033 = NOT(WX9960)
--	WX10034 = NOT(WX10033)
--	WX10035 = NOT(WX9961)
--	WX10036 = NOT(WX10035)
--	WX10037 = NOT(WX9962)
--	WX10038 = NOT(WX10037)
--	WX10039 = NOT(WX9963)
--	WX10040 = NOT(WX10039)
--	WX10041 = NOT(WX9964)
--	WX10042 = NOT(WX10041)
--	WX10043 = NOT(WX9965)
--	WX10044 = NOT(WX10043)
--	WX10045 = NOT(WX9966)
--	WX10046 = NOT(WX10045)
--	WX10047 = NOT(TM0)
--	WX10048 = NOT(TM0)
--	WX10049 = NOT(TM0)
--	WX10050 = NOT(TM1)
--	WX10051 = NOT(TM1)
--	WX10052 = NOT(WX10051)
--	WX10053 = NOT(WX10049)
--	WX10054 = NOT(WX10050)
--	WX10055 = NOT(WX10048)
--	WX10056 = NOT(WX10047)
--	WX10060 = NOT(WX10056)
--	WX10062 = NOT(WX10061)
--	WX10063 = NOT(WX10062)
--	WX10067 = NOT(WX10056)
--	WX10069 = NOT(WX10068)
--	WX10070 = NOT(WX10069)
--	WX10074 = NOT(WX10056)
--	WX10076 = NOT(WX10075)
--	WX10077 = NOT(WX10076)
--	WX10081 = NOT(WX10056)
--	WX10083 = NOT(WX10082)
--	WX10084 = NOT(WX10083)
--	WX10088 = NOT(WX10056)
--	WX10090 = NOT(WX10089)
--	WX10091 = NOT(WX10090)
--	WX10095 = NOT(WX10056)
--	WX10097 = NOT(WX10096)
--	WX10098 = NOT(WX10097)
--	WX10102 = NOT(WX10056)
--	WX10104 = NOT(WX10103)
--	WX10105 = NOT(WX10104)
--	WX10109 = NOT(WX10056)
--	WX10111 = NOT(WX10110)
--	WX10112 = NOT(WX10111)
--	WX10116 = NOT(WX10056)
--	WX10118 = NOT(WX10117)
--	WX10119 = NOT(WX10118)
--	WX10123 = NOT(WX10056)
--	WX10125 = NOT(WX10124)
--	WX10126 = NOT(WX10125)
--	WX10130 = NOT(WX10056)
--	WX10132 = NOT(WX10131)
--	WX10133 = NOT(WX10132)
--	WX10137 = NOT(WX10056)
--	WX10139 = NOT(WX10138)
--	WX10140 = NOT(WX10139)
--	WX10144 = NOT(WX10056)
--	WX10146 = NOT(WX10145)
--	WX10147 = NOT(WX10146)
--	WX10151 = NOT(WX10056)
--	WX10153 = NOT(WX10152)
--	WX10154 = NOT(WX10153)
--	WX10158 = NOT(WX10056)
--	WX10160 = NOT(WX10159)
--	WX10161 = NOT(WX10160)
--	WX10165 = NOT(WX10056)
--	WX10167 = NOT(WX10166)
--	WX10168 = NOT(WX10167)
--	WX10172 = NOT(WX10056)
--	WX10174 = NOT(WX10173)
--	WX10175 = NOT(WX10174)
--	WX10179 = NOT(WX10056)
--	WX10181 = NOT(WX10180)
--	WX10182 = NOT(WX10181)
--	WX10186 = NOT(WX10056)
--	WX10188 = NOT(WX10187)
--	WX10189 = NOT(WX10188)
--	WX10193 = NOT(WX10056)
--	WX10195 = NOT(WX10194)
--	WX10196 = NOT(WX10195)
--	WX10200 = NOT(WX10056)
--	WX10202 = NOT(WX10201)
--	WX10203 = NOT(WX10202)
--	WX10207 = NOT(WX10056)
--	WX10209 = NOT(WX10208)
--	WX10210 = NOT(WX10209)
--	WX10214 = NOT(WX10056)
--	WX10216 = NOT(WX10215)
--	WX10217 = NOT(WX10216)
--	WX10221 = NOT(WX10056)
--	WX10223 = NOT(WX10222)
--	WX10224 = NOT(WX10223)
--	WX10228 = NOT(WX10056)
--	WX10230 = NOT(WX10229)
--	WX10231 = NOT(WX10230)
--	WX10235 = NOT(WX10056)
--	WX10237 = NOT(WX10236)
--	WX10238 = NOT(WX10237)
--	WX10242 = NOT(WX10056)
--	WX10244 = NOT(WX10243)
--	WX10245 = NOT(WX10244)
--	WX10249 = NOT(WX10056)
--	WX10251 = NOT(WX10250)
--	WX10252 = NOT(WX10251)
--	WX10256 = NOT(WX10056)
--	WX10258 = NOT(WX10257)
--	WX10259 = NOT(WX10258)
--	WX10263 = NOT(WX10056)
--	WX10265 = NOT(WX10264)
--	WX10266 = NOT(WX10265)
--	WX10270 = NOT(WX10056)
--	WX10272 = NOT(WX10271)
--	WX10273 = NOT(WX10272)
--	WX10277 = NOT(WX10056)
--	WX10279 = NOT(WX10278)
--	WX10280 = NOT(WX10279)
--	WX10281 = NOT(RESET)
--	WX10314 = NOT(WX10281)
--	WX10381 = NOT(WX11347)
--	WX10385 = NOT(WX11348)
--	WX10389 = NOT(WX11348)
--	WX10391 = NOT(WX10382)
--	WX10392 = NOT(WX10391)
--	WX10395 = NOT(WX11347)
--	WX10399 = NOT(WX11348)
--	WX10403 = NOT(WX11348)
--	WX10405 = NOT(WX10396)
--	WX10406 = NOT(WX10405)
--	WX10409 = NOT(WX11347)
--	WX10413 = NOT(WX11348)
--	WX10417 = NOT(WX11348)
--	WX10419 = NOT(WX10410)
--	WX10420 = NOT(WX10419)
--	WX10423 = NOT(WX11347)
--	WX10427 = NOT(WX11348)
--	WX10431 = NOT(WX11348)
--	WX10433 = NOT(WX10424)
--	WX10434 = NOT(WX10433)
--	WX10437 = NOT(WX11347)
--	WX10441 = NOT(WX11348)
--	WX10445 = NOT(WX11348)
--	WX10447 = NOT(WX10438)
--	WX10448 = NOT(WX10447)
--	WX10451 = NOT(WX11347)
--	WX10455 = NOT(WX11348)
--	WX10459 = NOT(WX11348)
--	WX10461 = NOT(WX10452)
--	WX10462 = NOT(WX10461)
--	WX10465 = NOT(WX11347)
--	WX10469 = NOT(WX11348)
--	WX10473 = NOT(WX11348)
--	WX10475 = NOT(WX10466)
--	WX10476 = NOT(WX10475)
--	WX10479 = NOT(WX11347)
--	WX10483 = NOT(WX11348)
--	WX10487 = NOT(WX11348)
--	WX10489 = NOT(WX10480)
--	WX10490 = NOT(WX10489)
--	WX10493 = NOT(WX11347)
--	WX10497 = NOT(WX11348)
--	WX10501 = NOT(WX11348)
--	WX10503 = NOT(WX10494)
--	WX10504 = NOT(WX10503)
--	WX10507 = NOT(WX11347)
--	WX10511 = NOT(WX11348)
--	WX10515 = NOT(WX11348)
--	WX10517 = NOT(WX10508)
--	WX10518 = NOT(WX10517)
--	WX10521 = NOT(WX11347)
--	WX10525 = NOT(WX11348)
--	WX10529 = NOT(WX11348)
--	WX10531 = NOT(WX10522)
--	WX10532 = NOT(WX10531)
--	WX10535 = NOT(WX11347)
--	WX10539 = NOT(WX11348)
--	WX10543 = NOT(WX11348)
--	WX10545 = NOT(WX10536)
--	WX10546 = NOT(WX10545)
--	WX10549 = NOT(WX11347)
--	WX10553 = NOT(WX11348)
--	WX10557 = NOT(WX11348)
--	WX10559 = NOT(WX10550)
--	WX10560 = NOT(WX10559)
--	WX10563 = NOT(WX11347)
--	WX10567 = NOT(WX11348)
--	WX10571 = NOT(WX11348)
--	WX10573 = NOT(WX10564)
--	WX10574 = NOT(WX10573)
--	WX10577 = NOT(WX11347)
--	WX10581 = NOT(WX11348)
--	WX10585 = NOT(WX11348)
--	WX10587 = NOT(WX10578)
--	WX10588 = NOT(WX10587)
--	WX10591 = NOT(WX11347)
--	WX10595 = NOT(WX11348)
--	WX10599 = NOT(WX11348)
--	WX10601 = NOT(WX10592)
--	WX10602 = NOT(WX10601)
--	WX10605 = NOT(WX11347)
--	WX10609 = NOT(WX11348)
--	WX10613 = NOT(WX11348)
--	WX10615 = NOT(WX10606)
--	WX10616 = NOT(WX10615)
--	WX10619 = NOT(WX11347)
--	WX10623 = NOT(WX11348)
--	WX10627 = NOT(WX11348)
--	WX10629 = NOT(WX10620)
--	WX10630 = NOT(WX10629)
--	WX10633 = NOT(WX11347)
--	WX10637 = NOT(WX11348)
--	WX10641 = NOT(WX11348)
--	WX10643 = NOT(WX10634)
--	WX10644 = NOT(WX10643)
--	WX10647 = NOT(WX11347)
--	WX10651 = NOT(WX11348)
--	WX10655 = NOT(WX11348)
--	WX10657 = NOT(WX10648)
--	WX10658 = NOT(WX10657)
--	WX10661 = NOT(WX11347)
--	WX10665 = NOT(WX11348)
--	WX10669 = NOT(WX11348)
--	WX10671 = NOT(WX10662)
--	WX10672 = NOT(WX10671)
--	WX10675 = NOT(WX11347)
--	WX10679 = NOT(WX11348)
--	WX10683 = NOT(WX11348)
--	WX10685 = NOT(WX10676)
--	WX10686 = NOT(WX10685)
--	WX10689 = NOT(WX11347)
--	WX10693 = NOT(WX11348)
--	WX10697 = NOT(WX11348)
--	WX10699 = NOT(WX10690)
--	WX10700 = NOT(WX10699)
--	WX10703 = NOT(WX11347)
--	WX10707 = NOT(WX11348)
--	WX10711 = NOT(WX11348)
--	WX10713 = NOT(WX10704)
--	WX10714 = NOT(WX10713)
--	WX10717 = NOT(WX11347)
--	WX10721 = NOT(WX11348)
--	WX10725 = NOT(WX11348)
--	WX10727 = NOT(WX10718)
--	WX10728 = NOT(WX10727)
--	WX10731 = NOT(WX11347)
--	WX10735 = NOT(WX11348)
--	WX10739 = NOT(WX11348)
--	WX10741 = NOT(WX10732)
--	WX10742 = NOT(WX10741)
--	WX10745 = NOT(WX11347)
--	WX10749 = NOT(WX11348)
--	WX10753 = NOT(WX11348)
--	WX10755 = NOT(WX10746)
--	WX10756 = NOT(WX10755)
--	WX10759 = NOT(WX11347)
--	WX10763 = NOT(WX11348)
--	WX10767 = NOT(WX11348)
--	WX10769 = NOT(WX10760)
--	WX10770 = NOT(WX10769)
--	WX10773 = NOT(WX11347)
--	WX10777 = NOT(WX11348)
--	WX10781 = NOT(WX11348)
--	WX10783 = NOT(WX10774)
--	WX10784 = NOT(WX10783)
--	WX10787 = NOT(WX11347)
--	WX10791 = NOT(WX11348)
--	WX10795 = NOT(WX11348)
--	WX10797 = NOT(WX10788)
--	WX10798 = NOT(WX10797)
--	WX10801 = NOT(WX11347)
--	WX10805 = NOT(WX11348)
--	WX10809 = NOT(WX11348)
--	WX10811 = NOT(WX10802)
--	WX10812 = NOT(WX10811)
--	WX10815 = NOT(WX11347)
--	WX10819 = NOT(WX11348)
--	WX10823 = NOT(WX11348)
--	WX10825 = NOT(WX10816)
--	WX10826 = NOT(WX10825)
--	WX10827 = NOT(WX10829)
--	WX10892 = NOT(WX11309)
--	WX10893 = NOT(WX11311)
--	WX10894 = NOT(WX11313)
--	WX10895 = NOT(WX11315)
--	WX10896 = NOT(WX11317)
--	WX10897 = NOT(WX11319)
--	WX10898 = NOT(WX11321)
--	WX10899 = NOT(WX11323)
--	WX10900 = NOT(WX11325)
--	WX10901 = NOT(WX11327)
--	WX10902 = NOT(WX11329)
--	WX10903 = NOT(WX11331)
--	WX10904 = NOT(WX11333)
--	WX10905 = NOT(WX11335)
--	WX10906 = NOT(WX11337)
--	WX10907 = NOT(WX11339)
--	WX10908 = NOT(WX11277)
--	WX10909 = NOT(WX11279)
--	WX10910 = NOT(WX11281)
--	WX10911 = NOT(WX11283)
--	WX10912 = NOT(WX11285)
--	WX10913 = NOT(WX11287)
--	WX10914 = NOT(WX11289)
--	WX10915 = NOT(WX11291)
--	WX10916 = NOT(WX11293)
--	WX10917 = NOT(WX11295)
--	WX10918 = NOT(WX11297)
--	WX10919 = NOT(WX11299)
--	WX10920 = NOT(WX11301)
--	WX10921 = NOT(WX11303)
--	WX10922 = NOT(WX11305)
--	WX10923 = NOT(WX11307)
--	WX10924 = NOT(WX10892)
--	WX10925 = NOT(WX10893)
--	WX10926 = NOT(WX10894)
--	WX10927 = NOT(WX10895)
--	WX10928 = NOT(WX10896)
--	WX10929 = NOT(WX10897)
--	WX10930 = NOT(WX10898)
--	WX10931 = NOT(WX10899)
--	WX10932 = NOT(WX10900)
--	WX10933 = NOT(WX10901)
--	WX10934 = NOT(WX10902)
--	WX10935 = NOT(WX10903)
--	WX10936 = NOT(WX10904)
--	WX10937 = NOT(WX10905)
--	WX10938 = NOT(WX10906)
--	WX10939 = NOT(WX10907)
--	WX10940 = NOT(WX10908)
--	WX10941 = NOT(WX10909)
--	WX10942 = NOT(WX10910)
--	WX10943 = NOT(WX10911)
--	WX10944 = NOT(WX10912)
--	WX10945 = NOT(WX10913)
--	WX10946 = NOT(WX10914)
--	WX10947 = NOT(WX10915)
--	WX10948 = NOT(WX10916)
--	WX10949 = NOT(WX10917)
--	WX10950 = NOT(WX10918)
--	WX10951 = NOT(WX10919)
--	WX10952 = NOT(WX10920)
--	WX10953 = NOT(WX10921)
--	WX10954 = NOT(WX10922)
--	WX10955 = NOT(WX10923)
--	WX10956 = NOT(WX11181)
--	WX10957 = NOT(WX11183)
--	WX10958 = NOT(WX11185)
--	WX10959 = NOT(WX11187)
--	WX10960 = NOT(WX11189)
--	WX10961 = NOT(WX11191)
--	WX10962 = NOT(WX11193)
--	WX10963 = NOT(WX11195)
--	WX10964 = NOT(WX11197)
--	WX10965 = NOT(WX11199)
--	WX10966 = NOT(WX11201)
--	WX10967 = NOT(WX11203)
--	WX10968 = NOT(WX11205)
--	WX10969 = NOT(WX11207)
--	WX10970 = NOT(WX11209)
--	WX10971 = NOT(WX11211)
--	WX10972 = NOT(WX11213)
--	WX10973 = NOT(WX11215)
--	WX10974 = NOT(WX11217)
--	WX10975 = NOT(WX11219)
--	WX10976 = NOT(WX11221)
--	WX10977 = NOT(WX11223)
--	WX10978 = NOT(WX11225)
--	WX10979 = NOT(WX11227)
--	WX10980 = NOT(WX11229)
--	WX10981 = NOT(WX11231)
--	WX10982 = NOT(WX11233)
--	WX10983 = NOT(WX11235)
--	WX10984 = NOT(WX11237)
--	WX10985 = NOT(WX11239)
--	WX10986 = NOT(WX11241)
--	WX10987 = NOT(WX11243)
--	WX11276 = NOT(WX11260)
--	WX11277 = NOT(WX11276)
--	WX11278 = NOT(WX11261)
--	WX11279 = NOT(WX11278)
--	WX11280 = NOT(WX11262)
--	WX11281 = NOT(WX11280)
--	WX11282 = NOT(WX11263)
--	WX11283 = NOT(WX11282)
--	WX11284 = NOT(WX11264)
--	WX11285 = NOT(WX11284)
--	WX11286 = NOT(WX11265)
--	WX11287 = NOT(WX11286)
--	WX11288 = NOT(WX11266)
--	WX11289 = NOT(WX11288)
--	WX11290 = NOT(WX11267)
--	WX11291 = NOT(WX11290)
--	WX11292 = NOT(WX11268)
--	WX11293 = NOT(WX11292)
--	WX11294 = NOT(WX11269)
--	WX11295 = NOT(WX11294)
--	WX11296 = NOT(WX11270)
--	WX11297 = NOT(WX11296)
--	WX11298 = NOT(WX11271)
--	WX11299 = NOT(WX11298)
--	WX11300 = NOT(WX11272)
--	WX11301 = NOT(WX11300)
--	WX11302 = NOT(WX11273)
--	WX11303 = NOT(WX11302)
--	WX11304 = NOT(WX11274)
--	WX11305 = NOT(WX11304)
--	WX11306 = NOT(WX11275)
--	WX11307 = NOT(WX11306)
--	WX11308 = NOT(WX11244)
--	WX11309 = NOT(WX11308)
--	WX11310 = NOT(WX11245)
--	WX11311 = NOT(WX11310)
--	WX11312 = NOT(WX11246)
--	WX11313 = NOT(WX11312)
--	WX11314 = NOT(WX11247)
--	WX11315 = NOT(WX11314)
--	WX11316 = NOT(WX11248)
--	WX11317 = NOT(WX11316)
--	WX11318 = NOT(WX11249)
--	WX11319 = NOT(WX11318)
--	WX11320 = NOT(WX11250)
--	WX11321 = NOT(WX11320)
--	WX11322 = NOT(WX11251)
--	WX11323 = NOT(WX11322)
--	WX11324 = NOT(WX11252)
--	WX11325 = NOT(WX11324)
--	WX11326 = NOT(WX11253)
--	WX11327 = NOT(WX11326)
--	WX11328 = NOT(WX11254)
--	WX11329 = NOT(WX11328)
--	WX11330 = NOT(WX11255)
--	WX11331 = NOT(WX11330)
--	WX11332 = NOT(WX11256)
--	WX11333 = NOT(WX11332)
--	WX11334 = NOT(WX11257)
--	WX11335 = NOT(WX11334)
--	WX11336 = NOT(WX11258)
--	WX11337 = NOT(WX11336)
--	WX11338 = NOT(WX11259)
--	WX11339 = NOT(WX11338)
--	WX11340 = NOT(TM0)
--	WX11341 = NOT(TM0)
--	WX11342 = NOT(TM0)
--	WX11343 = NOT(TM1)
--	WX11344 = NOT(TM1)
--	WX11345 = NOT(WX11344)
--	WX11346 = NOT(WX11342)
--	WX11347 = NOT(WX11343)
--	WX11348 = NOT(WX11341)
--	WX11349 = NOT(WX11340)
--	WX11353 = NOT(WX11349)
--	WX11355 = NOT(WX11354)
--	WX11356 = NOT(WX11355)
--	WX11360 = NOT(WX11349)
--	WX11362 = NOT(WX11361)
--	WX11363 = NOT(WX11362)
--	WX11367 = NOT(WX11349)
--	WX11369 = NOT(WX11368)
--	WX11370 = NOT(WX11369)
--	WX11374 = NOT(WX11349)
--	WX11376 = NOT(WX11375)
--	WX11377 = NOT(WX11376)
--	WX11381 = NOT(WX11349)
--	WX11383 = NOT(WX11382)
--	WX11384 = NOT(WX11383)
--	WX11388 = NOT(WX11349)
--	WX11390 = NOT(WX11389)
--	WX11391 = NOT(WX11390)
--	WX11395 = NOT(WX11349)
--	WX11397 = NOT(WX11396)
--	WX11398 = NOT(WX11397)
--	WX11402 = NOT(WX11349)
--	WX11404 = NOT(WX11403)
--	WX11405 = NOT(WX11404)
--	WX11409 = NOT(WX11349)
--	WX11411 = NOT(WX11410)
--	WX11412 = NOT(WX11411)
--	WX11416 = NOT(WX11349)
--	WX11418 = NOT(WX11417)
--	WX11419 = NOT(WX11418)
--	WX11423 = NOT(WX11349)
--	WX11425 = NOT(WX11424)
--	WX11426 = NOT(WX11425)
--	WX11430 = NOT(WX11349)
--	WX11432 = NOT(WX11431)
--	WX11433 = NOT(WX11432)
--	WX11437 = NOT(WX11349)
--	WX11439 = NOT(WX11438)
--	WX11440 = NOT(WX11439)
--	WX11444 = NOT(WX11349)
--	WX11446 = NOT(WX11445)
--	WX11447 = NOT(WX11446)
--	WX11451 = NOT(WX11349)
--	WX11453 = NOT(WX11452)
--	WX11454 = NOT(WX11453)
--	WX11458 = NOT(WX11349)
--	WX11460 = NOT(WX11459)
--	WX11461 = NOT(WX11460)
--	WX11465 = NOT(WX11349)
--	WX11467 = NOT(WX11466)
--	WX11468 = NOT(WX11467)
--	WX11472 = NOT(WX11349)
--	WX11474 = NOT(WX11473)
--	WX11475 = NOT(WX11474)
--	WX11479 = NOT(WX11349)
--	WX11481 = NOT(WX11480)
--	WX11482 = NOT(WX11481)
--	WX11486 = NOT(WX11349)
--	WX11488 = NOT(WX11487)
--	WX11489 = NOT(WX11488)
--	WX11493 = NOT(WX11349)
--	WX11495 = NOT(WX11494)
--	WX11496 = NOT(WX11495)
--	WX11500 = NOT(WX11349)
--	WX11502 = NOT(WX11501)
--	WX11503 = NOT(WX11502)
--	WX11507 = NOT(WX11349)
--	WX11509 = NOT(WX11508)
--	WX11510 = NOT(WX11509)
--	WX11514 = NOT(WX11349)
--	WX11516 = NOT(WX11515)
--	WX11517 = NOT(WX11516)
--	WX11521 = NOT(WX11349)
--	WX11523 = NOT(WX11522)
--	WX11524 = NOT(WX11523)
--	WX11528 = NOT(WX11349)
--	WX11530 = NOT(WX11529)
--	WX11531 = NOT(WX11530)
--	WX11535 = NOT(WX11349)
--	WX11537 = NOT(WX11536)
--	WX11538 = NOT(WX11537)
--	WX11542 = NOT(WX11349)
--	WX11544 = NOT(WX11543)
--	WX11545 = NOT(WX11544)
--	WX11549 = NOT(WX11349)
--	WX11551 = NOT(WX11550)
--	WX11552 = NOT(WX11551)
--	WX11556 = NOT(WX11349)
--	WX11558 = NOT(WX11557)
--	WX11559 = NOT(WX11558)
--	WX11563 = NOT(WX11349)
--	WX11565 = NOT(WX11564)
--	WX11566 = NOT(WX11565)
--	WX11570 = NOT(WX11349)
--	WX11572 = NOT(WX11571)
--	WX11573 = NOT(WX11572)
--	WX11574 = NOT(RESET)
--	WX11607 = NOT(WX11574)
--	
--	WX35 = AND(WX46, WX1003)
--	WX36 = AND(WX42, WX37)
--	WX39 = AND(CRC_OUT_9_31, WX1004)
--	WX40 = AND(WX2305, WX41)
--	WX43 = AND(WX485, WX1004)
--	WX44 = AND(DATA_9_31, WX45)
--	WX49 = AND(WX60, WX1003)
--	WX50 = AND(WX56, WX51)
--	WX53 = AND(CRC_OUT_9_30, WX1004)
--	WX54 = AND(WX2312, WX55)
--	WX57 = AND(WX487, WX1004)
--	WX58 = AND(DATA_9_30, WX59)
--	WX63 = AND(WX74, WX1003)
--	WX64 = AND(WX70, WX65)
--	WX67 = AND(CRC_OUT_9_29, WX1004)
--	WX68 = AND(WX2319, WX69)
--	WX71 = AND(WX489, WX1004)
--	WX72 = AND(DATA_9_29, WX73)
--	WX77 = AND(WX88, WX1003)
--	WX78 = AND(WX84, WX79)
--	WX81 = AND(CRC_OUT_9_28, WX1004)
--	WX82 = AND(WX2326, WX83)
--	WX85 = AND(WX491, WX1004)
--	WX86 = AND(DATA_9_28, WX87)
--	WX91 = AND(WX102, WX1003)
--	WX92 = AND(WX98, WX93)
--	WX95 = AND(CRC_OUT_9_27, WX1004)
--	WX96 = AND(WX2333, WX97)
--	WX99 = AND(WX493, WX1004)
--	WX100 = AND(DATA_9_27, WX101)
--	WX105 = AND(WX116, WX1003)
--	WX106 = AND(WX112, WX107)
--	WX109 = AND(CRC_OUT_9_26, WX1004)
--	WX110 = AND(WX2340, WX111)
--	WX113 = AND(WX495, WX1004)
--	WX114 = AND(DATA_9_26, WX115)
--	WX119 = AND(WX130, WX1003)
--	WX120 = AND(WX126, WX121)
--	WX123 = AND(CRC_OUT_9_25, WX1004)
--	WX124 = AND(WX2347, WX125)
--	WX127 = AND(WX497, WX1004)
--	WX128 = AND(DATA_9_25, WX129)
--	WX133 = AND(WX144, WX1003)
--	WX134 = AND(WX140, WX135)
--	WX137 = AND(CRC_OUT_9_24, WX1004)
--	WX138 = AND(WX2354, WX139)
--	WX141 = AND(WX499, WX1004)
--	WX142 = AND(DATA_9_24, WX143)
--	WX147 = AND(WX158, WX1003)
--	WX148 = AND(WX154, WX149)
--	WX151 = AND(CRC_OUT_9_23, WX1004)
--	WX152 = AND(WX2361, WX153)
--	WX155 = AND(WX501, WX1004)
--	WX156 = AND(DATA_9_23, WX157)
--	WX161 = AND(WX172, WX1003)
--	WX162 = AND(WX168, WX163)
--	WX165 = AND(CRC_OUT_9_22, WX1004)
--	WX166 = AND(WX2368, WX167)
--	WX169 = AND(WX503, WX1004)
--	WX170 = AND(DATA_9_22, WX171)
--	WX175 = AND(WX186, WX1003)
--	WX176 = AND(WX182, WX177)
--	WX179 = AND(CRC_OUT_9_21, WX1004)
--	WX180 = AND(WX2375, WX181)
--	WX183 = AND(WX505, WX1004)
--	WX184 = AND(DATA_9_21, WX185)
--	WX189 = AND(WX200, WX1003)
--	WX190 = AND(WX196, WX191)
--	WX193 = AND(CRC_OUT_9_20, WX1004)
--	WX194 = AND(WX2382, WX195)
--	WX197 = AND(WX507, WX1004)
--	WX198 = AND(DATA_9_20, WX199)
--	WX203 = AND(WX214, WX1003)
--	WX204 = AND(WX210, WX205)
--	WX207 = AND(CRC_OUT_9_19, WX1004)
--	WX208 = AND(WX2389, WX209)
--	WX211 = AND(WX509, WX1004)
--	WX212 = AND(DATA_9_19, WX213)
--	WX217 = AND(WX228, WX1003)
--	WX218 = AND(WX224, WX219)
--	WX221 = AND(CRC_OUT_9_18, WX1004)
--	WX222 = AND(WX2396, WX223)
--	WX225 = AND(WX511, WX1004)
--	WX226 = AND(DATA_9_18, WX227)
--	WX231 = AND(WX242, WX1003)
--	WX232 = AND(WX238, WX233)
--	WX235 = AND(CRC_OUT_9_17, WX1004)
--	WX236 = AND(WX2403, WX237)
--	WX239 = AND(WX513, WX1004)
--	WX240 = AND(DATA_9_17, WX241)
--	WX245 = AND(WX256, WX1003)
--	WX246 = AND(WX252, WX247)
--	WX249 = AND(CRC_OUT_9_16, WX1004)
--	WX250 = AND(WX2410, WX251)
--	WX253 = AND(WX515, WX1004)
--	WX254 = AND(DATA_9_16, WX255)
--	WX259 = AND(WX270, WX1003)
--	WX260 = AND(WX266, WX261)
--	WX263 = AND(CRC_OUT_9_15, WX1004)
--	WX264 = AND(WX2417, WX265)
--	WX267 = AND(WX517, WX1004)
--	WX268 = AND(DATA_9_15, WX269)
--	WX273 = AND(WX284, WX1003)
--	WX274 = AND(WX280, WX275)
--	WX277 = AND(CRC_OUT_9_14, WX1004)
--	WX278 = AND(WX2424, WX279)
--	WX281 = AND(WX519, WX1004)
--	WX282 = AND(DATA_9_14, WX283)
--	WX287 = AND(WX298, WX1003)
--	WX288 = AND(WX294, WX289)
--	WX291 = AND(CRC_OUT_9_13, WX1004)
--	WX292 = AND(WX2431, WX293)
--	WX295 = AND(WX521, WX1004)
--	WX296 = AND(DATA_9_13, WX297)
--	WX301 = AND(WX312, WX1003)
--	WX302 = AND(WX308, WX303)
--	WX305 = AND(CRC_OUT_9_12, WX1004)
--	WX306 = AND(WX2438, WX307)
--	WX309 = AND(WX523, WX1004)
--	WX310 = AND(DATA_9_12, WX311)
--	WX315 = AND(WX326, WX1003)
--	WX316 = AND(WX322, WX317)
--	WX319 = AND(CRC_OUT_9_11, WX1004)
--	WX320 = AND(WX2445, WX321)
--	WX323 = AND(WX525, WX1004)
--	WX324 = AND(DATA_9_11, WX325)
--	WX329 = AND(WX340, WX1003)
--	WX330 = AND(WX336, WX331)
--	WX333 = AND(CRC_OUT_9_10, WX1004)
--	WX334 = AND(WX2452, WX335)
--	WX337 = AND(WX527, WX1004)
--	WX338 = AND(DATA_9_10, WX339)
--	WX343 = AND(WX354, WX1003)
--	WX344 = AND(WX350, WX345)
--	WX347 = AND(CRC_OUT_9_9, WX1004)
--	WX348 = AND(WX2459, WX349)
--	WX351 = AND(WX529, WX1004)
--	WX352 = AND(DATA_9_9, WX353)
--	WX357 = AND(WX368, WX1003)
--	WX358 = AND(WX364, WX359)
--	WX361 = AND(CRC_OUT_9_8, WX1004)
--	WX362 = AND(WX2466, WX363)
--	WX365 = AND(WX531, WX1004)
--	WX366 = AND(DATA_9_8, WX367)
--	WX371 = AND(WX382, WX1003)
--	WX372 = AND(WX378, WX373)
--	WX375 = AND(CRC_OUT_9_7, WX1004)
--	WX376 = AND(WX2473, WX377)
--	WX379 = AND(WX533, WX1004)
--	WX380 = AND(DATA_9_7, WX381)
--	WX385 = AND(WX396, WX1003)
--	WX386 = AND(WX392, WX387)
--	WX389 = AND(CRC_OUT_9_6, WX1004)
--	WX390 = AND(WX2480, WX391)
--	WX393 = AND(WX535, WX1004)
--	WX394 = AND(DATA_9_6, WX395)
--	WX399 = AND(WX410, WX1003)
--	WX400 = AND(WX406, WX401)
--	WX403 = AND(CRC_OUT_9_5, WX1004)
--	WX404 = AND(WX2487, WX405)
--	WX407 = AND(WX537, WX1004)
--	WX408 = AND(DATA_9_5, WX409)
--	WX413 = AND(WX424, WX1003)
--	WX414 = AND(WX420, WX415)
--	WX417 = AND(CRC_OUT_9_4, WX1004)
--	WX418 = AND(WX2494, WX419)
--	WX421 = AND(WX539, WX1004)
--	WX422 = AND(DATA_9_4, WX423)
--	WX427 = AND(WX438, WX1003)
--	WX428 = AND(WX434, WX429)
--	WX431 = AND(CRC_OUT_9_3, WX1004)
--	WX432 = AND(WX2501, WX433)
--	WX435 = AND(WX541, WX1004)
--	WX436 = AND(DATA_9_3, WX437)
--	WX441 = AND(WX452, WX1003)
--	WX442 = AND(WX448, WX443)
--	WX445 = AND(CRC_OUT_9_2, WX1004)
--	WX446 = AND(WX2508, WX447)
--	WX449 = AND(WX543, WX1004)
--	WX450 = AND(DATA_9_2, WX451)
--	WX455 = AND(WX466, WX1003)
--	WX456 = AND(WX462, WX457)
--	WX459 = AND(CRC_OUT_9_1, WX1004)
--	WX460 = AND(WX2515, WX461)
--	WX463 = AND(WX545, WX1004)
--	WX464 = AND(DATA_9_1, WX465)
--	WX469 = AND(WX480, WX1003)
--	WX470 = AND(WX476, WX471)
--	WX473 = AND(CRC_OUT_9_0, WX1004)
--	WX474 = AND(WX2522, WX475)
--	WX477 = AND(WX547, WX1004)
--	WX478 = AND(DATA_9_0, WX479)
--	WX484 = AND(WX487, RESET)
--	WX486 = AND(WX489, RESET)
--	WX488 = AND(WX491, RESET)
--	WX490 = AND(WX493, RESET)
--	WX492 = AND(WX495, RESET)
--	WX494 = AND(WX497, RESET)
--	WX496 = AND(WX499, RESET)
--	WX498 = AND(WX501, RESET)
--	WX500 = AND(WX503, RESET)
--	WX502 = AND(WX505, RESET)
--	WX504 = AND(WX507, RESET)
--	WX506 = AND(WX509, RESET)
--	WX508 = AND(WX511, RESET)
--	WX510 = AND(WX513, RESET)
--	WX512 = AND(WX515, RESET)
--	WX514 = AND(WX517, RESET)
--	WX516 = AND(WX519, RESET)
--	WX518 = AND(WX521, RESET)
--	WX520 = AND(WX523, RESET)
--	WX522 = AND(WX525, RESET)
--	WX524 = AND(WX527, RESET)
--	WX526 = AND(WX529, RESET)
--	WX528 = AND(WX531, RESET)
--	WX530 = AND(WX533, RESET)
--	WX532 = AND(WX535, RESET)
--	WX534 = AND(WX537, RESET)
--	WX536 = AND(WX539, RESET)
--	WX538 = AND(WX541, RESET)
--	WX540 = AND(WX543, RESET)
--	WX542 = AND(WX545, RESET)
--	WX544 = AND(WX547, RESET)
--	WX546 = AND(WX483, RESET)
--	WX644 = AND(WX48, RESET)
--	WX646 = AND(WX62, RESET)
--	WX648 = AND(WX76, RESET)
--	WX650 = AND(WX90, RESET)
--	WX652 = AND(WX104, RESET)
--	WX654 = AND(WX118, RESET)
--	WX656 = AND(WX132, RESET)
--	WX658 = AND(WX146, RESET)
--	WX660 = AND(WX160, RESET)
--	WX662 = AND(WX174, RESET)
--	WX664 = AND(WX188, RESET)
--	WX666 = AND(WX202, RESET)
--	WX668 = AND(WX216, RESET)
--	WX670 = AND(WX230, RESET)
--	WX672 = AND(WX244, RESET)
--	WX674 = AND(WX258, RESET)
--	WX676 = AND(WX272, RESET)
--	WX678 = AND(WX286, RESET)
--	WX680 = AND(WX300, RESET)
--	WX682 = AND(WX314, RESET)
--	WX684 = AND(WX328, RESET)
--	WX686 = AND(WX342, RESET)
--	WX688 = AND(WX356, RESET)
--	WX690 = AND(WX370, RESET)
--	WX692 = AND(WX384, RESET)
--	WX694 = AND(WX398, RESET)
--	WX696 = AND(WX412, RESET)
--	WX698 = AND(WX426, RESET)
--	WX700 = AND(WX440, RESET)
--	WX702 = AND(WX454, RESET)
--	WX704 = AND(WX468, RESET)
--	WX706 = AND(WX482, RESET)
--	WX708 = AND(WX645, RESET)
--	WX710 = AND(WX647, RESET)
--	WX712 = AND(WX649, RESET)
--	WX714 = AND(WX651, RESET)
--	WX716 = AND(WX653, RESET)
--	WX718 = AND(WX655, RESET)
--	WX720 = AND(WX657, RESET)
--	WX722 = AND(WX659, RESET)
--	WX724 = AND(WX661, RESET)
--	WX726 = AND(WX663, RESET)
--	WX728 = AND(WX665, RESET)
--	WX730 = AND(WX667, RESET)
--	WX732 = AND(WX669, RESET)
--	WX734 = AND(WX671, RESET)
--	WX736 = AND(WX673, RESET)
--	WX738 = AND(WX675, RESET)
--	WX740 = AND(WX677, RESET)
--	WX742 = AND(WX679, RESET)
--	WX744 = AND(WX681, RESET)
--	WX746 = AND(WX683, RESET)
--	WX748 = AND(WX685, RESET)
--	WX750 = AND(WX687, RESET)
--	WX752 = AND(WX689, RESET)
--	WX754 = AND(WX691, RESET)
--	WX756 = AND(WX693, RESET)
--	WX758 = AND(WX695, RESET)
--	WX760 = AND(WX697, RESET)
--	WX762 = AND(WX699, RESET)
--	WX764 = AND(WX701, RESET)
--	WX766 = AND(WX703, RESET)
--	WX768 = AND(WX705, RESET)
--	WX770 = AND(WX707, RESET)
--	WX772 = AND(WX709, RESET)
--	WX774 = AND(WX711, RESET)
--	WX776 = AND(WX713, RESET)
--	WX778 = AND(WX715, RESET)
--	WX780 = AND(WX717, RESET)
--	WX782 = AND(WX719, RESET)
--	WX784 = AND(WX721, RESET)
--	WX786 = AND(WX723, RESET)
--	WX788 = AND(WX725, RESET)
--	WX790 = AND(WX727, RESET)
--	WX792 = AND(WX729, RESET)
--	WX794 = AND(WX731, RESET)
--	WX796 = AND(WX733, RESET)
--	WX798 = AND(WX735, RESET)
--	WX800 = AND(WX737, RESET)
--	WX802 = AND(WX739, RESET)
--	WX804 = AND(WX741, RESET)
--	WX806 = AND(WX743, RESET)
--	WX808 = AND(WX745, RESET)
--	WX810 = AND(WX747, RESET)
--	WX812 = AND(WX749, RESET)
--	WX814 = AND(WX751, RESET)
--	WX816 = AND(WX753, RESET)
--	WX818 = AND(WX755, RESET)
--	WX820 = AND(WX757, RESET)
--	WX822 = AND(WX759, RESET)
--	WX824 = AND(WX761, RESET)
--	WX826 = AND(WX763, RESET)
--	WX828 = AND(WX765, RESET)
--	WX830 = AND(WX767, RESET)
--	WX832 = AND(WX769, RESET)
--	WX834 = AND(WX771, RESET)
--	WX836 = AND(WX773, RESET)
--	WX838 = AND(WX775, RESET)
--	WX840 = AND(WX777, RESET)
--	WX842 = AND(WX779, RESET)
--	WX844 = AND(WX781, RESET)
--	WX846 = AND(WX783, RESET)
--	WX848 = AND(WX785, RESET)
--	WX850 = AND(WX787, RESET)
--	WX852 = AND(WX789, RESET)
--	WX854 = AND(WX791, RESET)
--	WX856 = AND(WX793, RESET)
--	WX858 = AND(WX795, RESET)
--	WX860 = AND(WX797, RESET)
--	WX862 = AND(WX799, RESET)
--	WX864 = AND(WX801, RESET)
--	WX866 = AND(WX803, RESET)
--	WX868 = AND(WX805, RESET)
--	WX870 = AND(WX807, RESET)
--	WX872 = AND(WX809, RESET)
--	WX874 = AND(WX811, RESET)
--	WX876 = AND(WX813, RESET)
--	WX878 = AND(WX815, RESET)
--	WX880 = AND(WX817, RESET)
--	WX882 = AND(WX819, RESET)
--	WX884 = AND(WX821, RESET)
--	WX886 = AND(WX823, RESET)
--	WX888 = AND(WX825, RESET)
--	WX890 = AND(WX827, RESET)
--	WX892 = AND(WX829, RESET)
--	WX894 = AND(WX831, RESET)
--	WX896 = AND(WX833, RESET)
--	WX898 = AND(WX835, RESET)
--	WX1007 = AND(WX1006, WX1005)
--	WX1008 = AND(WX580, WX1009)
--	WX1014 = AND(WX1013, WX1005)
--	WX1015 = AND(WX581, WX1016)
--	WX1021 = AND(WX1020, WX1005)
--	WX1022 = AND(WX582, WX1023)
--	WX1028 = AND(WX1027, WX1005)
--	WX1029 = AND(WX583, WX1030)
--	WX1035 = AND(WX1034, WX1005)
--	WX1036 = AND(WX584, WX1037)
--	WX1042 = AND(WX1041, WX1005)
--	WX1043 = AND(WX585, WX1044)
--	WX1049 = AND(WX1048, WX1005)
--	WX1050 = AND(WX586, WX1051)
--	WX1056 = AND(WX1055, WX1005)
--	WX1057 = AND(WX587, WX1058)
--	WX1063 = AND(WX1062, WX1005)
--	WX1064 = AND(WX588, WX1065)
--	WX1070 = AND(WX1069, WX1005)
--	WX1071 = AND(WX589, WX1072)
--	WX1077 = AND(WX1076, WX1005)
--	WX1078 = AND(WX590, WX1079)
--	WX1084 = AND(WX1083, WX1005)
--	WX1085 = AND(WX591, WX1086)
--	WX1091 = AND(WX1090, WX1005)
--	WX1092 = AND(WX592, WX1093)
--	WX1098 = AND(WX1097, WX1005)
--	WX1099 = AND(WX593, WX1100)
--	WX1105 = AND(WX1104, WX1005)
--	WX1106 = AND(WX594, WX1107)
--	WX1112 = AND(WX1111, WX1005)
--	WX1113 = AND(WX595, WX1114)
--	WX1119 = AND(WX1118, WX1005)
--	WX1120 = AND(WX596, WX1121)
--	WX1126 = AND(WX1125, WX1005)
--	WX1127 = AND(WX597, WX1128)
--	WX1133 = AND(WX1132, WX1005)
--	WX1134 = AND(WX598, WX1135)
--	WX1140 = AND(WX1139, WX1005)
--	WX1141 = AND(WX599, WX1142)
--	WX1147 = AND(WX1146, WX1005)
--	WX1148 = AND(WX600, WX1149)
--	WX1154 = AND(WX1153, WX1005)
--	WX1155 = AND(WX601, WX1156)
--	WX1161 = AND(WX1160, WX1005)
--	WX1162 = AND(WX602, WX1163)
--	WX1168 = AND(WX1167, WX1005)
--	WX1169 = AND(WX603, WX1170)
--	WX1175 = AND(WX1174, WX1005)
--	WX1176 = AND(WX604, WX1177)
--	WX1182 = AND(WX1181, WX1005)
--	WX1183 = AND(WX605, WX1184)
--	WX1189 = AND(WX1188, WX1005)
--	WX1190 = AND(WX606, WX1191)
--	WX1196 = AND(WX1195, WX1005)
--	WX1197 = AND(WX607, WX1198)
--	WX1203 = AND(WX1202, WX1005)
--	WX1204 = AND(WX608, WX1205)
--	WX1210 = AND(WX1209, WX1005)
--	WX1211 = AND(WX609, WX1212)
--	WX1217 = AND(WX1216, WX1005)
--	WX1218 = AND(WX610, WX1219)
--	WX1224 = AND(WX1223, WX1005)
--	WX1225 = AND(WX611, WX1226)
--	WX1264 = AND(WX1234, WX1263)
--	WX1266 = AND(WX1262, WX1263)
--	WX1268 = AND(WX1261, WX1263)
--	WX1270 = AND(WX1260, WX1263)
--	WX1272 = AND(WX1233, WX1263)
--	WX1274 = AND(WX1259, WX1263)
--	WX1276 = AND(WX1258, WX1263)
--	WX1278 = AND(WX1257, WX1263)
--	WX1280 = AND(WX1256, WX1263)
--	WX1282 = AND(WX1255, WX1263)
--	WX1284 = AND(WX1254, WX1263)
--	WX1286 = AND(WX1232, WX1263)
--	WX1288 = AND(WX1253, WX1263)
--	WX1290 = AND(WX1252, WX1263)
--	WX1292 = AND(WX1251, WX1263)
--	WX1294 = AND(WX1250, WX1263)
--	WX1296 = AND(WX1231, WX1263)
--	WX1298 = AND(WX1249, WX1263)
--	WX1300 = AND(WX1248, WX1263)
--	WX1302 = AND(WX1247, WX1263)
--	WX1304 = AND(WX1246, WX1263)
--	WX1306 = AND(WX1245, WX1263)
--	WX1308 = AND(WX1244, WX1263)
--	WX1310 = AND(WX1243, WX1263)
--	WX1312 = AND(WX1242, WX1263)
--	WX1314 = AND(WX1241, WX1263)
--	WX1316 = AND(WX1240, WX1263)
--	WX1318 = AND(WX1239, WX1263)
--	WX1320 = AND(WX1238, WX1263)
--	WX1322 = AND(WX1237, WX1263)
--	WX1324 = AND(WX1236, WX1263)
--	WX1326 = AND(WX1235, WX1263)
--	WX1328 = AND(WX1339, WX2296)
--	WX1329 = AND(WX1335, WX1330)
--	WX1332 = AND(CRC_OUT_8_31, WX2297)
--	WX1333 = AND(WX3598, WX1334)
--	WX1336 = AND(WX1778, WX2297)
--	WX1337 = AND(WX2305, WX1338)
--	WX1342 = AND(WX1353, WX2296)
--	WX1343 = AND(WX1349, WX1344)
--	WX1346 = AND(CRC_OUT_8_30, WX2297)
--	WX1347 = AND(WX3605, WX1348)
--	WX1350 = AND(WX1780, WX2297)
--	WX1351 = AND(WX2312, WX1352)
--	WX1356 = AND(WX1367, WX2296)
--	WX1357 = AND(WX1363, WX1358)
--	WX1360 = AND(CRC_OUT_8_29, WX2297)
--	WX1361 = AND(WX3612, WX1362)
--	WX1364 = AND(WX1782, WX2297)
--	WX1365 = AND(WX2319, WX1366)
--	WX1370 = AND(WX1381, WX2296)
--	WX1371 = AND(WX1377, WX1372)
--	WX1374 = AND(CRC_OUT_8_28, WX2297)
--	WX1375 = AND(WX3619, WX1376)
--	WX1378 = AND(WX1784, WX2297)
--	WX1379 = AND(WX2326, WX1380)
--	WX1384 = AND(WX1395, WX2296)
--	WX1385 = AND(WX1391, WX1386)
--	WX1388 = AND(CRC_OUT_8_27, WX2297)
--	WX1389 = AND(WX3626, WX1390)
--	WX1392 = AND(WX1786, WX2297)
--	WX1393 = AND(WX2333, WX1394)
--	WX1398 = AND(WX1409, WX2296)
--	WX1399 = AND(WX1405, WX1400)
--	WX1402 = AND(CRC_OUT_8_26, WX2297)
--	WX1403 = AND(WX3633, WX1404)
--	WX1406 = AND(WX1788, WX2297)
--	WX1407 = AND(WX2340, WX1408)
--	WX1412 = AND(WX1423, WX2296)
--	WX1413 = AND(WX1419, WX1414)
--	WX1416 = AND(CRC_OUT_8_25, WX2297)
--	WX1417 = AND(WX3640, WX1418)
--	WX1420 = AND(WX1790, WX2297)
--	WX1421 = AND(WX2347, WX1422)
--	WX1426 = AND(WX1437, WX2296)
--	WX1427 = AND(WX1433, WX1428)
--	WX1430 = AND(CRC_OUT_8_24, WX2297)
--	WX1431 = AND(WX3647, WX1432)
--	WX1434 = AND(WX1792, WX2297)
--	WX1435 = AND(WX2354, WX1436)
--	WX1440 = AND(WX1451, WX2296)
--	WX1441 = AND(WX1447, WX1442)
--	WX1444 = AND(CRC_OUT_8_23, WX2297)
--	WX1445 = AND(WX3654, WX1446)
--	WX1448 = AND(WX1794, WX2297)
--	WX1449 = AND(WX2361, WX1450)
--	WX1454 = AND(WX1465, WX2296)
--	WX1455 = AND(WX1461, WX1456)
--	WX1458 = AND(CRC_OUT_8_22, WX2297)
--	WX1459 = AND(WX3661, WX1460)
--	WX1462 = AND(WX1796, WX2297)
--	WX1463 = AND(WX2368, WX1464)
--	WX1468 = AND(WX1479, WX2296)
--	WX1469 = AND(WX1475, WX1470)
--	WX1472 = AND(CRC_OUT_8_21, WX2297)
--	WX1473 = AND(WX3668, WX1474)
--	WX1476 = AND(WX1798, WX2297)
--	WX1477 = AND(WX2375, WX1478)
--	WX1482 = AND(WX1493, WX2296)
--	WX1483 = AND(WX1489, WX1484)
--	WX1486 = AND(CRC_OUT_8_20, WX2297)
--	WX1487 = AND(WX3675, WX1488)
--	WX1490 = AND(WX1800, WX2297)
--	WX1491 = AND(WX2382, WX1492)
--	WX1496 = AND(WX1507, WX2296)
--	WX1497 = AND(WX1503, WX1498)
--	WX1500 = AND(CRC_OUT_8_19, WX2297)
--	WX1501 = AND(WX3682, WX1502)
--	WX1504 = AND(WX1802, WX2297)
--	WX1505 = AND(WX2389, WX1506)
--	WX1510 = AND(WX1521, WX2296)
--	WX1511 = AND(WX1517, WX1512)
--	WX1514 = AND(CRC_OUT_8_18, WX2297)
--	WX1515 = AND(WX3689, WX1516)
--	WX1518 = AND(WX1804, WX2297)
--	WX1519 = AND(WX2396, WX1520)
--	WX1524 = AND(WX1535, WX2296)
--	WX1525 = AND(WX1531, WX1526)
--	WX1528 = AND(CRC_OUT_8_17, WX2297)
--	WX1529 = AND(WX3696, WX1530)
--	WX1532 = AND(WX1806, WX2297)
--	WX1533 = AND(WX2403, WX1534)
--	WX1538 = AND(WX1549, WX2296)
--	WX1539 = AND(WX1545, WX1540)
--	WX1542 = AND(CRC_OUT_8_16, WX2297)
--	WX1543 = AND(WX3703, WX1544)
--	WX1546 = AND(WX1808, WX2297)
--	WX1547 = AND(WX2410, WX1548)
--	WX1552 = AND(WX1563, WX2296)
--	WX1553 = AND(WX1559, WX1554)
--	WX1556 = AND(CRC_OUT_8_15, WX2297)
--	WX1557 = AND(WX3710, WX1558)
--	WX1560 = AND(WX1810, WX2297)
--	WX1561 = AND(WX2417, WX1562)
--	WX1566 = AND(WX1577, WX2296)
--	WX1567 = AND(WX1573, WX1568)
--	WX1570 = AND(CRC_OUT_8_14, WX2297)
--	WX1571 = AND(WX3717, WX1572)
--	WX1574 = AND(WX1812, WX2297)
--	WX1575 = AND(WX2424, WX1576)
--	WX1580 = AND(WX1591, WX2296)
--	WX1581 = AND(WX1587, WX1582)
--	WX1584 = AND(CRC_OUT_8_13, WX2297)
--	WX1585 = AND(WX3724, WX1586)
--	WX1588 = AND(WX1814, WX2297)
--	WX1589 = AND(WX2431, WX1590)
--	WX1594 = AND(WX1605, WX2296)
--	WX1595 = AND(WX1601, WX1596)
--	WX1598 = AND(CRC_OUT_8_12, WX2297)
--	WX1599 = AND(WX3731, WX1600)
--	WX1602 = AND(WX1816, WX2297)
--	WX1603 = AND(WX2438, WX1604)
--	WX1608 = AND(WX1619, WX2296)
--	WX1609 = AND(WX1615, WX1610)
--	WX1612 = AND(CRC_OUT_8_11, WX2297)
--	WX1613 = AND(WX3738, WX1614)
--	WX1616 = AND(WX1818, WX2297)
--	WX1617 = AND(WX2445, WX1618)
--	WX1622 = AND(WX1633, WX2296)
--	WX1623 = AND(WX1629, WX1624)
--	WX1626 = AND(CRC_OUT_8_10, WX2297)
--	WX1627 = AND(WX3745, WX1628)
--	WX1630 = AND(WX1820, WX2297)
--	WX1631 = AND(WX2452, WX1632)
--	WX1636 = AND(WX1647, WX2296)
--	WX1637 = AND(WX1643, WX1638)
--	WX1640 = AND(CRC_OUT_8_9, WX2297)
--	WX1641 = AND(WX3752, WX1642)
--	WX1644 = AND(WX1822, WX2297)
--	WX1645 = AND(WX2459, WX1646)
--	WX1650 = AND(WX1661, WX2296)
--	WX1651 = AND(WX1657, WX1652)
--	WX1654 = AND(CRC_OUT_8_8, WX2297)
--	WX1655 = AND(WX3759, WX1656)
--	WX1658 = AND(WX1824, WX2297)
--	WX1659 = AND(WX2466, WX1660)
--	WX1664 = AND(WX1675, WX2296)
--	WX1665 = AND(WX1671, WX1666)
--	WX1668 = AND(CRC_OUT_8_7, WX2297)
--	WX1669 = AND(WX3766, WX1670)
--	WX1672 = AND(WX1826, WX2297)
--	WX1673 = AND(WX2473, WX1674)
--	WX1678 = AND(WX1689, WX2296)
--	WX1679 = AND(WX1685, WX1680)
--	WX1682 = AND(CRC_OUT_8_6, WX2297)
--	WX1683 = AND(WX3773, WX1684)
--	WX1686 = AND(WX1828, WX2297)
--	WX1687 = AND(WX2480, WX1688)
--	WX1692 = AND(WX1703, WX2296)
--	WX1693 = AND(WX1699, WX1694)
--	WX1696 = AND(CRC_OUT_8_5, WX2297)
--	WX1697 = AND(WX3780, WX1698)
--	WX1700 = AND(WX1830, WX2297)
--	WX1701 = AND(WX2487, WX1702)
--	WX1706 = AND(WX1717, WX2296)
--	WX1707 = AND(WX1713, WX1708)
--	WX1710 = AND(CRC_OUT_8_4, WX2297)
--	WX1711 = AND(WX3787, WX1712)
--	WX1714 = AND(WX1832, WX2297)
--	WX1715 = AND(WX2494, WX1716)
--	WX1720 = AND(WX1731, WX2296)
--	WX1721 = AND(WX1727, WX1722)
--	WX1724 = AND(CRC_OUT_8_3, WX2297)
--	WX1725 = AND(WX3794, WX1726)
--	WX1728 = AND(WX1834, WX2297)
--	WX1729 = AND(WX2501, WX1730)
--	WX1734 = AND(WX1745, WX2296)
--	WX1735 = AND(WX1741, WX1736)
--	WX1738 = AND(CRC_OUT_8_2, WX2297)
--	WX1739 = AND(WX3801, WX1740)
--	WX1742 = AND(WX1836, WX2297)
--	WX1743 = AND(WX2508, WX1744)
--	WX1748 = AND(WX1759, WX2296)
--	WX1749 = AND(WX1755, WX1750)
--	WX1752 = AND(CRC_OUT_8_1, WX2297)
--	WX1753 = AND(WX3808, WX1754)
--	WX1756 = AND(WX1838, WX2297)
--	WX1757 = AND(WX2515, WX1758)
--	WX1762 = AND(WX1773, WX2296)
--	WX1763 = AND(WX1769, WX1764)
--	WX1766 = AND(CRC_OUT_8_0, WX2297)
--	WX1767 = AND(WX3815, WX1768)
--	WX1770 = AND(WX1840, WX2297)
--	WX1771 = AND(WX2522, WX1772)
--	WX1777 = AND(WX1780, RESET)
--	WX1779 = AND(WX1782, RESET)
--	WX1781 = AND(WX1784, RESET)
--	WX1783 = AND(WX1786, RESET)
--	WX1785 = AND(WX1788, RESET)
--	WX1787 = AND(WX1790, RESET)
--	WX1789 = AND(WX1792, RESET)
--	WX1791 = AND(WX1794, RESET)
--	WX1793 = AND(WX1796, RESET)
--	WX1795 = AND(WX1798, RESET)
--	WX1797 = AND(WX1800, RESET)
--	WX1799 = AND(WX1802, RESET)
--	WX1801 = AND(WX1804, RESET)
--	WX1803 = AND(WX1806, RESET)
--	WX1805 = AND(WX1808, RESET)
--	WX1807 = AND(WX1810, RESET)
--	WX1809 = AND(WX1812, RESET)
--	WX1811 = AND(WX1814, RESET)
--	WX1813 = AND(WX1816, RESET)
--	WX1815 = AND(WX1818, RESET)
--	WX1817 = AND(WX1820, RESET)
--	WX1819 = AND(WX1822, RESET)
--	WX1821 = AND(WX1824, RESET)
--	WX1823 = AND(WX1826, RESET)
--	WX1825 = AND(WX1828, RESET)
--	WX1827 = AND(WX1830, RESET)
--	WX1829 = AND(WX1832, RESET)
--	WX1831 = AND(WX1834, RESET)
--	WX1833 = AND(WX1836, RESET)
--	WX1835 = AND(WX1838, RESET)
--	WX1837 = AND(WX1840, RESET)
--	WX1839 = AND(WX1776, RESET)
--	WX1937 = AND(WX1341, RESET)
--	WX1939 = AND(WX1355, RESET)
--	WX1941 = AND(WX1369, RESET)
--	WX1943 = AND(WX1383, RESET)
--	WX1945 = AND(WX1397, RESET)
--	WX1947 = AND(WX1411, RESET)
--	WX1949 = AND(WX1425, RESET)
--	WX1951 = AND(WX1439, RESET)
--	WX1953 = AND(WX1453, RESET)
--	WX1955 = AND(WX1467, RESET)
--	WX1957 = AND(WX1481, RESET)
--	WX1959 = AND(WX1495, RESET)
--	WX1961 = AND(WX1509, RESET)
--	WX1963 = AND(WX1523, RESET)
--	WX1965 = AND(WX1537, RESET)
--	WX1967 = AND(WX1551, RESET)
--	WX1969 = AND(WX1565, RESET)
--	WX1971 = AND(WX1579, RESET)
--	WX1973 = AND(WX1593, RESET)
--	WX1975 = AND(WX1607, RESET)
--	WX1977 = AND(WX1621, RESET)
--	WX1979 = AND(WX1635, RESET)
--	WX1981 = AND(WX1649, RESET)
--	WX1983 = AND(WX1663, RESET)
--	WX1985 = AND(WX1677, RESET)
--	WX1987 = AND(WX1691, RESET)
--	WX1989 = AND(WX1705, RESET)
--	WX1991 = AND(WX1719, RESET)
--	WX1993 = AND(WX1733, RESET)
--	WX1995 = AND(WX1747, RESET)
--	WX1997 = AND(WX1761, RESET)
--	WX1999 = AND(WX1775, RESET)
--	WX2001 = AND(WX1938, RESET)
--	WX2003 = AND(WX1940, RESET)
--	WX2005 = AND(WX1942, RESET)
--	WX2007 = AND(WX1944, RESET)
--	WX2009 = AND(WX1946, RESET)
--	WX2011 = AND(WX1948, RESET)
--	WX2013 = AND(WX1950, RESET)
--	WX2015 = AND(WX1952, RESET)
--	WX2017 = AND(WX1954, RESET)
--	WX2019 = AND(WX1956, RESET)
--	WX2021 = AND(WX1958, RESET)
--	WX2023 = AND(WX1960, RESET)
--	WX2025 = AND(WX1962, RESET)
--	WX2027 = AND(WX1964, RESET)
--	WX2029 = AND(WX1966, RESET)
--	WX2031 = AND(WX1968, RESET)
--	WX2033 = AND(WX1970, RESET)
--	WX2035 = AND(WX1972, RESET)
--	WX2037 = AND(WX1974, RESET)
--	WX2039 = AND(WX1976, RESET)
--	WX2041 = AND(WX1978, RESET)
--	WX2043 = AND(WX1980, RESET)
--	WX2045 = AND(WX1982, RESET)
--	WX2047 = AND(WX1984, RESET)
--	WX2049 = AND(WX1986, RESET)
--	WX2051 = AND(WX1988, RESET)
--	WX2053 = AND(WX1990, RESET)
--	WX2055 = AND(WX1992, RESET)
--	WX2057 = AND(WX1994, RESET)
--	WX2059 = AND(WX1996, RESET)
--	WX2061 = AND(WX1998, RESET)
--	WX2063 = AND(WX2000, RESET)
--	WX2065 = AND(WX2002, RESET)
--	WX2067 = AND(WX2004, RESET)
--	WX2069 = AND(WX2006, RESET)
--	WX2071 = AND(WX2008, RESET)
--	WX2073 = AND(WX2010, RESET)
--	WX2075 = AND(WX2012, RESET)
--	WX2077 = AND(WX2014, RESET)
--	WX2079 = AND(WX2016, RESET)
--	WX2081 = AND(WX2018, RESET)
--	WX2083 = AND(WX2020, RESET)
--	WX2085 = AND(WX2022, RESET)
--	WX2087 = AND(WX2024, RESET)
--	WX2089 = AND(WX2026, RESET)
--	WX2091 = AND(WX2028, RESET)
--	WX2093 = AND(WX2030, RESET)
--	WX2095 = AND(WX2032, RESET)
--	WX2097 = AND(WX2034, RESET)
--	WX2099 = AND(WX2036, RESET)
--	WX2101 = AND(WX2038, RESET)
--	WX2103 = AND(WX2040, RESET)
--	WX2105 = AND(WX2042, RESET)
--	WX2107 = AND(WX2044, RESET)
--	WX2109 = AND(WX2046, RESET)
--	WX2111 = AND(WX2048, RESET)
--	WX2113 = AND(WX2050, RESET)
--	WX2115 = AND(WX2052, RESET)
--	WX2117 = AND(WX2054, RESET)
--	WX2119 = AND(WX2056, RESET)
--	WX2121 = AND(WX2058, RESET)
--	WX2123 = AND(WX2060, RESET)
--	WX2125 = AND(WX2062, RESET)
--	WX2127 = AND(WX2064, RESET)
--	WX2129 = AND(WX2066, RESET)
--	WX2131 = AND(WX2068, RESET)
--	WX2133 = AND(WX2070, RESET)
--	WX2135 = AND(WX2072, RESET)
--	WX2137 = AND(WX2074, RESET)
--	WX2139 = AND(WX2076, RESET)
--	WX2141 = AND(WX2078, RESET)
--	WX2143 = AND(WX2080, RESET)
--	WX2145 = AND(WX2082, RESET)
--	WX2147 = AND(WX2084, RESET)
--	WX2149 = AND(WX2086, RESET)
--	WX2151 = AND(WX2088, RESET)
--	WX2153 = AND(WX2090, RESET)
--	WX2155 = AND(WX2092, RESET)
--	WX2157 = AND(WX2094, RESET)
--	WX2159 = AND(WX2096, RESET)
--	WX2161 = AND(WX2098, RESET)
--	WX2163 = AND(WX2100, RESET)
--	WX2165 = AND(WX2102, RESET)
--	WX2167 = AND(WX2104, RESET)
--	WX2169 = AND(WX2106, RESET)
--	WX2171 = AND(WX2108, RESET)
--	WX2173 = AND(WX2110, RESET)
--	WX2175 = AND(WX2112, RESET)
--	WX2177 = AND(WX2114, RESET)
--	WX2179 = AND(WX2116, RESET)
--	WX2181 = AND(WX2118, RESET)
--	WX2183 = AND(WX2120, RESET)
--	WX2185 = AND(WX2122, RESET)
--	WX2187 = AND(WX2124, RESET)
--	WX2189 = AND(WX2126, RESET)
--	WX2191 = AND(WX2128, RESET)
--	WX2300 = AND(WX2299, WX2298)
--	WX2301 = AND(WX1873, WX2302)
--	WX2307 = AND(WX2306, WX2298)
--	WX2308 = AND(WX1874, WX2309)
--	WX2314 = AND(WX2313, WX2298)
--	WX2315 = AND(WX1875, WX2316)
--	WX2321 = AND(WX2320, WX2298)
--	WX2322 = AND(WX1876, WX2323)
--	WX2328 = AND(WX2327, WX2298)
--	WX2329 = AND(WX1877, WX2330)
--	WX2335 = AND(WX2334, WX2298)
--	WX2336 = AND(WX1878, WX2337)
--	WX2342 = AND(WX2341, WX2298)
--	WX2343 = AND(WX1879, WX2344)
--	WX2349 = AND(WX2348, WX2298)
--	WX2350 = AND(WX1880, WX2351)
--	WX2356 = AND(WX2355, WX2298)
--	WX2357 = AND(WX1881, WX2358)
--	WX2363 = AND(WX2362, WX2298)
--	WX2364 = AND(WX1882, WX2365)
--	WX2370 = AND(WX2369, WX2298)
--	WX2371 = AND(WX1883, WX2372)
--	WX2377 = AND(WX2376, WX2298)
--	WX2378 = AND(WX1884, WX2379)
--	WX2384 = AND(WX2383, WX2298)
--	WX2385 = AND(WX1885, WX2386)
--	WX2391 = AND(WX2390, WX2298)
--	WX2392 = AND(WX1886, WX2393)
--	WX2398 = AND(WX2397, WX2298)
--	WX2399 = AND(WX1887, WX2400)
--	WX2405 = AND(WX2404, WX2298)
--	WX2406 = AND(WX1888, WX2407)
--	WX2412 = AND(WX2411, WX2298)
--	WX2413 = AND(WX1889, WX2414)
--	WX2419 = AND(WX2418, WX2298)
--	WX2420 = AND(WX1890, WX2421)
--	WX2426 = AND(WX2425, WX2298)
--	WX2427 = AND(WX1891, WX2428)
--	WX2433 = AND(WX2432, WX2298)
--	WX2434 = AND(WX1892, WX2435)
--	WX2440 = AND(WX2439, WX2298)
--	WX2441 = AND(WX1893, WX2442)
--	WX2447 = AND(WX2446, WX2298)
--	WX2448 = AND(WX1894, WX2449)
--	WX2454 = AND(WX2453, WX2298)
--	WX2455 = AND(WX1895, WX2456)
--	WX2461 = AND(WX2460, WX2298)
--	WX2462 = AND(WX1896, WX2463)
--	WX2468 = AND(WX2467, WX2298)
--	WX2469 = AND(WX1897, WX2470)
--	WX2475 = AND(WX2474, WX2298)
--	WX2476 = AND(WX1898, WX2477)
--	WX2482 = AND(WX2481, WX2298)
--	WX2483 = AND(WX1899, WX2484)
--	WX2489 = AND(WX2488, WX2298)
--	WX2490 = AND(WX1900, WX2491)
--	WX2496 = AND(WX2495, WX2298)
--	WX2497 = AND(WX1901, WX2498)
--	WX2503 = AND(WX2502, WX2298)
--	WX2504 = AND(WX1902, WX2505)
--	WX2510 = AND(WX2509, WX2298)
--	WX2511 = AND(WX1903, WX2512)
--	WX2517 = AND(WX2516, WX2298)
--	WX2518 = AND(WX1904, WX2519)
--	WX2557 = AND(WX2527, WX2556)
--	WX2559 = AND(WX2555, WX2556)
--	WX2561 = AND(WX2554, WX2556)
--	WX2563 = AND(WX2553, WX2556)
--	WX2565 = AND(WX2526, WX2556)
--	WX2567 = AND(WX2552, WX2556)
--	WX2569 = AND(WX2551, WX2556)
--	WX2571 = AND(WX2550, WX2556)
--	WX2573 = AND(WX2549, WX2556)
--	WX2575 = AND(WX2548, WX2556)
--	WX2577 = AND(WX2547, WX2556)
--	WX2579 = AND(WX2525, WX2556)
--	WX2581 = AND(WX2546, WX2556)
--	WX2583 = AND(WX2545, WX2556)
--	WX2585 = AND(WX2544, WX2556)
--	WX2587 = AND(WX2543, WX2556)
--	WX2589 = AND(WX2524, WX2556)
--	WX2591 = AND(WX2542, WX2556)
--	WX2593 = AND(WX2541, WX2556)
--	WX2595 = AND(WX2540, WX2556)
--	WX2597 = AND(WX2539, WX2556)
--	WX2599 = AND(WX2538, WX2556)
--	WX2601 = AND(WX2537, WX2556)
--	WX2603 = AND(WX2536, WX2556)
--	WX2605 = AND(WX2535, WX2556)
--	WX2607 = AND(WX2534, WX2556)
--	WX2609 = AND(WX2533, WX2556)
--	WX2611 = AND(WX2532, WX2556)
--	WX2613 = AND(WX2531, WX2556)
--	WX2615 = AND(WX2530, WX2556)
--	WX2617 = AND(WX2529, WX2556)
--	WX2619 = AND(WX2528, WX2556)
--	WX2621 = AND(WX2632, WX3589)
--	WX2622 = AND(WX2628, WX2623)
--	WX2625 = AND(CRC_OUT_7_31, WX3590)
--	WX2626 = AND(WX4891, WX2627)
--	WX2629 = AND(WX3071, WX3590)
--	WX2630 = AND(WX3598, WX2631)
--	WX2635 = AND(WX2646, WX3589)
--	WX2636 = AND(WX2642, WX2637)
--	WX2639 = AND(CRC_OUT_7_30, WX3590)
--	WX2640 = AND(WX4898, WX2641)
--	WX2643 = AND(WX3073, WX3590)
--	WX2644 = AND(WX3605, WX2645)
--	WX2649 = AND(WX2660, WX3589)
--	WX2650 = AND(WX2656, WX2651)
--	WX2653 = AND(CRC_OUT_7_29, WX3590)
--	WX2654 = AND(WX4905, WX2655)
--	WX2657 = AND(WX3075, WX3590)
--	WX2658 = AND(WX3612, WX2659)
--	WX2663 = AND(WX2674, WX3589)
--	WX2664 = AND(WX2670, WX2665)
--	WX2667 = AND(CRC_OUT_7_28, WX3590)
--	WX2668 = AND(WX4912, WX2669)
--	WX2671 = AND(WX3077, WX3590)
--	WX2672 = AND(WX3619, WX2673)
--	WX2677 = AND(WX2688, WX3589)
--	WX2678 = AND(WX2684, WX2679)
--	WX2681 = AND(CRC_OUT_7_27, WX3590)
--	WX2682 = AND(WX4919, WX2683)
--	WX2685 = AND(WX3079, WX3590)
--	WX2686 = AND(WX3626, WX2687)
--	WX2691 = AND(WX2702, WX3589)
--	WX2692 = AND(WX2698, WX2693)
--	WX2695 = AND(CRC_OUT_7_26, WX3590)
--	WX2696 = AND(WX4926, WX2697)
--	WX2699 = AND(WX3081, WX3590)
--	WX2700 = AND(WX3633, WX2701)
--	WX2705 = AND(WX2716, WX3589)
--	WX2706 = AND(WX2712, WX2707)
--	WX2709 = AND(CRC_OUT_7_25, WX3590)
--	WX2710 = AND(WX4933, WX2711)
--	WX2713 = AND(WX3083, WX3590)
--	WX2714 = AND(WX3640, WX2715)
--	WX2719 = AND(WX2730, WX3589)
--	WX2720 = AND(WX2726, WX2721)
--	WX2723 = AND(CRC_OUT_7_24, WX3590)
--	WX2724 = AND(WX4940, WX2725)
--	WX2727 = AND(WX3085, WX3590)
--	WX2728 = AND(WX3647, WX2729)
--	WX2733 = AND(WX2744, WX3589)
--	WX2734 = AND(WX2740, WX2735)
--	WX2737 = AND(CRC_OUT_7_23, WX3590)
--	WX2738 = AND(WX4947, WX2739)
--	WX2741 = AND(WX3087, WX3590)
--	WX2742 = AND(WX3654, WX2743)
--	WX2747 = AND(WX2758, WX3589)
--	WX2748 = AND(WX2754, WX2749)
--	WX2751 = AND(CRC_OUT_7_22, WX3590)
--	WX2752 = AND(WX4954, WX2753)
--	WX2755 = AND(WX3089, WX3590)
--	WX2756 = AND(WX3661, WX2757)
--	WX2761 = AND(WX2772, WX3589)
--	WX2762 = AND(WX2768, WX2763)
--	WX2765 = AND(CRC_OUT_7_21, WX3590)
--	WX2766 = AND(WX4961, WX2767)
--	WX2769 = AND(WX3091, WX3590)
--	WX2770 = AND(WX3668, WX2771)
--	WX2775 = AND(WX2786, WX3589)
--	WX2776 = AND(WX2782, WX2777)
--	WX2779 = AND(CRC_OUT_7_20, WX3590)
--	WX2780 = AND(WX4968, WX2781)
--	WX2783 = AND(WX3093, WX3590)
--	WX2784 = AND(WX3675, WX2785)
--	WX2789 = AND(WX2800, WX3589)
--	WX2790 = AND(WX2796, WX2791)
--	WX2793 = AND(CRC_OUT_7_19, WX3590)
--	WX2794 = AND(WX4975, WX2795)
--	WX2797 = AND(WX3095, WX3590)
--	WX2798 = AND(WX3682, WX2799)
--	WX2803 = AND(WX2814, WX3589)
--	WX2804 = AND(WX2810, WX2805)
--	WX2807 = AND(CRC_OUT_7_18, WX3590)
--	WX2808 = AND(WX4982, WX2809)
--	WX2811 = AND(WX3097, WX3590)
--	WX2812 = AND(WX3689, WX2813)
--	WX2817 = AND(WX2828, WX3589)
--	WX2818 = AND(WX2824, WX2819)
--	WX2821 = AND(CRC_OUT_7_17, WX3590)
--	WX2822 = AND(WX4989, WX2823)
--	WX2825 = AND(WX3099, WX3590)
--	WX2826 = AND(WX3696, WX2827)
--	WX2831 = AND(WX2842, WX3589)
--	WX2832 = AND(WX2838, WX2833)
--	WX2835 = AND(CRC_OUT_7_16, WX3590)
--	WX2836 = AND(WX4996, WX2837)
--	WX2839 = AND(WX3101, WX3590)
--	WX2840 = AND(WX3703, WX2841)
--	WX2845 = AND(WX2856, WX3589)
--	WX2846 = AND(WX2852, WX2847)
--	WX2849 = AND(CRC_OUT_7_15, WX3590)
--	WX2850 = AND(WX5003, WX2851)
--	WX2853 = AND(WX3103, WX3590)
--	WX2854 = AND(WX3710, WX2855)
--	WX2859 = AND(WX2870, WX3589)
--	WX2860 = AND(WX2866, WX2861)
--	WX2863 = AND(CRC_OUT_7_14, WX3590)
--	WX2864 = AND(WX5010, WX2865)
--	WX2867 = AND(WX3105, WX3590)
--	WX2868 = AND(WX3717, WX2869)
--	WX2873 = AND(WX2884, WX3589)
--	WX2874 = AND(WX2880, WX2875)
--	WX2877 = AND(CRC_OUT_7_13, WX3590)
--	WX2878 = AND(WX5017, WX2879)
--	WX2881 = AND(WX3107, WX3590)
--	WX2882 = AND(WX3724, WX2883)
--	WX2887 = AND(WX2898, WX3589)
--	WX2888 = AND(WX2894, WX2889)
--	WX2891 = AND(CRC_OUT_7_12, WX3590)
--	WX2892 = AND(WX5024, WX2893)
--	WX2895 = AND(WX3109, WX3590)
--	WX2896 = AND(WX3731, WX2897)
--	WX2901 = AND(WX2912, WX3589)
--	WX2902 = AND(WX2908, WX2903)
--	WX2905 = AND(CRC_OUT_7_11, WX3590)
--	WX2906 = AND(WX5031, WX2907)
--	WX2909 = AND(WX3111, WX3590)
--	WX2910 = AND(WX3738, WX2911)
--	WX2915 = AND(WX2926, WX3589)
--	WX2916 = AND(WX2922, WX2917)
--	WX2919 = AND(CRC_OUT_7_10, WX3590)
--	WX2920 = AND(WX5038, WX2921)
--	WX2923 = AND(WX3113, WX3590)
--	WX2924 = AND(WX3745, WX2925)
--	WX2929 = AND(WX2940, WX3589)
--	WX2930 = AND(WX2936, WX2931)
--	WX2933 = AND(CRC_OUT_7_9, WX3590)
--	WX2934 = AND(WX5045, WX2935)
--	WX2937 = AND(WX3115, WX3590)
--	WX2938 = AND(WX3752, WX2939)
--	WX2943 = AND(WX2954, WX3589)
--	WX2944 = AND(WX2950, WX2945)
--	WX2947 = AND(CRC_OUT_7_8, WX3590)
--	WX2948 = AND(WX5052, WX2949)
--	WX2951 = AND(WX3117, WX3590)
--	WX2952 = AND(WX3759, WX2953)
--	WX2957 = AND(WX2968, WX3589)
--	WX2958 = AND(WX2964, WX2959)
--	WX2961 = AND(CRC_OUT_7_7, WX3590)
--	WX2962 = AND(WX5059, WX2963)
--	WX2965 = AND(WX3119, WX3590)
--	WX2966 = AND(WX3766, WX2967)
--	WX2971 = AND(WX2982, WX3589)
--	WX2972 = AND(WX2978, WX2973)
--	WX2975 = AND(CRC_OUT_7_6, WX3590)
--	WX2976 = AND(WX5066, WX2977)
--	WX2979 = AND(WX3121, WX3590)
--	WX2980 = AND(WX3773, WX2981)
--	WX2985 = AND(WX2996, WX3589)
--	WX2986 = AND(WX2992, WX2987)
--	WX2989 = AND(CRC_OUT_7_5, WX3590)
--	WX2990 = AND(WX5073, WX2991)
--	WX2993 = AND(WX3123, WX3590)
--	WX2994 = AND(WX3780, WX2995)
--	WX2999 = AND(WX3010, WX3589)
--	WX3000 = AND(WX3006, WX3001)
--	WX3003 = AND(CRC_OUT_7_4, WX3590)
--	WX3004 = AND(WX5080, WX3005)
--	WX3007 = AND(WX3125, WX3590)
--	WX3008 = AND(WX3787, WX3009)
--	WX3013 = AND(WX3024, WX3589)
--	WX3014 = AND(WX3020, WX3015)
--	WX3017 = AND(CRC_OUT_7_3, WX3590)
--	WX3018 = AND(WX5087, WX3019)
--	WX3021 = AND(WX3127, WX3590)
--	WX3022 = AND(WX3794, WX3023)
--	WX3027 = AND(WX3038, WX3589)
--	WX3028 = AND(WX3034, WX3029)
--	WX3031 = AND(CRC_OUT_7_2, WX3590)
--	WX3032 = AND(WX5094, WX3033)
--	WX3035 = AND(WX3129, WX3590)
--	WX3036 = AND(WX3801, WX3037)
--	WX3041 = AND(WX3052, WX3589)
--	WX3042 = AND(WX3048, WX3043)
--	WX3045 = AND(CRC_OUT_7_1, WX3590)
--	WX3046 = AND(WX5101, WX3047)
--	WX3049 = AND(WX3131, WX3590)
--	WX3050 = AND(WX3808, WX3051)
--	WX3055 = AND(WX3066, WX3589)
--	WX3056 = AND(WX3062, WX3057)
--	WX3059 = AND(CRC_OUT_7_0, WX3590)
--	WX3060 = AND(WX5108, WX3061)
--	WX3063 = AND(WX3133, WX3590)
--	WX3064 = AND(WX3815, WX3065)
--	WX3070 = AND(WX3073, RESET)
--	WX3072 = AND(WX3075, RESET)
--	WX3074 = AND(WX3077, RESET)
--	WX3076 = AND(WX3079, RESET)
--	WX3078 = AND(WX3081, RESET)
--	WX3080 = AND(WX3083, RESET)
--	WX3082 = AND(WX3085, RESET)
--	WX3084 = AND(WX3087, RESET)
--	WX3086 = AND(WX3089, RESET)
--	WX3088 = AND(WX3091, RESET)
--	WX3090 = AND(WX3093, RESET)
--	WX3092 = AND(WX3095, RESET)
--	WX3094 = AND(WX3097, RESET)
--	WX3096 = AND(WX3099, RESET)
--	WX3098 = AND(WX3101, RESET)
--	WX3100 = AND(WX3103, RESET)
--	WX3102 = AND(WX3105, RESET)
--	WX3104 = AND(WX3107, RESET)
--	WX3106 = AND(WX3109, RESET)
--	WX3108 = AND(WX3111, RESET)
--	WX3110 = AND(WX3113, RESET)
--	WX3112 = AND(WX3115, RESET)
--	WX3114 = AND(WX3117, RESET)
--	WX3116 = AND(WX3119, RESET)
--	WX3118 = AND(WX3121, RESET)
--	WX3120 = AND(WX3123, RESET)
--	WX3122 = AND(WX3125, RESET)
--	WX3124 = AND(WX3127, RESET)
--	WX3126 = AND(WX3129, RESET)
--	WX3128 = AND(WX3131, RESET)
--	WX3130 = AND(WX3133, RESET)
--	WX3132 = AND(WX3069, RESET)
--	WX3230 = AND(WX2634, RESET)
--	WX3232 = AND(WX2648, RESET)
--	WX3234 = AND(WX2662, RESET)
--	WX3236 = AND(WX2676, RESET)
--	WX3238 = AND(WX2690, RESET)
--	WX3240 = AND(WX2704, RESET)
--	WX3242 = AND(WX2718, RESET)
--	WX3244 = AND(WX2732, RESET)
--	WX3246 = AND(WX2746, RESET)
--	WX3248 = AND(WX2760, RESET)
--	WX3250 = AND(WX2774, RESET)
--	WX3252 = AND(WX2788, RESET)
--	WX3254 = AND(WX2802, RESET)
--	WX3256 = AND(WX2816, RESET)
--	WX3258 = AND(WX2830, RESET)
--	WX3260 = AND(WX2844, RESET)
--	WX3262 = AND(WX2858, RESET)
--	WX3264 = AND(WX2872, RESET)
--	WX3266 = AND(WX2886, RESET)
--	WX3268 = AND(WX2900, RESET)
--	WX3270 = AND(WX2914, RESET)
--	WX3272 = AND(WX2928, RESET)
--	WX3274 = AND(WX2942, RESET)
--	WX3276 = AND(WX2956, RESET)
--	WX3278 = AND(WX2970, RESET)
--	WX3280 = AND(WX2984, RESET)
--	WX3282 = AND(WX2998, RESET)
--	WX3284 = AND(WX3012, RESET)
--	WX3286 = AND(WX3026, RESET)
--	WX3288 = AND(WX3040, RESET)
--	WX3290 = AND(WX3054, RESET)
--	WX3292 = AND(WX3068, RESET)
--	WX3294 = AND(WX3231, RESET)
--	WX3296 = AND(WX3233, RESET)
--	WX3298 = AND(WX3235, RESET)
--	WX3300 = AND(WX3237, RESET)
--	WX3302 = AND(WX3239, RESET)
--	WX3304 = AND(WX3241, RESET)
--	WX3306 = AND(WX3243, RESET)
--	WX3308 = AND(WX3245, RESET)
--	WX3310 = AND(WX3247, RESET)
--	WX3312 = AND(WX3249, RESET)
--	WX3314 = AND(WX3251, RESET)
--	WX3316 = AND(WX3253, RESET)
--	WX3318 = AND(WX3255, RESET)
--	WX3320 = AND(WX3257, RESET)
--	WX3322 = AND(WX3259, RESET)
--	WX3324 = AND(WX3261, RESET)
--	WX3326 = AND(WX3263, RESET)
--	WX3328 = AND(WX3265, RESET)
--	WX3330 = AND(WX3267, RESET)
--	WX3332 = AND(WX3269, RESET)
--	WX3334 = AND(WX3271, RESET)
--	WX3336 = AND(WX3273, RESET)
--	WX3338 = AND(WX3275, RESET)
--	WX3340 = AND(WX3277, RESET)
--	WX3342 = AND(WX3279, RESET)
--	WX3344 = AND(WX3281, RESET)
--	WX3346 = AND(WX3283, RESET)
--	WX3348 = AND(WX3285, RESET)
--	WX3350 = AND(WX3287, RESET)
--	WX3352 = AND(WX3289, RESET)
--	WX3354 = AND(WX3291, RESET)
--	WX3356 = AND(WX3293, RESET)
--	WX3358 = AND(WX3295, RESET)
--	WX3360 = AND(WX3297, RESET)
--	WX3362 = AND(WX3299, RESET)
--	WX3364 = AND(WX3301, RESET)
--	WX3366 = AND(WX3303, RESET)
--	WX3368 = AND(WX3305, RESET)
--	WX3370 = AND(WX3307, RESET)
--	WX3372 = AND(WX3309, RESET)
--	WX3374 = AND(WX3311, RESET)
--	WX3376 = AND(WX3313, RESET)
--	WX3378 = AND(WX3315, RESET)
--	WX3380 = AND(WX3317, RESET)
--	WX3382 = AND(WX3319, RESET)
--	WX3384 = AND(WX3321, RESET)
--	WX3386 = AND(WX3323, RESET)
--	WX3388 = AND(WX3325, RESET)
--	WX3390 = AND(WX3327, RESET)
--	WX3392 = AND(WX3329, RESET)
--	WX3394 = AND(WX3331, RESET)
--	WX3396 = AND(WX3333, RESET)
--	WX3398 = AND(WX3335, RESET)
--	WX3400 = AND(WX3337, RESET)
--	WX3402 = AND(WX3339, RESET)
--	WX3404 = AND(WX3341, RESET)
--	WX3406 = AND(WX3343, RESET)
--	WX3408 = AND(WX3345, RESET)
--	WX3410 = AND(WX3347, RESET)
--	WX3412 = AND(WX3349, RESET)
--	WX3414 = AND(WX3351, RESET)
--	WX3416 = AND(WX3353, RESET)
--	WX3418 = AND(WX3355, RESET)
--	WX3420 = AND(WX3357, RESET)
--	WX3422 = AND(WX3359, RESET)
--	WX3424 = AND(WX3361, RESET)
--	WX3426 = AND(WX3363, RESET)
--	WX3428 = AND(WX3365, RESET)
--	WX3430 = AND(WX3367, RESET)
--	WX3432 = AND(WX3369, RESET)
--	WX3434 = AND(WX3371, RESET)
--	WX3436 = AND(WX3373, RESET)
--	WX3438 = AND(WX3375, RESET)
--	WX3440 = AND(WX3377, RESET)
--	WX3442 = AND(WX3379, RESET)
--	WX3444 = AND(WX3381, RESET)
--	WX3446 = AND(WX3383, RESET)
--	WX3448 = AND(WX3385, RESET)
--	WX3450 = AND(WX3387, RESET)
--	WX3452 = AND(WX3389, RESET)
--	WX3454 = AND(WX3391, RESET)
--	WX3456 = AND(WX3393, RESET)
--	WX3458 = AND(WX3395, RESET)
--	WX3460 = AND(WX3397, RESET)
--	WX3462 = AND(WX3399, RESET)
--	WX3464 = AND(WX3401, RESET)
--	WX3466 = AND(WX3403, RESET)
--	WX3468 = AND(WX3405, RESET)
--	WX3470 = AND(WX3407, RESET)
--	WX3472 = AND(WX3409, RESET)
--	WX3474 = AND(WX3411, RESET)
--	WX3476 = AND(WX3413, RESET)
--	WX3478 = AND(WX3415, RESET)
--	WX3480 = AND(WX3417, RESET)
--	WX3482 = AND(WX3419, RESET)
--	WX3484 = AND(WX3421, RESET)
--	WX3593 = AND(WX3592, WX3591)
--	WX3594 = AND(WX3166, WX3595)
--	WX3600 = AND(WX3599, WX3591)
--	WX3601 = AND(WX3167, WX3602)
--	WX3607 = AND(WX3606, WX3591)
--	WX3608 = AND(WX3168, WX3609)
--	WX3614 = AND(WX3613, WX3591)
--	WX3615 = AND(WX3169, WX3616)
--	WX3621 = AND(WX3620, WX3591)
--	WX3622 = AND(WX3170, WX3623)
--	WX3628 = AND(WX3627, WX3591)
--	WX3629 = AND(WX3171, WX3630)
--	WX3635 = AND(WX3634, WX3591)
--	WX3636 = AND(WX3172, WX3637)
--	WX3642 = AND(WX3641, WX3591)
--	WX3643 = AND(WX3173, WX3644)
--	WX3649 = AND(WX3648, WX3591)
--	WX3650 = AND(WX3174, WX3651)
--	WX3656 = AND(WX3655, WX3591)
--	WX3657 = AND(WX3175, WX3658)
--	WX3663 = AND(WX3662, WX3591)
--	WX3664 = AND(WX3176, WX3665)
--	WX3670 = AND(WX3669, WX3591)
--	WX3671 = AND(WX3177, WX3672)
--	WX3677 = AND(WX3676, WX3591)
--	WX3678 = AND(WX3178, WX3679)
--	WX3684 = AND(WX3683, WX3591)
--	WX3685 = AND(WX3179, WX3686)
--	WX3691 = AND(WX3690, WX3591)
--	WX3692 = AND(WX3180, WX3693)
--	WX3698 = AND(WX3697, WX3591)
--	WX3699 = AND(WX3181, WX3700)
--	WX3705 = AND(WX3704, WX3591)
--	WX3706 = AND(WX3182, WX3707)
--	WX3712 = AND(WX3711, WX3591)
--	WX3713 = AND(WX3183, WX3714)
--	WX3719 = AND(WX3718, WX3591)
--	WX3720 = AND(WX3184, WX3721)
--	WX3726 = AND(WX3725, WX3591)
--	WX3727 = AND(WX3185, WX3728)
--	WX3733 = AND(WX3732, WX3591)
--	WX3734 = AND(WX3186, WX3735)
--	WX3740 = AND(WX3739, WX3591)
--	WX3741 = AND(WX3187, WX3742)
--	WX3747 = AND(WX3746, WX3591)
--	WX3748 = AND(WX3188, WX3749)
--	WX3754 = AND(WX3753, WX3591)
--	WX3755 = AND(WX3189, WX3756)
--	WX3761 = AND(WX3760, WX3591)
--	WX3762 = AND(WX3190, WX3763)
--	WX3768 = AND(WX3767, WX3591)
--	WX3769 = AND(WX3191, WX3770)
--	WX3775 = AND(WX3774, WX3591)
--	WX3776 = AND(WX3192, WX3777)
--	WX3782 = AND(WX3781, WX3591)
--	WX3783 = AND(WX3193, WX3784)
--	WX3789 = AND(WX3788, WX3591)
--	WX3790 = AND(WX3194, WX3791)
--	WX3796 = AND(WX3795, WX3591)
--	WX3797 = AND(WX3195, WX3798)
--	WX3803 = AND(WX3802, WX3591)
--	WX3804 = AND(WX3196, WX3805)
--	WX3810 = AND(WX3809, WX3591)
--	WX3811 = AND(WX3197, WX3812)
--	WX3850 = AND(WX3820, WX3849)
--	WX3852 = AND(WX3848, WX3849)
--	WX3854 = AND(WX3847, WX3849)
--	WX3856 = AND(WX3846, WX3849)
--	WX3858 = AND(WX3819, WX3849)
--	WX3860 = AND(WX3845, WX3849)
--	WX3862 = AND(WX3844, WX3849)
--	WX3864 = AND(WX3843, WX3849)
--	WX3866 = AND(WX3842, WX3849)
--	WX3868 = AND(WX3841, WX3849)
--	WX3870 = AND(WX3840, WX3849)
--	WX3872 = AND(WX3818, WX3849)
--	WX3874 = AND(WX3839, WX3849)
--	WX3876 = AND(WX3838, WX3849)
--	WX3878 = AND(WX3837, WX3849)
--	WX3880 = AND(WX3836, WX3849)
--	WX3882 = AND(WX3817, WX3849)
--	WX3884 = AND(WX3835, WX3849)
--	WX3886 = AND(WX3834, WX3849)
--	WX3888 = AND(WX3833, WX3849)
--	WX3890 = AND(WX3832, WX3849)
--	WX3892 = AND(WX3831, WX3849)
--	WX3894 = AND(WX3830, WX3849)
--	WX3896 = AND(WX3829, WX3849)
--	WX3898 = AND(WX3828, WX3849)
--	WX3900 = AND(WX3827, WX3849)
--	WX3902 = AND(WX3826, WX3849)
--	WX3904 = AND(WX3825, WX3849)
--	WX3906 = AND(WX3824, WX3849)
--	WX3908 = AND(WX3823, WX3849)
--	WX3910 = AND(WX3822, WX3849)
--	WX3912 = AND(WX3821, WX3849)
--	WX3914 = AND(WX3925, WX4882)
--	WX3915 = AND(WX3921, WX3916)
--	WX3918 = AND(CRC_OUT_6_31, WX4883)
--	WX3919 = AND(WX6184, WX3920)
--	WX3922 = AND(WX4364, WX4883)
--	WX3923 = AND(WX4891, WX3924)
--	WX3928 = AND(WX3939, WX4882)
--	WX3929 = AND(WX3935, WX3930)
--	WX3932 = AND(CRC_OUT_6_30, WX4883)
--	WX3933 = AND(WX6191, WX3934)
--	WX3936 = AND(WX4366, WX4883)
--	WX3937 = AND(WX4898, WX3938)
--	WX3942 = AND(WX3953, WX4882)
--	WX3943 = AND(WX3949, WX3944)
--	WX3946 = AND(CRC_OUT_6_29, WX4883)
--	WX3947 = AND(WX6198, WX3948)
--	WX3950 = AND(WX4368, WX4883)
--	WX3951 = AND(WX4905, WX3952)
--	WX3956 = AND(WX3967, WX4882)
--	WX3957 = AND(WX3963, WX3958)
--	WX3960 = AND(CRC_OUT_6_28, WX4883)
--	WX3961 = AND(WX6205, WX3962)
--	WX3964 = AND(WX4370, WX4883)
--	WX3965 = AND(WX4912, WX3966)
--	WX3970 = AND(WX3981, WX4882)
--	WX3971 = AND(WX3977, WX3972)
--	WX3974 = AND(CRC_OUT_6_27, WX4883)
--	WX3975 = AND(WX6212, WX3976)
--	WX3978 = AND(WX4372, WX4883)
--	WX3979 = AND(WX4919, WX3980)
--	WX3984 = AND(WX3995, WX4882)
--	WX3985 = AND(WX3991, WX3986)
--	WX3988 = AND(CRC_OUT_6_26, WX4883)
--	WX3989 = AND(WX6219, WX3990)
--	WX3992 = AND(WX4374, WX4883)
--	WX3993 = AND(WX4926, WX3994)
--	WX3998 = AND(WX4009, WX4882)
--	WX3999 = AND(WX4005, WX4000)
--	WX4002 = AND(CRC_OUT_6_25, WX4883)
--	WX4003 = AND(WX6226, WX4004)
--	WX4006 = AND(WX4376, WX4883)
--	WX4007 = AND(WX4933, WX4008)
--	WX4012 = AND(WX4023, WX4882)
--	WX4013 = AND(WX4019, WX4014)
--	WX4016 = AND(CRC_OUT_6_24, WX4883)
--	WX4017 = AND(WX6233, WX4018)
--	WX4020 = AND(WX4378, WX4883)
--	WX4021 = AND(WX4940, WX4022)
--	WX4026 = AND(WX4037, WX4882)
--	WX4027 = AND(WX4033, WX4028)
--	WX4030 = AND(CRC_OUT_6_23, WX4883)
--	WX4031 = AND(WX6240, WX4032)
--	WX4034 = AND(WX4380, WX4883)
--	WX4035 = AND(WX4947, WX4036)
--	WX4040 = AND(WX4051, WX4882)
--	WX4041 = AND(WX4047, WX4042)
--	WX4044 = AND(CRC_OUT_6_22, WX4883)
--	WX4045 = AND(WX6247, WX4046)
--	WX4048 = AND(WX4382, WX4883)
--	WX4049 = AND(WX4954, WX4050)
--	WX4054 = AND(WX4065, WX4882)
--	WX4055 = AND(WX4061, WX4056)
--	WX4058 = AND(CRC_OUT_6_21, WX4883)
--	WX4059 = AND(WX6254, WX4060)
--	WX4062 = AND(WX4384, WX4883)
--	WX4063 = AND(WX4961, WX4064)
--	WX4068 = AND(WX4079, WX4882)
--	WX4069 = AND(WX4075, WX4070)
--	WX4072 = AND(CRC_OUT_6_20, WX4883)
--	WX4073 = AND(WX6261, WX4074)
--	WX4076 = AND(WX4386, WX4883)
--	WX4077 = AND(WX4968, WX4078)
--	WX4082 = AND(WX4093, WX4882)
--	WX4083 = AND(WX4089, WX4084)
--	WX4086 = AND(CRC_OUT_6_19, WX4883)
--	WX4087 = AND(WX6268, WX4088)
--	WX4090 = AND(WX4388, WX4883)
--	WX4091 = AND(WX4975, WX4092)
--	WX4096 = AND(WX4107, WX4882)
--	WX4097 = AND(WX4103, WX4098)
--	WX4100 = AND(CRC_OUT_6_18, WX4883)
--	WX4101 = AND(WX6275, WX4102)
--	WX4104 = AND(WX4390, WX4883)
--	WX4105 = AND(WX4982, WX4106)
--	WX4110 = AND(WX4121, WX4882)
--	WX4111 = AND(WX4117, WX4112)
--	WX4114 = AND(CRC_OUT_6_17, WX4883)
--	WX4115 = AND(WX6282, WX4116)
--	WX4118 = AND(WX4392, WX4883)
--	WX4119 = AND(WX4989, WX4120)
--	WX4124 = AND(WX4135, WX4882)
--	WX4125 = AND(WX4131, WX4126)
--	WX4128 = AND(CRC_OUT_6_16, WX4883)
--	WX4129 = AND(WX6289, WX4130)
--	WX4132 = AND(WX4394, WX4883)
--	WX4133 = AND(WX4996, WX4134)
--	WX4138 = AND(WX4149, WX4882)
--	WX4139 = AND(WX4145, WX4140)
--	WX4142 = AND(CRC_OUT_6_15, WX4883)
--	WX4143 = AND(WX6296, WX4144)
--	WX4146 = AND(WX4396, WX4883)
--	WX4147 = AND(WX5003, WX4148)
--	WX4152 = AND(WX4163, WX4882)
--	WX4153 = AND(WX4159, WX4154)
--	WX4156 = AND(CRC_OUT_6_14, WX4883)
--	WX4157 = AND(WX6303, WX4158)
--	WX4160 = AND(WX4398, WX4883)
--	WX4161 = AND(WX5010, WX4162)
--	WX4166 = AND(WX4177, WX4882)
--	WX4167 = AND(WX4173, WX4168)
--	WX4170 = AND(CRC_OUT_6_13, WX4883)
--	WX4171 = AND(WX6310, WX4172)
--	WX4174 = AND(WX4400, WX4883)
--	WX4175 = AND(WX5017, WX4176)
--	WX4180 = AND(WX4191, WX4882)
--	WX4181 = AND(WX4187, WX4182)
--	WX4184 = AND(CRC_OUT_6_12, WX4883)
--	WX4185 = AND(WX6317, WX4186)
--	WX4188 = AND(WX4402, WX4883)
--	WX4189 = AND(WX5024, WX4190)
--	WX4194 = AND(WX4205, WX4882)
--	WX4195 = AND(WX4201, WX4196)
--	WX4198 = AND(CRC_OUT_6_11, WX4883)
--	WX4199 = AND(WX6324, WX4200)
--	WX4202 = AND(WX4404, WX4883)
--	WX4203 = AND(WX5031, WX4204)
--	WX4208 = AND(WX4219, WX4882)
--	WX4209 = AND(WX4215, WX4210)
--	WX4212 = AND(CRC_OUT_6_10, WX4883)
--	WX4213 = AND(WX6331, WX4214)
--	WX4216 = AND(WX4406, WX4883)
--	WX4217 = AND(WX5038, WX4218)
--	WX4222 = AND(WX4233, WX4882)
--	WX4223 = AND(WX4229, WX4224)
--	WX4226 = AND(CRC_OUT_6_9, WX4883)
--	WX4227 = AND(WX6338, WX4228)
--	WX4230 = AND(WX4408, WX4883)
--	WX4231 = AND(WX5045, WX4232)
--	WX4236 = AND(WX4247, WX4882)
--	WX4237 = AND(WX4243, WX4238)
--	WX4240 = AND(CRC_OUT_6_8, WX4883)
--	WX4241 = AND(WX6345, WX4242)
--	WX4244 = AND(WX4410, WX4883)
--	WX4245 = AND(WX5052, WX4246)
--	WX4250 = AND(WX4261, WX4882)
--	WX4251 = AND(WX4257, WX4252)
--	WX4254 = AND(CRC_OUT_6_7, WX4883)
--	WX4255 = AND(WX6352, WX4256)
--	WX4258 = AND(WX4412, WX4883)
--	WX4259 = AND(WX5059, WX4260)
--	WX4264 = AND(WX4275, WX4882)
--	WX4265 = AND(WX4271, WX4266)
--	WX4268 = AND(CRC_OUT_6_6, WX4883)
--	WX4269 = AND(WX6359, WX4270)
--	WX4272 = AND(WX4414, WX4883)
--	WX4273 = AND(WX5066, WX4274)
--	WX4278 = AND(WX4289, WX4882)
--	WX4279 = AND(WX4285, WX4280)
--	WX4282 = AND(CRC_OUT_6_5, WX4883)
--	WX4283 = AND(WX6366, WX4284)
--	WX4286 = AND(WX4416, WX4883)
--	WX4287 = AND(WX5073, WX4288)
--	WX4292 = AND(WX4303, WX4882)
--	WX4293 = AND(WX4299, WX4294)
--	WX4296 = AND(CRC_OUT_6_4, WX4883)
--	WX4297 = AND(WX6373, WX4298)
--	WX4300 = AND(WX4418, WX4883)
--	WX4301 = AND(WX5080, WX4302)
--	WX4306 = AND(WX4317, WX4882)
--	WX4307 = AND(WX4313, WX4308)
--	WX4310 = AND(CRC_OUT_6_3, WX4883)
--	WX4311 = AND(WX6380, WX4312)
--	WX4314 = AND(WX4420, WX4883)
--	WX4315 = AND(WX5087, WX4316)
--	WX4320 = AND(WX4331, WX4882)
--	WX4321 = AND(WX4327, WX4322)
--	WX4324 = AND(CRC_OUT_6_2, WX4883)
--	WX4325 = AND(WX6387, WX4326)
--	WX4328 = AND(WX4422, WX4883)
--	WX4329 = AND(WX5094, WX4330)
--	WX4334 = AND(WX4345, WX4882)
--	WX4335 = AND(WX4341, WX4336)
--	WX4338 = AND(CRC_OUT_6_1, WX4883)
--	WX4339 = AND(WX6394, WX4340)
--	WX4342 = AND(WX4424, WX4883)
--	WX4343 = AND(WX5101, WX4344)
--	WX4348 = AND(WX4359, WX4882)
--	WX4349 = AND(WX4355, WX4350)
--	WX4352 = AND(CRC_OUT_6_0, WX4883)
--	WX4353 = AND(WX6401, WX4354)
--	WX4356 = AND(WX4426, WX4883)
--	WX4357 = AND(WX5108, WX4358)
--	WX4363 = AND(WX4366, RESET)
--	WX4365 = AND(WX4368, RESET)
--	WX4367 = AND(WX4370, RESET)
--	WX4369 = AND(WX4372, RESET)
--	WX4371 = AND(WX4374, RESET)
--	WX4373 = AND(WX4376, RESET)
--	WX4375 = AND(WX4378, RESET)
--	WX4377 = AND(WX4380, RESET)
--	WX4379 = AND(WX4382, RESET)
--	WX4381 = AND(WX4384, RESET)
--	WX4383 = AND(WX4386, RESET)
--	WX4385 = AND(WX4388, RESET)
--	WX4387 = AND(WX4390, RESET)
--	WX4389 = AND(WX4392, RESET)
--	WX4391 = AND(WX4394, RESET)
--	WX4393 = AND(WX4396, RESET)
--	WX4395 = AND(WX4398, RESET)
--	WX4397 = AND(WX4400, RESET)
--	WX4399 = AND(WX4402, RESET)
--	WX4401 = AND(WX4404, RESET)
--	WX4403 = AND(WX4406, RESET)
--	WX4405 = AND(WX4408, RESET)
--	WX4407 = AND(WX4410, RESET)
--	WX4409 = AND(WX4412, RESET)
--	WX4411 = AND(WX4414, RESET)
--	WX4413 = AND(WX4416, RESET)
--	WX4415 = AND(WX4418, RESET)
--	WX4417 = AND(WX4420, RESET)
--	WX4419 = AND(WX4422, RESET)
--	WX4421 = AND(WX4424, RESET)
--	WX4423 = AND(WX4426, RESET)
--	WX4425 = AND(WX4362, RESET)
--	WX4523 = AND(WX3927, RESET)
--	WX4525 = AND(WX3941, RESET)
--	WX4527 = AND(WX3955, RESET)
--	WX4529 = AND(WX3969, RESET)
--	WX4531 = AND(WX3983, RESET)
--	WX4533 = AND(WX3997, RESET)
--	WX4535 = AND(WX4011, RESET)
--	WX4537 = AND(WX4025, RESET)
--	WX4539 = AND(WX4039, RESET)
--	WX4541 = AND(WX4053, RESET)
--	WX4543 = AND(WX4067, RESET)
--	WX4545 = AND(WX4081, RESET)
--	WX4547 = AND(WX4095, RESET)
--	WX4549 = AND(WX4109, RESET)
--	WX4551 = AND(WX4123, RESET)
--	WX4553 = AND(WX4137, RESET)
--	WX4555 = AND(WX4151, RESET)
--	WX4557 = AND(WX4165, RESET)
--	WX4559 = AND(WX4179, RESET)
--	WX4561 = AND(WX4193, RESET)
--	WX4563 = AND(WX4207, RESET)
--	WX4565 = AND(WX4221, RESET)
--	WX4567 = AND(WX4235, RESET)
--	WX4569 = AND(WX4249, RESET)
--	WX4571 = AND(WX4263, RESET)
--	WX4573 = AND(WX4277, RESET)
--	WX4575 = AND(WX4291, RESET)
--	WX4577 = AND(WX4305, RESET)
--	WX4579 = AND(WX4319, RESET)
--	WX4581 = AND(WX4333, RESET)
--	WX4583 = AND(WX4347, RESET)
--	WX4585 = AND(WX4361, RESET)
--	WX4587 = AND(WX4524, RESET)
--	WX4589 = AND(WX4526, RESET)
--	WX4591 = AND(WX4528, RESET)
--	WX4593 = AND(WX4530, RESET)
--	WX4595 = AND(WX4532, RESET)
--	WX4597 = AND(WX4534, RESET)
--	WX4599 = AND(WX4536, RESET)
--	WX4601 = AND(WX4538, RESET)
--	WX4603 = AND(WX4540, RESET)
--	WX4605 = AND(WX4542, RESET)
--	WX4607 = AND(WX4544, RESET)
--	WX4609 = AND(WX4546, RESET)
--	WX4611 = AND(WX4548, RESET)
--	WX4613 = AND(WX4550, RESET)
--	WX4615 = AND(WX4552, RESET)
--	WX4617 = AND(WX4554, RESET)
--	WX4619 = AND(WX4556, RESET)
--	WX4621 = AND(WX4558, RESET)
--	WX4623 = AND(WX4560, RESET)
--	WX4625 = AND(WX4562, RESET)
--	WX4627 = AND(WX4564, RESET)
--	WX4629 = AND(WX4566, RESET)
--	WX4631 = AND(WX4568, RESET)
--	WX4633 = AND(WX4570, RESET)
--	WX4635 = AND(WX4572, RESET)
--	WX4637 = AND(WX4574, RESET)
--	WX4639 = AND(WX4576, RESET)
--	WX4641 = AND(WX4578, RESET)
--	WX4643 = AND(WX4580, RESET)
--	WX4645 = AND(WX4582, RESET)
--	WX4647 = AND(WX4584, RESET)
--	WX4649 = AND(WX4586, RESET)
--	WX4651 = AND(WX4588, RESET)
--	WX4653 = AND(WX4590, RESET)
--	WX4655 = AND(WX4592, RESET)
--	WX4657 = AND(WX4594, RESET)
--	WX4659 = AND(WX4596, RESET)
--	WX4661 = AND(WX4598, RESET)
--	WX4663 = AND(WX4600, RESET)
--	WX4665 = AND(WX4602, RESET)
--	WX4667 = AND(WX4604, RESET)
--	WX4669 = AND(WX4606, RESET)
--	WX4671 = AND(WX4608, RESET)
--	WX4673 = AND(WX4610, RESET)
--	WX4675 = AND(WX4612, RESET)
--	WX4677 = AND(WX4614, RESET)
--	WX4679 = AND(WX4616, RESET)
--	WX4681 = AND(WX4618, RESET)
--	WX4683 = AND(WX4620, RESET)
--	WX4685 = AND(WX4622, RESET)
--	WX4687 = AND(WX4624, RESET)
--	WX4689 = AND(WX4626, RESET)
--	WX4691 = AND(WX4628, RESET)
--	WX4693 = AND(WX4630, RESET)
--	WX4695 = AND(WX4632, RESET)
--	WX4697 = AND(WX4634, RESET)
--	WX4699 = AND(WX4636, RESET)
--	WX4701 = AND(WX4638, RESET)
--	WX4703 = AND(WX4640, RESET)
--	WX4705 = AND(WX4642, RESET)
--	WX4707 = AND(WX4644, RESET)
--	WX4709 = AND(WX4646, RESET)
--	WX4711 = AND(WX4648, RESET)
--	WX4713 = AND(WX4650, RESET)
--	WX4715 = AND(WX4652, RESET)
--	WX4717 = AND(WX4654, RESET)
--	WX4719 = AND(WX4656, RESET)
--	WX4721 = AND(WX4658, RESET)
--	WX4723 = AND(WX4660, RESET)
--	WX4725 = AND(WX4662, RESET)
--	WX4727 = AND(WX4664, RESET)
--	WX4729 = AND(WX4666, RESET)
--	WX4731 = AND(WX4668, RESET)
--	WX4733 = AND(WX4670, RESET)
--	WX4735 = AND(WX4672, RESET)
--	WX4737 = AND(WX4674, RESET)
--	WX4739 = AND(WX4676, RESET)
--	WX4741 = AND(WX4678, RESET)
--	WX4743 = AND(WX4680, RESET)
--	WX4745 = AND(WX4682, RESET)
--	WX4747 = AND(WX4684, RESET)
--	WX4749 = AND(WX4686, RESET)
--	WX4751 = AND(WX4688, RESET)
--	WX4753 = AND(WX4690, RESET)
--	WX4755 = AND(WX4692, RESET)
--	WX4757 = AND(WX4694, RESET)
--	WX4759 = AND(WX4696, RESET)
--	WX4761 = AND(WX4698, RESET)
--	WX4763 = AND(WX4700, RESET)
--	WX4765 = AND(WX4702, RESET)
--	WX4767 = AND(WX4704, RESET)
--	WX4769 = AND(WX4706, RESET)
--	WX4771 = AND(WX4708, RESET)
--	WX4773 = AND(WX4710, RESET)
--	WX4775 = AND(WX4712, RESET)
--	WX4777 = AND(WX4714, RESET)
--	WX4886 = AND(WX4885, WX4884)
--	WX4887 = AND(WX4459, WX4888)
--	WX4893 = AND(WX4892, WX4884)
--	WX4894 = AND(WX4460, WX4895)
--	WX4900 = AND(WX4899, WX4884)
--	WX4901 = AND(WX4461, WX4902)
--	WX4907 = AND(WX4906, WX4884)
--	WX4908 = AND(WX4462, WX4909)
--	WX4914 = AND(WX4913, WX4884)
--	WX4915 = AND(WX4463, WX4916)
--	WX4921 = AND(WX4920, WX4884)
--	WX4922 = AND(WX4464, WX4923)
--	WX4928 = AND(WX4927, WX4884)
--	WX4929 = AND(WX4465, WX4930)
--	WX4935 = AND(WX4934, WX4884)
--	WX4936 = AND(WX4466, WX4937)
--	WX4942 = AND(WX4941, WX4884)
--	WX4943 = AND(WX4467, WX4944)
--	WX4949 = AND(WX4948, WX4884)
--	WX4950 = AND(WX4468, WX4951)
--	WX4956 = AND(WX4955, WX4884)
--	WX4957 = AND(WX4469, WX4958)
--	WX4963 = AND(WX4962, WX4884)
--	WX4964 = AND(WX4470, WX4965)
--	WX4970 = AND(WX4969, WX4884)
--	WX4971 = AND(WX4471, WX4972)
--	WX4977 = AND(WX4976, WX4884)
--	WX4978 = AND(WX4472, WX4979)
--	WX4984 = AND(WX4983, WX4884)
--	WX4985 = AND(WX4473, WX4986)
--	WX4991 = AND(WX4990, WX4884)
--	WX4992 = AND(WX4474, WX4993)
--	WX4998 = AND(WX4997, WX4884)
--	WX4999 = AND(WX4475, WX5000)
--	WX5005 = AND(WX5004, WX4884)
--	WX5006 = AND(WX4476, WX5007)
--	WX5012 = AND(WX5011, WX4884)
--	WX5013 = AND(WX4477, WX5014)
--	WX5019 = AND(WX5018, WX4884)
--	WX5020 = AND(WX4478, WX5021)
--	WX5026 = AND(WX5025, WX4884)
--	WX5027 = AND(WX4479, WX5028)
--	WX5033 = AND(WX5032, WX4884)
--	WX5034 = AND(WX4480, WX5035)
--	WX5040 = AND(WX5039, WX4884)
--	WX5041 = AND(WX4481, WX5042)
--	WX5047 = AND(WX5046, WX4884)
--	WX5048 = AND(WX4482, WX5049)
--	WX5054 = AND(WX5053, WX4884)
--	WX5055 = AND(WX4483, WX5056)
--	WX5061 = AND(WX5060, WX4884)
--	WX5062 = AND(WX4484, WX5063)
--	WX5068 = AND(WX5067, WX4884)
--	WX5069 = AND(WX4485, WX5070)
--	WX5075 = AND(WX5074, WX4884)
--	WX5076 = AND(WX4486, WX5077)
--	WX5082 = AND(WX5081, WX4884)
--	WX5083 = AND(WX4487, WX5084)
--	WX5089 = AND(WX5088, WX4884)
--	WX5090 = AND(WX4488, WX5091)
--	WX5096 = AND(WX5095, WX4884)
--	WX5097 = AND(WX4489, WX5098)
--	WX5103 = AND(WX5102, WX4884)
--	WX5104 = AND(WX4490, WX5105)
--	WX5143 = AND(WX5113, WX5142)
--	WX5145 = AND(WX5141, WX5142)
--	WX5147 = AND(WX5140, WX5142)
--	WX5149 = AND(WX5139, WX5142)
--	WX5151 = AND(WX5112, WX5142)
--	WX5153 = AND(WX5138, WX5142)
--	WX5155 = AND(WX5137, WX5142)
--	WX5157 = AND(WX5136, WX5142)
--	WX5159 = AND(WX5135, WX5142)
--	WX5161 = AND(WX5134, WX5142)
--	WX5163 = AND(WX5133, WX5142)
--	WX5165 = AND(WX5111, WX5142)
--	WX5167 = AND(WX5132, WX5142)
--	WX5169 = AND(WX5131, WX5142)
--	WX5171 = AND(WX5130, WX5142)
--	WX5173 = AND(WX5129, WX5142)
--	WX5175 = AND(WX5110, WX5142)
--	WX5177 = AND(WX5128, WX5142)
--	WX5179 = AND(WX5127, WX5142)
--	WX5181 = AND(WX5126, WX5142)
--	WX5183 = AND(WX5125, WX5142)
--	WX5185 = AND(WX5124, WX5142)
--	WX5187 = AND(WX5123, WX5142)
--	WX5189 = AND(WX5122, WX5142)
--	WX5191 = AND(WX5121, WX5142)
--	WX5193 = AND(WX5120, WX5142)
--	WX5195 = AND(WX5119, WX5142)
--	WX5197 = AND(WX5118, WX5142)
--	WX5199 = AND(WX5117, WX5142)
--	WX5201 = AND(WX5116, WX5142)
--	WX5203 = AND(WX5115, WX5142)
--	WX5205 = AND(WX5114, WX5142)
--	WX5207 = AND(WX5218, WX6175)
--	WX5208 = AND(WX5214, WX5209)
--	WX5211 = AND(CRC_OUT_5_31, WX6176)
--	WX5212 = AND(WX7477, WX5213)
--	WX5215 = AND(WX5657, WX6176)
--	WX5216 = AND(WX6184, WX5217)
--	WX5221 = AND(WX5232, WX6175)
--	WX5222 = AND(WX5228, WX5223)
--	WX5225 = AND(CRC_OUT_5_30, WX6176)
--	WX5226 = AND(WX7484, WX5227)
--	WX5229 = AND(WX5659, WX6176)
--	WX5230 = AND(WX6191, WX5231)
--	WX5235 = AND(WX5246, WX6175)
--	WX5236 = AND(WX5242, WX5237)
--	WX5239 = AND(CRC_OUT_5_29, WX6176)
--	WX5240 = AND(WX7491, WX5241)
--	WX5243 = AND(WX5661, WX6176)
--	WX5244 = AND(WX6198, WX5245)
--	WX5249 = AND(WX5260, WX6175)
--	WX5250 = AND(WX5256, WX5251)
--	WX5253 = AND(CRC_OUT_5_28, WX6176)
--	WX5254 = AND(WX7498, WX5255)
--	WX5257 = AND(WX5663, WX6176)
--	WX5258 = AND(WX6205, WX5259)
--	WX5263 = AND(WX5274, WX6175)
--	WX5264 = AND(WX5270, WX5265)
--	WX5267 = AND(CRC_OUT_5_27, WX6176)
--	WX5268 = AND(WX7505, WX5269)
--	WX5271 = AND(WX5665, WX6176)
--	WX5272 = AND(WX6212, WX5273)
--	WX5277 = AND(WX5288, WX6175)
--	WX5278 = AND(WX5284, WX5279)
--	WX5281 = AND(CRC_OUT_5_26, WX6176)
--	WX5282 = AND(WX7512, WX5283)
--	WX5285 = AND(WX5667, WX6176)
--	WX5286 = AND(WX6219, WX5287)
--	WX5291 = AND(WX5302, WX6175)
--	WX5292 = AND(WX5298, WX5293)
--	WX5295 = AND(CRC_OUT_5_25, WX6176)
--	WX5296 = AND(WX7519, WX5297)
--	WX5299 = AND(WX5669, WX6176)
--	WX5300 = AND(WX6226, WX5301)
--	WX5305 = AND(WX5316, WX6175)
--	WX5306 = AND(WX5312, WX5307)
--	WX5309 = AND(CRC_OUT_5_24, WX6176)
--	WX5310 = AND(WX7526, WX5311)
--	WX5313 = AND(WX5671, WX6176)
--	WX5314 = AND(WX6233, WX5315)
--	WX5319 = AND(WX5330, WX6175)
--	WX5320 = AND(WX5326, WX5321)
--	WX5323 = AND(CRC_OUT_5_23, WX6176)
--	WX5324 = AND(WX7533, WX5325)
--	WX5327 = AND(WX5673, WX6176)
--	WX5328 = AND(WX6240, WX5329)
--	WX5333 = AND(WX5344, WX6175)
--	WX5334 = AND(WX5340, WX5335)
--	WX5337 = AND(CRC_OUT_5_22, WX6176)
--	WX5338 = AND(WX7540, WX5339)
--	WX5341 = AND(WX5675, WX6176)
--	WX5342 = AND(WX6247, WX5343)
--	WX5347 = AND(WX5358, WX6175)
--	WX5348 = AND(WX5354, WX5349)
--	WX5351 = AND(CRC_OUT_5_21, WX6176)
--	WX5352 = AND(WX7547, WX5353)
--	WX5355 = AND(WX5677, WX6176)
--	WX5356 = AND(WX6254, WX5357)
--	WX5361 = AND(WX5372, WX6175)
--	WX5362 = AND(WX5368, WX5363)
--	WX5365 = AND(CRC_OUT_5_20, WX6176)
--	WX5366 = AND(WX7554, WX5367)
--	WX5369 = AND(WX5679, WX6176)
--	WX5370 = AND(WX6261, WX5371)
--	WX5375 = AND(WX5386, WX6175)
--	WX5376 = AND(WX5382, WX5377)
--	WX5379 = AND(CRC_OUT_5_19, WX6176)
--	WX5380 = AND(WX7561, WX5381)
--	WX5383 = AND(WX5681, WX6176)
--	WX5384 = AND(WX6268, WX5385)
--	WX5389 = AND(WX5400, WX6175)
--	WX5390 = AND(WX5396, WX5391)
--	WX5393 = AND(CRC_OUT_5_18, WX6176)
--	WX5394 = AND(WX7568, WX5395)
--	WX5397 = AND(WX5683, WX6176)
--	WX5398 = AND(WX6275, WX5399)
--	WX5403 = AND(WX5414, WX6175)
--	WX5404 = AND(WX5410, WX5405)
--	WX5407 = AND(CRC_OUT_5_17, WX6176)
--	WX5408 = AND(WX7575, WX5409)
--	WX5411 = AND(WX5685, WX6176)
--	WX5412 = AND(WX6282, WX5413)
--	WX5417 = AND(WX5428, WX6175)
--	WX5418 = AND(WX5424, WX5419)
--	WX5421 = AND(CRC_OUT_5_16, WX6176)
--	WX5422 = AND(WX7582, WX5423)
--	WX5425 = AND(WX5687, WX6176)
--	WX5426 = AND(WX6289, WX5427)
--	WX5431 = AND(WX5442, WX6175)
--	WX5432 = AND(WX5438, WX5433)
--	WX5435 = AND(CRC_OUT_5_15, WX6176)
--	WX5436 = AND(WX7589, WX5437)
--	WX5439 = AND(WX5689, WX6176)
--	WX5440 = AND(WX6296, WX5441)
--	WX5445 = AND(WX5456, WX6175)
--	WX5446 = AND(WX5452, WX5447)
--	WX5449 = AND(CRC_OUT_5_14, WX6176)
--	WX5450 = AND(WX7596, WX5451)
--	WX5453 = AND(WX5691, WX6176)
--	WX5454 = AND(WX6303, WX5455)
--	WX5459 = AND(WX5470, WX6175)
--	WX5460 = AND(WX5466, WX5461)
--	WX5463 = AND(CRC_OUT_5_13, WX6176)
--	WX5464 = AND(WX7603, WX5465)
--	WX5467 = AND(WX5693, WX6176)
--	WX5468 = AND(WX6310, WX5469)
--	WX5473 = AND(WX5484, WX6175)
--	WX5474 = AND(WX5480, WX5475)
--	WX5477 = AND(CRC_OUT_5_12, WX6176)
--	WX5478 = AND(WX7610, WX5479)
--	WX5481 = AND(WX5695, WX6176)
--	WX5482 = AND(WX6317, WX5483)
--	WX5487 = AND(WX5498, WX6175)
--	WX5488 = AND(WX5494, WX5489)
--	WX5491 = AND(CRC_OUT_5_11, WX6176)
--	WX5492 = AND(WX7617, WX5493)
--	WX5495 = AND(WX5697, WX6176)
--	WX5496 = AND(WX6324, WX5497)
--	WX5501 = AND(WX5512, WX6175)
--	WX5502 = AND(WX5508, WX5503)
--	WX5505 = AND(CRC_OUT_5_10, WX6176)
--	WX5506 = AND(WX7624, WX5507)
--	WX5509 = AND(WX5699, WX6176)
--	WX5510 = AND(WX6331, WX5511)
--	WX5515 = AND(WX5526, WX6175)
--	WX5516 = AND(WX5522, WX5517)
--	WX5519 = AND(CRC_OUT_5_9, WX6176)
--	WX5520 = AND(WX7631, WX5521)
--	WX5523 = AND(WX5701, WX6176)
--	WX5524 = AND(WX6338, WX5525)
--	WX5529 = AND(WX5540, WX6175)
--	WX5530 = AND(WX5536, WX5531)
--	WX5533 = AND(CRC_OUT_5_8, WX6176)
--	WX5534 = AND(WX7638, WX5535)
--	WX5537 = AND(WX5703, WX6176)
--	WX5538 = AND(WX6345, WX5539)
--	WX5543 = AND(WX5554, WX6175)
--	WX5544 = AND(WX5550, WX5545)
--	WX5547 = AND(CRC_OUT_5_7, WX6176)
--	WX5548 = AND(WX7645, WX5549)
--	WX5551 = AND(WX5705, WX6176)
--	WX5552 = AND(WX6352, WX5553)
--	WX5557 = AND(WX5568, WX6175)
--	WX5558 = AND(WX5564, WX5559)
--	WX5561 = AND(CRC_OUT_5_6, WX6176)
--	WX5562 = AND(WX7652, WX5563)
--	WX5565 = AND(WX5707, WX6176)
--	WX5566 = AND(WX6359, WX5567)
--	WX5571 = AND(WX5582, WX6175)
--	WX5572 = AND(WX5578, WX5573)
--	WX5575 = AND(CRC_OUT_5_5, WX6176)
--	WX5576 = AND(WX7659, WX5577)
--	WX5579 = AND(WX5709, WX6176)
--	WX5580 = AND(WX6366, WX5581)
--	WX5585 = AND(WX5596, WX6175)
--	WX5586 = AND(WX5592, WX5587)
--	WX5589 = AND(CRC_OUT_5_4, WX6176)
--	WX5590 = AND(WX7666, WX5591)
--	WX5593 = AND(WX5711, WX6176)
--	WX5594 = AND(WX6373, WX5595)
--	WX5599 = AND(WX5610, WX6175)
--	WX5600 = AND(WX5606, WX5601)
--	WX5603 = AND(CRC_OUT_5_3, WX6176)
--	WX5604 = AND(WX7673, WX5605)
--	WX5607 = AND(WX5713, WX6176)
--	WX5608 = AND(WX6380, WX5609)
--	WX5613 = AND(WX5624, WX6175)
--	WX5614 = AND(WX5620, WX5615)
--	WX5617 = AND(CRC_OUT_5_2, WX6176)
--	WX5618 = AND(WX7680, WX5619)
--	WX5621 = AND(WX5715, WX6176)
--	WX5622 = AND(WX6387, WX5623)
--	WX5627 = AND(WX5638, WX6175)
--	WX5628 = AND(WX5634, WX5629)
--	WX5631 = AND(CRC_OUT_5_1, WX6176)
--	WX5632 = AND(WX7687, WX5633)
--	WX5635 = AND(WX5717, WX6176)
--	WX5636 = AND(WX6394, WX5637)
--	WX5641 = AND(WX5652, WX6175)
--	WX5642 = AND(WX5648, WX5643)
--	WX5645 = AND(CRC_OUT_5_0, WX6176)
--	WX5646 = AND(WX7694, WX5647)
--	WX5649 = AND(WX5719, WX6176)
--	WX5650 = AND(WX6401, WX5651)
--	WX5656 = AND(WX5659, RESET)
--	WX5658 = AND(WX5661, RESET)
--	WX5660 = AND(WX5663, RESET)
--	WX5662 = AND(WX5665, RESET)
--	WX5664 = AND(WX5667, RESET)
--	WX5666 = AND(WX5669, RESET)
--	WX5668 = AND(WX5671, RESET)
--	WX5670 = AND(WX5673, RESET)
--	WX5672 = AND(WX5675, RESET)
--	WX5674 = AND(WX5677, RESET)
--	WX5676 = AND(WX5679, RESET)
--	WX5678 = AND(WX5681, RESET)
--	WX5680 = AND(WX5683, RESET)
--	WX5682 = AND(WX5685, RESET)
--	WX5684 = AND(WX5687, RESET)
--	WX5686 = AND(WX5689, RESET)
--	WX5688 = AND(WX5691, RESET)
--	WX5690 = AND(WX5693, RESET)
--	WX5692 = AND(WX5695, RESET)
--	WX5694 = AND(WX5697, RESET)
--	WX5696 = AND(WX5699, RESET)
--	WX5698 = AND(WX5701, RESET)
--	WX5700 = AND(WX5703, RESET)
--	WX5702 = AND(WX5705, RESET)
--	WX5704 = AND(WX5707, RESET)
--	WX5706 = AND(WX5709, RESET)
--	WX5708 = AND(WX5711, RESET)
--	WX5710 = AND(WX5713, RESET)
--	WX5712 = AND(WX5715, RESET)
--	WX5714 = AND(WX5717, RESET)
--	WX5716 = AND(WX5719, RESET)
--	WX5718 = AND(WX5655, RESET)
--	WX5816 = AND(WX5220, RESET)
--	WX5818 = AND(WX5234, RESET)
--	WX5820 = AND(WX5248, RESET)
--	WX5822 = AND(WX5262, RESET)
--	WX5824 = AND(WX5276, RESET)
--	WX5826 = AND(WX5290, RESET)
--	WX5828 = AND(WX5304, RESET)
--	WX5830 = AND(WX5318, RESET)
--	WX5832 = AND(WX5332, RESET)
--	WX5834 = AND(WX5346, RESET)
--	WX5836 = AND(WX5360, RESET)
--	WX5838 = AND(WX5374, RESET)
--	WX5840 = AND(WX5388, RESET)
--	WX5842 = AND(WX5402, RESET)
--	WX5844 = AND(WX5416, RESET)
--	WX5846 = AND(WX5430, RESET)
--	WX5848 = AND(WX5444, RESET)
--	WX5850 = AND(WX5458, RESET)
--	WX5852 = AND(WX5472, RESET)
--	WX5854 = AND(WX5486, RESET)
--	WX5856 = AND(WX5500, RESET)
--	WX5858 = AND(WX5514, RESET)
--	WX5860 = AND(WX5528, RESET)
--	WX5862 = AND(WX5542, RESET)
--	WX5864 = AND(WX5556, RESET)
--	WX5866 = AND(WX5570, RESET)
--	WX5868 = AND(WX5584, RESET)
--	WX5870 = AND(WX5598, RESET)
--	WX5872 = AND(WX5612, RESET)
--	WX5874 = AND(WX5626, RESET)
--	WX5876 = AND(WX5640, RESET)
--	WX5878 = AND(WX5654, RESET)
--	WX5880 = AND(WX5817, RESET)
--	WX5882 = AND(WX5819, RESET)
--	WX5884 = AND(WX5821, RESET)
--	WX5886 = AND(WX5823, RESET)
--	WX5888 = AND(WX5825, RESET)
--	WX5890 = AND(WX5827, RESET)
--	WX5892 = AND(WX5829, RESET)
--	WX5894 = AND(WX5831, RESET)
--	WX5896 = AND(WX5833, RESET)
--	WX5898 = AND(WX5835, RESET)
--	WX5900 = AND(WX5837, RESET)
--	WX5902 = AND(WX5839, RESET)
--	WX5904 = AND(WX5841, RESET)
--	WX5906 = AND(WX5843, RESET)
--	WX5908 = AND(WX5845, RESET)
--	WX5910 = AND(WX5847, RESET)
--	WX5912 = AND(WX5849, RESET)
--	WX5914 = AND(WX5851, RESET)
--	WX5916 = AND(WX5853, RESET)
--	WX5918 = AND(WX5855, RESET)
--	WX5920 = AND(WX5857, RESET)
--	WX5922 = AND(WX5859, RESET)
--	WX5924 = AND(WX5861, RESET)
--	WX5926 = AND(WX5863, RESET)
--	WX5928 = AND(WX5865, RESET)
--	WX5930 = AND(WX5867, RESET)
--	WX5932 = AND(WX5869, RESET)
--	WX5934 = AND(WX5871, RESET)
--	WX5936 = AND(WX5873, RESET)
--	WX5938 = AND(WX5875, RESET)
--	WX5940 = AND(WX5877, RESET)
--	WX5942 = AND(WX5879, RESET)
--	WX5944 = AND(WX5881, RESET)
--	WX5946 = AND(WX5883, RESET)
--	WX5948 = AND(WX5885, RESET)
--	WX5950 = AND(WX5887, RESET)
--	WX5952 = AND(WX5889, RESET)
--	WX5954 = AND(WX5891, RESET)
--	WX5956 = AND(WX5893, RESET)
--	WX5958 = AND(WX5895, RESET)
--	WX5960 = AND(WX5897, RESET)
--	WX5962 = AND(WX5899, RESET)
--	WX5964 = AND(WX5901, RESET)
--	WX5966 = AND(WX5903, RESET)
--	WX5968 = AND(WX5905, RESET)
--	WX5970 = AND(WX5907, RESET)
--	WX5972 = AND(WX5909, RESET)
--	WX5974 = AND(WX5911, RESET)
--	WX5976 = AND(WX5913, RESET)
--	WX5978 = AND(WX5915, RESET)
--	WX5980 = AND(WX5917, RESET)
--	WX5982 = AND(WX5919, RESET)
--	WX5984 = AND(WX5921, RESET)
--	WX5986 = AND(WX5923, RESET)
--	WX5988 = AND(WX5925, RESET)
--	WX5990 = AND(WX5927, RESET)
--	WX5992 = AND(WX5929, RESET)
--	WX5994 = AND(WX5931, RESET)
--	WX5996 = AND(WX5933, RESET)
--	WX5998 = AND(WX5935, RESET)
--	WX6000 = AND(WX5937, RESET)
--	WX6002 = AND(WX5939, RESET)
--	WX6004 = AND(WX5941, RESET)
--	WX6006 = AND(WX5943, RESET)
--	WX6008 = AND(WX5945, RESET)
--	WX6010 = AND(WX5947, RESET)
--	WX6012 = AND(WX5949, RESET)
--	WX6014 = AND(WX5951, RESET)
--	WX6016 = AND(WX5953, RESET)
--	WX6018 = AND(WX5955, RESET)
--	WX6020 = AND(WX5957, RESET)
--	WX6022 = AND(WX5959, RESET)
--	WX6024 = AND(WX5961, RESET)
--	WX6026 = AND(WX5963, RESET)
--	WX6028 = AND(WX5965, RESET)
--	WX6030 = AND(WX5967, RESET)
--	WX6032 = AND(WX5969, RESET)
--	WX6034 = AND(WX5971, RESET)
--	WX6036 = AND(WX5973, RESET)
--	WX6038 = AND(WX5975, RESET)
--	WX6040 = AND(WX5977, RESET)
--	WX6042 = AND(WX5979, RESET)
--	WX6044 = AND(WX5981, RESET)
--	WX6046 = AND(WX5983, RESET)
--	WX6048 = AND(WX5985, RESET)
--	WX6050 = AND(WX5987, RESET)
--	WX6052 = AND(WX5989, RESET)
--	WX6054 = AND(WX5991, RESET)
--	WX6056 = AND(WX5993, RESET)
--	WX6058 = AND(WX5995, RESET)
--	WX6060 = AND(WX5997, RESET)
--	WX6062 = AND(WX5999, RESET)
--	WX6064 = AND(WX6001, RESET)
--	WX6066 = AND(WX6003, RESET)
--	WX6068 = AND(WX6005, RESET)
--	WX6070 = AND(WX6007, RESET)
--	WX6179 = AND(WX6178, WX6177)
--	WX6180 = AND(WX5752, WX6181)
--	WX6186 = AND(WX6185, WX6177)
--	WX6187 = AND(WX5753, WX6188)
--	WX6193 = AND(WX6192, WX6177)
--	WX6194 = AND(WX5754, WX6195)
--	WX6200 = AND(WX6199, WX6177)
--	WX6201 = AND(WX5755, WX6202)
--	WX6207 = AND(WX6206, WX6177)
--	WX6208 = AND(WX5756, WX6209)
--	WX6214 = AND(WX6213, WX6177)
--	WX6215 = AND(WX5757, WX6216)
--	WX6221 = AND(WX6220, WX6177)
--	WX6222 = AND(WX5758, WX6223)
--	WX6228 = AND(WX6227, WX6177)
--	WX6229 = AND(WX5759, WX6230)
--	WX6235 = AND(WX6234, WX6177)
--	WX6236 = AND(WX5760, WX6237)
--	WX6242 = AND(WX6241, WX6177)
--	WX6243 = AND(WX5761, WX6244)
--	WX6249 = AND(WX6248, WX6177)
--	WX6250 = AND(WX5762, WX6251)
--	WX6256 = AND(WX6255, WX6177)
--	WX6257 = AND(WX5763, WX6258)
--	WX6263 = AND(WX6262, WX6177)
--	WX6264 = AND(WX5764, WX6265)
--	WX6270 = AND(WX6269, WX6177)
--	WX6271 = AND(WX5765, WX6272)
--	WX6277 = AND(WX6276, WX6177)
--	WX6278 = AND(WX5766, WX6279)
--	WX6284 = AND(WX6283, WX6177)
--	WX6285 = AND(WX5767, WX6286)
--	WX6291 = AND(WX6290, WX6177)
--	WX6292 = AND(WX5768, WX6293)
--	WX6298 = AND(WX6297, WX6177)
--	WX6299 = AND(WX5769, WX6300)
--	WX6305 = AND(WX6304, WX6177)
--	WX6306 = AND(WX5770, WX6307)
--	WX6312 = AND(WX6311, WX6177)
--	WX6313 = AND(WX5771, WX6314)
--	WX6319 = AND(WX6318, WX6177)
--	WX6320 = AND(WX5772, WX6321)
--	WX6326 = AND(WX6325, WX6177)
--	WX6327 = AND(WX5773, WX6328)
--	WX6333 = AND(WX6332, WX6177)
--	WX6334 = AND(WX5774, WX6335)
--	WX6340 = AND(WX6339, WX6177)
--	WX6341 = AND(WX5775, WX6342)
--	WX6347 = AND(WX6346, WX6177)
--	WX6348 = AND(WX5776, WX6349)
--	WX6354 = AND(WX6353, WX6177)
--	WX6355 = AND(WX5777, WX6356)
--	WX6361 = AND(WX6360, WX6177)
--	WX6362 = AND(WX5778, WX6363)
--	WX6368 = AND(WX6367, WX6177)
--	WX6369 = AND(WX5779, WX6370)
--	WX6375 = AND(WX6374, WX6177)
--	WX6376 = AND(WX5780, WX6377)
--	WX6382 = AND(WX6381, WX6177)
--	WX6383 = AND(WX5781, WX6384)
--	WX6389 = AND(WX6388, WX6177)
--	WX6390 = AND(WX5782, WX6391)
--	WX6396 = AND(WX6395, WX6177)
--	WX6397 = AND(WX5783, WX6398)
--	WX6436 = AND(WX6406, WX6435)
--	WX6438 = AND(WX6434, WX6435)
--	WX6440 = AND(WX6433, WX6435)
--	WX6442 = AND(WX6432, WX6435)
--	WX6444 = AND(WX6405, WX6435)
--	WX6446 = AND(WX6431, WX6435)
--	WX6448 = AND(WX6430, WX6435)
--	WX6450 = AND(WX6429, WX6435)
--	WX6452 = AND(WX6428, WX6435)
--	WX6454 = AND(WX6427, WX6435)
--	WX6456 = AND(WX6426, WX6435)
--	WX6458 = AND(WX6404, WX6435)
--	WX6460 = AND(WX6425, WX6435)
--	WX6462 = AND(WX6424, WX6435)
--	WX6464 = AND(WX6423, WX6435)
--	WX6466 = AND(WX6422, WX6435)
--	WX6468 = AND(WX6403, WX6435)
--	WX6470 = AND(WX6421, WX6435)
--	WX6472 = AND(WX6420, WX6435)
--	WX6474 = AND(WX6419, WX6435)
--	WX6476 = AND(WX6418, WX6435)
--	WX6478 = AND(WX6417, WX6435)
--	WX6480 = AND(WX6416, WX6435)
--	WX6482 = AND(WX6415, WX6435)
--	WX6484 = AND(WX6414, WX6435)
--	WX6486 = AND(WX6413, WX6435)
--	WX6488 = AND(WX6412, WX6435)
--	WX6490 = AND(WX6411, WX6435)
--	WX6492 = AND(WX6410, WX6435)
--	WX6494 = AND(WX6409, WX6435)
--	WX6496 = AND(WX6408, WX6435)
--	WX6498 = AND(WX6407, WX6435)
--	WX6500 = AND(WX6511, WX7468)
--	WX6501 = AND(WX6507, WX6502)
--	WX6504 = AND(CRC_OUT_4_31, WX7469)
--	WX6505 = AND(WX8770, WX6506)
--	WX6508 = AND(WX6950, WX7469)
--	WX6509 = AND(WX7477, WX6510)
--	WX6514 = AND(WX6525, WX7468)
--	WX6515 = AND(WX6521, WX6516)
--	WX6518 = AND(CRC_OUT_4_30, WX7469)
--	WX6519 = AND(WX8777, WX6520)
--	WX6522 = AND(WX6952, WX7469)
--	WX6523 = AND(WX7484, WX6524)
--	WX6528 = AND(WX6539, WX7468)
--	WX6529 = AND(WX6535, WX6530)
--	WX6532 = AND(CRC_OUT_4_29, WX7469)
--	WX6533 = AND(WX8784, WX6534)
--	WX6536 = AND(WX6954, WX7469)
--	WX6537 = AND(WX7491, WX6538)
--	WX6542 = AND(WX6553, WX7468)
--	WX6543 = AND(WX6549, WX6544)
--	WX6546 = AND(CRC_OUT_4_28, WX7469)
--	WX6547 = AND(WX8791, WX6548)
--	WX6550 = AND(WX6956, WX7469)
--	WX6551 = AND(WX7498, WX6552)
--	WX6556 = AND(WX6567, WX7468)
--	WX6557 = AND(WX6563, WX6558)
--	WX6560 = AND(CRC_OUT_4_27, WX7469)
--	WX6561 = AND(WX8798, WX6562)
--	WX6564 = AND(WX6958, WX7469)
--	WX6565 = AND(WX7505, WX6566)
--	WX6570 = AND(WX6581, WX7468)
--	WX6571 = AND(WX6577, WX6572)
--	WX6574 = AND(CRC_OUT_4_26, WX7469)
--	WX6575 = AND(WX8805, WX6576)
--	WX6578 = AND(WX6960, WX7469)
--	WX6579 = AND(WX7512, WX6580)
--	WX6584 = AND(WX6595, WX7468)
--	WX6585 = AND(WX6591, WX6586)
--	WX6588 = AND(CRC_OUT_4_25, WX7469)
--	WX6589 = AND(WX8812, WX6590)
--	WX6592 = AND(WX6962, WX7469)
--	WX6593 = AND(WX7519, WX6594)
--	WX6598 = AND(WX6609, WX7468)
--	WX6599 = AND(WX6605, WX6600)
--	WX6602 = AND(CRC_OUT_4_24, WX7469)
--	WX6603 = AND(WX8819, WX6604)
--	WX6606 = AND(WX6964, WX7469)
--	WX6607 = AND(WX7526, WX6608)
--	WX6612 = AND(WX6623, WX7468)
--	WX6613 = AND(WX6619, WX6614)
--	WX6616 = AND(CRC_OUT_4_23, WX7469)
--	WX6617 = AND(WX8826, WX6618)
--	WX6620 = AND(WX6966, WX7469)
--	WX6621 = AND(WX7533, WX6622)
--	WX6626 = AND(WX6637, WX7468)
--	WX6627 = AND(WX6633, WX6628)
--	WX6630 = AND(CRC_OUT_4_22, WX7469)
--	WX6631 = AND(WX8833, WX6632)
--	WX6634 = AND(WX6968, WX7469)
--	WX6635 = AND(WX7540, WX6636)
--	WX6640 = AND(WX6651, WX7468)
--	WX6641 = AND(WX6647, WX6642)
--	WX6644 = AND(CRC_OUT_4_21, WX7469)
--	WX6645 = AND(WX8840, WX6646)
--	WX6648 = AND(WX6970, WX7469)
--	WX6649 = AND(WX7547, WX6650)
--	WX6654 = AND(WX6665, WX7468)
--	WX6655 = AND(WX6661, WX6656)
--	WX6658 = AND(CRC_OUT_4_20, WX7469)
--	WX6659 = AND(WX8847, WX6660)
--	WX6662 = AND(WX6972, WX7469)
--	WX6663 = AND(WX7554, WX6664)
--	WX6668 = AND(WX6679, WX7468)
--	WX6669 = AND(WX6675, WX6670)
--	WX6672 = AND(CRC_OUT_4_19, WX7469)
--	WX6673 = AND(WX8854, WX6674)
--	WX6676 = AND(WX6974, WX7469)
--	WX6677 = AND(WX7561, WX6678)
--	WX6682 = AND(WX6693, WX7468)
--	WX6683 = AND(WX6689, WX6684)
--	WX6686 = AND(CRC_OUT_4_18, WX7469)
--	WX6687 = AND(WX8861, WX6688)
--	WX6690 = AND(WX6976, WX7469)
--	WX6691 = AND(WX7568, WX6692)
--	WX6696 = AND(WX6707, WX7468)
--	WX6697 = AND(WX6703, WX6698)
--	WX6700 = AND(CRC_OUT_4_17, WX7469)
--	WX6701 = AND(WX8868, WX6702)
--	WX6704 = AND(WX6978, WX7469)
--	WX6705 = AND(WX7575, WX6706)
--	WX6710 = AND(WX6721, WX7468)
--	WX6711 = AND(WX6717, WX6712)
--	WX6714 = AND(CRC_OUT_4_16, WX7469)
--	WX6715 = AND(WX8875, WX6716)
--	WX6718 = AND(WX6980, WX7469)
--	WX6719 = AND(WX7582, WX6720)
--	WX6724 = AND(WX6735, WX7468)
--	WX6725 = AND(WX6731, WX6726)
--	WX6728 = AND(CRC_OUT_4_15, WX7469)
--	WX6729 = AND(WX8882, WX6730)
--	WX6732 = AND(WX6982, WX7469)
--	WX6733 = AND(WX7589, WX6734)
--	WX6738 = AND(WX6749, WX7468)
--	WX6739 = AND(WX6745, WX6740)
--	WX6742 = AND(CRC_OUT_4_14, WX7469)
--	WX6743 = AND(WX8889, WX6744)
--	WX6746 = AND(WX6984, WX7469)
--	WX6747 = AND(WX7596, WX6748)
--	WX6752 = AND(WX6763, WX7468)
--	WX6753 = AND(WX6759, WX6754)
--	WX6756 = AND(CRC_OUT_4_13, WX7469)
--	WX6757 = AND(WX8896, WX6758)
--	WX6760 = AND(WX6986, WX7469)
--	WX6761 = AND(WX7603, WX6762)
--	WX6766 = AND(WX6777, WX7468)
--	WX6767 = AND(WX6773, WX6768)
--	WX6770 = AND(CRC_OUT_4_12, WX7469)
--	WX6771 = AND(WX8903, WX6772)
--	WX6774 = AND(WX6988, WX7469)
--	WX6775 = AND(WX7610, WX6776)
--	WX6780 = AND(WX6791, WX7468)
--	WX6781 = AND(WX6787, WX6782)
--	WX6784 = AND(CRC_OUT_4_11, WX7469)
--	WX6785 = AND(WX8910, WX6786)
--	WX6788 = AND(WX6990, WX7469)
--	WX6789 = AND(WX7617, WX6790)
--	WX6794 = AND(WX6805, WX7468)
--	WX6795 = AND(WX6801, WX6796)
--	WX6798 = AND(CRC_OUT_4_10, WX7469)
--	WX6799 = AND(WX8917, WX6800)
--	WX6802 = AND(WX6992, WX7469)
--	WX6803 = AND(WX7624, WX6804)
--	WX6808 = AND(WX6819, WX7468)
--	WX6809 = AND(WX6815, WX6810)
--	WX6812 = AND(CRC_OUT_4_9, WX7469)
--	WX6813 = AND(WX8924, WX6814)
--	WX6816 = AND(WX6994, WX7469)
--	WX6817 = AND(WX7631, WX6818)
--	WX6822 = AND(WX6833, WX7468)
--	WX6823 = AND(WX6829, WX6824)
--	WX6826 = AND(CRC_OUT_4_8, WX7469)
--	WX6827 = AND(WX8931, WX6828)
--	WX6830 = AND(WX6996, WX7469)
--	WX6831 = AND(WX7638, WX6832)
--	WX6836 = AND(WX6847, WX7468)
--	WX6837 = AND(WX6843, WX6838)
--	WX6840 = AND(CRC_OUT_4_7, WX7469)
--	WX6841 = AND(WX8938, WX6842)
--	WX6844 = AND(WX6998, WX7469)
--	WX6845 = AND(WX7645, WX6846)
--	WX6850 = AND(WX6861, WX7468)
--	WX6851 = AND(WX6857, WX6852)
--	WX6854 = AND(CRC_OUT_4_6, WX7469)
--	WX6855 = AND(WX8945, WX6856)
--	WX6858 = AND(WX7000, WX7469)
--	WX6859 = AND(WX7652, WX6860)
--	WX6864 = AND(WX6875, WX7468)
--	WX6865 = AND(WX6871, WX6866)
--	WX6868 = AND(CRC_OUT_4_5, WX7469)
--	WX6869 = AND(WX8952, WX6870)
--	WX6872 = AND(WX7002, WX7469)
--	WX6873 = AND(WX7659, WX6874)
--	WX6878 = AND(WX6889, WX7468)
--	WX6879 = AND(WX6885, WX6880)
--	WX6882 = AND(CRC_OUT_4_4, WX7469)
--	WX6883 = AND(WX8959, WX6884)
--	WX6886 = AND(WX7004, WX7469)
--	WX6887 = AND(WX7666, WX6888)
--	WX6892 = AND(WX6903, WX7468)
--	WX6893 = AND(WX6899, WX6894)
--	WX6896 = AND(CRC_OUT_4_3, WX7469)
--	WX6897 = AND(WX8966, WX6898)
--	WX6900 = AND(WX7006, WX7469)
--	WX6901 = AND(WX7673, WX6902)
--	WX6906 = AND(WX6917, WX7468)
--	WX6907 = AND(WX6913, WX6908)
--	WX6910 = AND(CRC_OUT_4_2, WX7469)
--	WX6911 = AND(WX8973, WX6912)
--	WX6914 = AND(WX7008, WX7469)
--	WX6915 = AND(WX7680, WX6916)
--	WX6920 = AND(WX6931, WX7468)
--	WX6921 = AND(WX6927, WX6922)
--	WX6924 = AND(CRC_OUT_4_1, WX7469)
--	WX6925 = AND(WX8980, WX6926)
--	WX6928 = AND(WX7010, WX7469)
--	WX6929 = AND(WX7687, WX6930)
--	WX6934 = AND(WX6945, WX7468)
--	WX6935 = AND(WX6941, WX6936)
--	WX6938 = AND(CRC_OUT_4_0, WX7469)
--	WX6939 = AND(WX8987, WX6940)
--	WX6942 = AND(WX7012, WX7469)
--	WX6943 = AND(WX7694, WX6944)
--	WX6949 = AND(WX6952, RESET)
--	WX6951 = AND(WX6954, RESET)
--	WX6953 = AND(WX6956, RESET)
--	WX6955 = AND(WX6958, RESET)
--	WX6957 = AND(WX6960, RESET)
--	WX6959 = AND(WX6962, RESET)
--	WX6961 = AND(WX6964, RESET)
--	WX6963 = AND(WX6966, RESET)
--	WX6965 = AND(WX6968, RESET)
--	WX6967 = AND(WX6970, RESET)
--	WX6969 = AND(WX6972, RESET)
--	WX6971 = AND(WX6974, RESET)
--	WX6973 = AND(WX6976, RESET)
--	WX6975 = AND(WX6978, RESET)
--	WX6977 = AND(WX6980, RESET)
--	WX6979 = AND(WX6982, RESET)
--	WX6981 = AND(WX6984, RESET)
--	WX6983 = AND(WX6986, RESET)
--	WX6985 = AND(WX6988, RESET)
--	WX6987 = AND(WX6990, RESET)
--	WX6989 = AND(WX6992, RESET)
--	WX6991 = AND(WX6994, RESET)
--	WX6993 = AND(WX6996, RESET)
--	WX6995 = AND(WX6998, RESET)
--	WX6997 = AND(WX7000, RESET)
--	WX6999 = AND(WX7002, RESET)
--	WX7001 = AND(WX7004, RESET)
--	WX7003 = AND(WX7006, RESET)
--	WX7005 = AND(WX7008, RESET)
--	WX7007 = AND(WX7010, RESET)
--	WX7009 = AND(WX7012, RESET)
--	WX7011 = AND(WX6948, RESET)
--	WX7109 = AND(WX6513, RESET)
--	WX7111 = AND(WX6527, RESET)
--	WX7113 = AND(WX6541, RESET)
--	WX7115 = AND(WX6555, RESET)
--	WX7117 = AND(WX6569, RESET)
--	WX7119 = AND(WX6583, RESET)
--	WX7121 = AND(WX6597, RESET)
--	WX7123 = AND(WX6611, RESET)
--	WX7125 = AND(WX6625, RESET)
--	WX7127 = AND(WX6639, RESET)
--	WX7129 = AND(WX6653, RESET)
--	WX7131 = AND(WX6667, RESET)
--	WX7133 = AND(WX6681, RESET)
--	WX7135 = AND(WX6695, RESET)
--	WX7137 = AND(WX6709, RESET)
--	WX7139 = AND(WX6723, RESET)
--	WX7141 = AND(WX6737, RESET)
--	WX7143 = AND(WX6751, RESET)
--	WX7145 = AND(WX6765, RESET)
--	WX7147 = AND(WX6779, RESET)
--	WX7149 = AND(WX6793, RESET)
--	WX7151 = AND(WX6807, RESET)
--	WX7153 = AND(WX6821, RESET)
--	WX7155 = AND(WX6835, RESET)
--	WX7157 = AND(WX6849, RESET)
--	WX7159 = AND(WX6863, RESET)
--	WX7161 = AND(WX6877, RESET)
--	WX7163 = AND(WX6891, RESET)
--	WX7165 = AND(WX6905, RESET)
--	WX7167 = AND(WX6919, RESET)
--	WX7169 = AND(WX6933, RESET)
--	WX7171 = AND(WX6947, RESET)
--	WX7173 = AND(WX7110, RESET)
--	WX7175 = AND(WX7112, RESET)
--	WX7177 = AND(WX7114, RESET)
--	WX7179 = AND(WX7116, RESET)
--	WX7181 = AND(WX7118, RESET)
--	WX7183 = AND(WX7120, RESET)
--	WX7185 = AND(WX7122, RESET)
--	WX7187 = AND(WX7124, RESET)
--	WX7189 = AND(WX7126, RESET)
--	WX7191 = AND(WX7128, RESET)
--	WX7193 = AND(WX7130, RESET)
--	WX7195 = AND(WX7132, RESET)
--	WX7197 = AND(WX7134, RESET)
--	WX7199 = AND(WX7136, RESET)
--	WX7201 = AND(WX7138, RESET)
--	WX7203 = AND(WX7140, RESET)
--	WX7205 = AND(WX7142, RESET)
--	WX7207 = AND(WX7144, RESET)
--	WX7209 = AND(WX7146, RESET)
--	WX7211 = AND(WX7148, RESET)
--	WX7213 = AND(WX7150, RESET)
--	WX7215 = AND(WX7152, RESET)
--	WX7217 = AND(WX7154, RESET)
--	WX7219 = AND(WX7156, RESET)
--	WX7221 = AND(WX7158, RESET)
--	WX7223 = AND(WX7160, RESET)
--	WX7225 = AND(WX7162, RESET)
--	WX7227 = AND(WX7164, RESET)
--	WX7229 = AND(WX7166, RESET)
--	WX7231 = AND(WX7168, RESET)
--	WX7233 = AND(WX7170, RESET)
--	WX7235 = AND(WX7172, RESET)
--	WX7237 = AND(WX7174, RESET)
--	WX7239 = AND(WX7176, RESET)
--	WX7241 = AND(WX7178, RESET)
--	WX7243 = AND(WX7180, RESET)
--	WX7245 = AND(WX7182, RESET)
--	WX7247 = AND(WX7184, RESET)
--	WX7249 = AND(WX7186, RESET)
--	WX7251 = AND(WX7188, RESET)
--	WX7253 = AND(WX7190, RESET)
--	WX7255 = AND(WX7192, RESET)
--	WX7257 = AND(WX7194, RESET)
--	WX7259 = AND(WX7196, RESET)
--	WX7261 = AND(WX7198, RESET)
--	WX7263 = AND(WX7200, RESET)
--	WX7265 = AND(WX7202, RESET)
--	WX7267 = AND(WX7204, RESET)
--	WX7269 = AND(WX7206, RESET)
--	WX7271 = AND(WX7208, RESET)
--	WX7273 = AND(WX7210, RESET)
--	WX7275 = AND(WX7212, RESET)
--	WX7277 = AND(WX7214, RESET)
--	WX7279 = AND(WX7216, RESET)
--	WX7281 = AND(WX7218, RESET)
--	WX7283 = AND(WX7220, RESET)
--	WX7285 = AND(WX7222, RESET)
--	WX7287 = AND(WX7224, RESET)
--	WX7289 = AND(WX7226, RESET)
--	WX7291 = AND(WX7228, RESET)
--	WX7293 = AND(WX7230, RESET)
--	WX7295 = AND(WX7232, RESET)
--	WX7297 = AND(WX7234, RESET)
--	WX7299 = AND(WX7236, RESET)
--	WX7301 = AND(WX7238, RESET)
--	WX7303 = AND(WX7240, RESET)
--	WX7305 = AND(WX7242, RESET)
--	WX7307 = AND(WX7244, RESET)
--	WX7309 = AND(WX7246, RESET)
--	WX7311 = AND(WX7248, RESET)
--	WX7313 = AND(WX7250, RESET)
--	WX7315 = AND(WX7252, RESET)
--	WX7317 = AND(WX7254, RESET)
--	WX7319 = AND(WX7256, RESET)
--	WX7321 = AND(WX7258, RESET)
--	WX7323 = AND(WX7260, RESET)
--	WX7325 = AND(WX7262, RESET)
--	WX7327 = AND(WX7264, RESET)
--	WX7329 = AND(WX7266, RESET)
--	WX7331 = AND(WX7268, RESET)
--	WX7333 = AND(WX7270, RESET)
--	WX7335 = AND(WX7272, RESET)
--	WX7337 = AND(WX7274, RESET)
--	WX7339 = AND(WX7276, RESET)
--	WX7341 = AND(WX7278, RESET)
--	WX7343 = AND(WX7280, RESET)
--	WX7345 = AND(WX7282, RESET)
--	WX7347 = AND(WX7284, RESET)
--	WX7349 = AND(WX7286, RESET)
--	WX7351 = AND(WX7288, RESET)
--	WX7353 = AND(WX7290, RESET)
--	WX7355 = AND(WX7292, RESET)
--	WX7357 = AND(WX7294, RESET)
--	WX7359 = AND(WX7296, RESET)
--	WX7361 = AND(WX7298, RESET)
--	WX7363 = AND(WX7300, RESET)
--	WX7472 = AND(WX7471, WX7470)
--	WX7473 = AND(WX7045, WX7474)
--	WX7479 = AND(WX7478, WX7470)
--	WX7480 = AND(WX7046, WX7481)
--	WX7486 = AND(WX7485, WX7470)
--	WX7487 = AND(WX7047, WX7488)
--	WX7493 = AND(WX7492, WX7470)
--	WX7494 = AND(WX7048, WX7495)
--	WX7500 = AND(WX7499, WX7470)
--	WX7501 = AND(WX7049, WX7502)
--	WX7507 = AND(WX7506, WX7470)
--	WX7508 = AND(WX7050, WX7509)
--	WX7514 = AND(WX7513, WX7470)
--	WX7515 = AND(WX7051, WX7516)
--	WX7521 = AND(WX7520, WX7470)
--	WX7522 = AND(WX7052, WX7523)
--	WX7528 = AND(WX7527, WX7470)
--	WX7529 = AND(WX7053, WX7530)
--	WX7535 = AND(WX7534, WX7470)
--	WX7536 = AND(WX7054, WX7537)
--	WX7542 = AND(WX7541, WX7470)
--	WX7543 = AND(WX7055, WX7544)
--	WX7549 = AND(WX7548, WX7470)
--	WX7550 = AND(WX7056, WX7551)
--	WX7556 = AND(WX7555, WX7470)
--	WX7557 = AND(WX7057, WX7558)
--	WX7563 = AND(WX7562, WX7470)
--	WX7564 = AND(WX7058, WX7565)
--	WX7570 = AND(WX7569, WX7470)
--	WX7571 = AND(WX7059, WX7572)
--	WX7577 = AND(WX7576, WX7470)
--	WX7578 = AND(WX7060, WX7579)
--	WX7584 = AND(WX7583, WX7470)
--	WX7585 = AND(WX7061, WX7586)
--	WX7591 = AND(WX7590, WX7470)
--	WX7592 = AND(WX7062, WX7593)
--	WX7598 = AND(WX7597, WX7470)
--	WX7599 = AND(WX7063, WX7600)
--	WX7605 = AND(WX7604, WX7470)
--	WX7606 = AND(WX7064, WX7607)
--	WX7612 = AND(WX7611, WX7470)
--	WX7613 = AND(WX7065, WX7614)
--	WX7619 = AND(WX7618, WX7470)
--	WX7620 = AND(WX7066, WX7621)
--	WX7626 = AND(WX7625, WX7470)
--	WX7627 = AND(WX7067, WX7628)
--	WX7633 = AND(WX7632, WX7470)
--	WX7634 = AND(WX7068, WX7635)
--	WX7640 = AND(WX7639, WX7470)
--	WX7641 = AND(WX7069, WX7642)
--	WX7647 = AND(WX7646, WX7470)
--	WX7648 = AND(WX7070, WX7649)
--	WX7654 = AND(WX7653, WX7470)
--	WX7655 = AND(WX7071, WX7656)
--	WX7661 = AND(WX7660, WX7470)
--	WX7662 = AND(WX7072, WX7663)
--	WX7668 = AND(WX7667, WX7470)
--	WX7669 = AND(WX7073, WX7670)
--	WX7675 = AND(WX7674, WX7470)
--	WX7676 = AND(WX7074, WX7677)
--	WX7682 = AND(WX7681, WX7470)
--	WX7683 = AND(WX7075, WX7684)
--	WX7689 = AND(WX7688, WX7470)
--	WX7690 = AND(WX7076, WX7691)
--	WX7729 = AND(WX7699, WX7728)
--	WX7731 = AND(WX7727, WX7728)
--	WX7733 = AND(WX7726, WX7728)
--	WX7735 = AND(WX7725, WX7728)
--	WX7737 = AND(WX7698, WX7728)
--	WX7739 = AND(WX7724, WX7728)
--	WX7741 = AND(WX7723, WX7728)
--	WX7743 = AND(WX7722, WX7728)
--	WX7745 = AND(WX7721, WX7728)
--	WX7747 = AND(WX7720, WX7728)
--	WX7749 = AND(WX7719, WX7728)
--	WX7751 = AND(WX7697, WX7728)
--	WX7753 = AND(WX7718, WX7728)
--	WX7755 = AND(WX7717, WX7728)
--	WX7757 = AND(WX7716, WX7728)
--	WX7759 = AND(WX7715, WX7728)
--	WX7761 = AND(WX7696, WX7728)
--	WX7763 = AND(WX7714, WX7728)
--	WX7765 = AND(WX7713, WX7728)
--	WX7767 = AND(WX7712, WX7728)
--	WX7769 = AND(WX7711, WX7728)
--	WX7771 = AND(WX7710, WX7728)
--	WX7773 = AND(WX7709, WX7728)
--	WX7775 = AND(WX7708, WX7728)
--	WX7777 = AND(WX7707, WX7728)
--	WX7779 = AND(WX7706, WX7728)
--	WX7781 = AND(WX7705, WX7728)
--	WX7783 = AND(WX7704, WX7728)
--	WX7785 = AND(WX7703, WX7728)
--	WX7787 = AND(WX7702, WX7728)
--	WX7789 = AND(WX7701, WX7728)
--	WX7791 = AND(WX7700, WX7728)
--	WX7793 = AND(WX7804, WX8761)
--	WX7794 = AND(WX7800, WX7795)
--	WX7797 = AND(CRC_OUT_3_31, WX8762)
--	WX7798 = AND(WX10063, WX7799)
--	WX7801 = AND(WX8243, WX8762)
--	WX7802 = AND(WX8770, WX7803)
--	WX7807 = AND(WX7818, WX8761)
--	WX7808 = AND(WX7814, WX7809)
--	WX7811 = AND(CRC_OUT_3_30, WX8762)
--	WX7812 = AND(WX10070, WX7813)
--	WX7815 = AND(WX8245, WX8762)
--	WX7816 = AND(WX8777, WX7817)
--	WX7821 = AND(WX7832, WX8761)
--	WX7822 = AND(WX7828, WX7823)
--	WX7825 = AND(CRC_OUT_3_29, WX8762)
--	WX7826 = AND(WX10077, WX7827)
--	WX7829 = AND(WX8247, WX8762)
--	WX7830 = AND(WX8784, WX7831)
--	WX7835 = AND(WX7846, WX8761)
--	WX7836 = AND(WX7842, WX7837)
--	WX7839 = AND(CRC_OUT_3_28, WX8762)
--	WX7840 = AND(WX10084, WX7841)
--	WX7843 = AND(WX8249, WX8762)
--	WX7844 = AND(WX8791, WX7845)
--	WX7849 = AND(WX7860, WX8761)
--	WX7850 = AND(WX7856, WX7851)
--	WX7853 = AND(CRC_OUT_3_27, WX8762)
--	WX7854 = AND(WX10091, WX7855)
--	WX7857 = AND(WX8251, WX8762)
--	WX7858 = AND(WX8798, WX7859)
--	WX7863 = AND(WX7874, WX8761)
--	WX7864 = AND(WX7870, WX7865)
--	WX7867 = AND(CRC_OUT_3_26, WX8762)
--	WX7868 = AND(WX10098, WX7869)
--	WX7871 = AND(WX8253, WX8762)
--	WX7872 = AND(WX8805, WX7873)
--	WX7877 = AND(WX7888, WX8761)
--	WX7878 = AND(WX7884, WX7879)
--	WX7881 = AND(CRC_OUT_3_25, WX8762)
--	WX7882 = AND(WX10105, WX7883)
--	WX7885 = AND(WX8255, WX8762)
--	WX7886 = AND(WX8812, WX7887)
--	WX7891 = AND(WX7902, WX8761)
--	WX7892 = AND(WX7898, WX7893)
--	WX7895 = AND(CRC_OUT_3_24, WX8762)
--	WX7896 = AND(WX10112, WX7897)
--	WX7899 = AND(WX8257, WX8762)
--	WX7900 = AND(WX8819, WX7901)
--	WX7905 = AND(WX7916, WX8761)
--	WX7906 = AND(WX7912, WX7907)
--	WX7909 = AND(CRC_OUT_3_23, WX8762)
--	WX7910 = AND(WX10119, WX7911)
--	WX7913 = AND(WX8259, WX8762)
--	WX7914 = AND(WX8826, WX7915)
--	WX7919 = AND(WX7930, WX8761)
--	WX7920 = AND(WX7926, WX7921)
--	WX7923 = AND(CRC_OUT_3_22, WX8762)
--	WX7924 = AND(WX10126, WX7925)
--	WX7927 = AND(WX8261, WX8762)
--	WX7928 = AND(WX8833, WX7929)
--	WX7933 = AND(WX7944, WX8761)
--	WX7934 = AND(WX7940, WX7935)
--	WX7937 = AND(CRC_OUT_3_21, WX8762)
--	WX7938 = AND(WX10133, WX7939)
--	WX7941 = AND(WX8263, WX8762)
--	WX7942 = AND(WX8840, WX7943)
--	WX7947 = AND(WX7958, WX8761)
--	WX7948 = AND(WX7954, WX7949)
--	WX7951 = AND(CRC_OUT_3_20, WX8762)
--	WX7952 = AND(WX10140, WX7953)
--	WX7955 = AND(WX8265, WX8762)
--	WX7956 = AND(WX8847, WX7957)
--	WX7961 = AND(WX7972, WX8761)
--	WX7962 = AND(WX7968, WX7963)
--	WX7965 = AND(CRC_OUT_3_19, WX8762)
--	WX7966 = AND(WX10147, WX7967)
--	WX7969 = AND(WX8267, WX8762)
--	WX7970 = AND(WX8854, WX7971)
--	WX7975 = AND(WX7986, WX8761)
--	WX7976 = AND(WX7982, WX7977)
--	WX7979 = AND(CRC_OUT_3_18, WX8762)
--	WX7980 = AND(WX10154, WX7981)
--	WX7983 = AND(WX8269, WX8762)
--	WX7984 = AND(WX8861, WX7985)
--	WX7989 = AND(WX8000, WX8761)
--	WX7990 = AND(WX7996, WX7991)
--	WX7993 = AND(CRC_OUT_3_17, WX8762)
--	WX7994 = AND(WX10161, WX7995)
--	WX7997 = AND(WX8271, WX8762)
--	WX7998 = AND(WX8868, WX7999)
--	WX8003 = AND(WX8014, WX8761)
--	WX8004 = AND(WX8010, WX8005)
--	WX8007 = AND(CRC_OUT_3_16, WX8762)
--	WX8008 = AND(WX10168, WX8009)
--	WX8011 = AND(WX8273, WX8762)
--	WX8012 = AND(WX8875, WX8013)
--	WX8017 = AND(WX8028, WX8761)
--	WX8018 = AND(WX8024, WX8019)
--	WX8021 = AND(CRC_OUT_3_15, WX8762)
--	WX8022 = AND(WX10175, WX8023)
--	WX8025 = AND(WX8275, WX8762)
--	WX8026 = AND(WX8882, WX8027)
--	WX8031 = AND(WX8042, WX8761)
--	WX8032 = AND(WX8038, WX8033)
--	WX8035 = AND(CRC_OUT_3_14, WX8762)
--	WX8036 = AND(WX10182, WX8037)
--	WX8039 = AND(WX8277, WX8762)
--	WX8040 = AND(WX8889, WX8041)
--	WX8045 = AND(WX8056, WX8761)
--	WX8046 = AND(WX8052, WX8047)
--	WX8049 = AND(CRC_OUT_3_13, WX8762)
--	WX8050 = AND(WX10189, WX8051)
--	WX8053 = AND(WX8279, WX8762)
--	WX8054 = AND(WX8896, WX8055)
--	WX8059 = AND(WX8070, WX8761)
--	WX8060 = AND(WX8066, WX8061)
--	WX8063 = AND(CRC_OUT_3_12, WX8762)
--	WX8064 = AND(WX10196, WX8065)
--	WX8067 = AND(WX8281, WX8762)
--	WX8068 = AND(WX8903, WX8069)
--	WX8073 = AND(WX8084, WX8761)
--	WX8074 = AND(WX8080, WX8075)
--	WX8077 = AND(CRC_OUT_3_11, WX8762)
--	WX8078 = AND(WX10203, WX8079)
--	WX8081 = AND(WX8283, WX8762)
--	WX8082 = AND(WX8910, WX8083)
--	WX8087 = AND(WX8098, WX8761)
--	WX8088 = AND(WX8094, WX8089)
--	WX8091 = AND(CRC_OUT_3_10, WX8762)
--	WX8092 = AND(WX10210, WX8093)
--	WX8095 = AND(WX8285, WX8762)
--	WX8096 = AND(WX8917, WX8097)
--	WX8101 = AND(WX8112, WX8761)
--	WX8102 = AND(WX8108, WX8103)
--	WX8105 = AND(CRC_OUT_3_9, WX8762)
--	WX8106 = AND(WX10217, WX8107)
--	WX8109 = AND(WX8287, WX8762)
--	WX8110 = AND(WX8924, WX8111)
--	WX8115 = AND(WX8126, WX8761)
--	WX8116 = AND(WX8122, WX8117)
--	WX8119 = AND(CRC_OUT_3_8, WX8762)
--	WX8120 = AND(WX10224, WX8121)
--	WX8123 = AND(WX8289, WX8762)
--	WX8124 = AND(WX8931, WX8125)
--	WX8129 = AND(WX8140, WX8761)
--	WX8130 = AND(WX8136, WX8131)
--	WX8133 = AND(CRC_OUT_3_7, WX8762)
--	WX8134 = AND(WX10231, WX8135)
--	WX8137 = AND(WX8291, WX8762)
--	WX8138 = AND(WX8938, WX8139)
--	WX8143 = AND(WX8154, WX8761)
--	WX8144 = AND(WX8150, WX8145)
--	WX8147 = AND(CRC_OUT_3_6, WX8762)
--	WX8148 = AND(WX10238, WX8149)
--	WX8151 = AND(WX8293, WX8762)
--	WX8152 = AND(WX8945, WX8153)
--	WX8157 = AND(WX8168, WX8761)
--	WX8158 = AND(WX8164, WX8159)
--	WX8161 = AND(CRC_OUT_3_5, WX8762)
--	WX8162 = AND(WX10245, WX8163)
--	WX8165 = AND(WX8295, WX8762)
--	WX8166 = AND(WX8952, WX8167)
--	WX8171 = AND(WX8182, WX8761)
--	WX8172 = AND(WX8178, WX8173)
--	WX8175 = AND(CRC_OUT_3_4, WX8762)
--	WX8176 = AND(WX10252, WX8177)
--	WX8179 = AND(WX8297, WX8762)
--	WX8180 = AND(WX8959, WX8181)
--	WX8185 = AND(WX8196, WX8761)
--	WX8186 = AND(WX8192, WX8187)
--	WX8189 = AND(CRC_OUT_3_3, WX8762)
--	WX8190 = AND(WX10259, WX8191)
--	WX8193 = AND(WX8299, WX8762)
--	WX8194 = AND(WX8966, WX8195)
--	WX8199 = AND(WX8210, WX8761)
--	WX8200 = AND(WX8206, WX8201)
--	WX8203 = AND(CRC_OUT_3_2, WX8762)
--	WX8204 = AND(WX10266, WX8205)
--	WX8207 = AND(WX8301, WX8762)
--	WX8208 = AND(WX8973, WX8209)
--	WX8213 = AND(WX8224, WX8761)
--	WX8214 = AND(WX8220, WX8215)
--	WX8217 = AND(CRC_OUT_3_1, WX8762)
--	WX8218 = AND(WX10273, WX8219)
--	WX8221 = AND(WX8303, WX8762)
--	WX8222 = AND(WX8980, WX8223)
--	WX8227 = AND(WX8238, WX8761)
--	WX8228 = AND(WX8234, WX8229)
--	WX8231 = AND(CRC_OUT_3_0, WX8762)
--	WX8232 = AND(WX10280, WX8233)
--	WX8235 = AND(WX8305, WX8762)
--	WX8236 = AND(WX8987, WX8237)
--	WX8242 = AND(WX8245, RESET)
--	WX8244 = AND(WX8247, RESET)
--	WX8246 = AND(WX8249, RESET)
--	WX8248 = AND(WX8251, RESET)
--	WX8250 = AND(WX8253, RESET)
--	WX8252 = AND(WX8255, RESET)
--	WX8254 = AND(WX8257, RESET)
--	WX8256 = AND(WX8259, RESET)
--	WX8258 = AND(WX8261, RESET)
--	WX8260 = AND(WX8263, RESET)
--	WX8262 = AND(WX8265, RESET)
--	WX8264 = AND(WX8267, RESET)
--	WX8266 = AND(WX8269, RESET)
--	WX8268 = AND(WX8271, RESET)
--	WX8270 = AND(WX8273, RESET)
--	WX8272 = AND(WX8275, RESET)
--	WX8274 = AND(WX8277, RESET)
--	WX8276 = AND(WX8279, RESET)
--	WX8278 = AND(WX8281, RESET)
--	WX8280 = AND(WX8283, RESET)
--	WX8282 = AND(WX8285, RESET)
--	WX8284 = AND(WX8287, RESET)
--	WX8286 = AND(WX8289, RESET)
--	WX8288 = AND(WX8291, RESET)
--	WX8290 = AND(WX8293, RESET)
--	WX8292 = AND(WX8295, RESET)
--	WX8294 = AND(WX8297, RESET)
--	WX8296 = AND(WX8299, RESET)
--	WX8298 = AND(WX8301, RESET)
--	WX8300 = AND(WX8303, RESET)
--	WX8302 = AND(WX8305, RESET)
--	WX8304 = AND(WX8241, RESET)
--	WX8402 = AND(WX7806, RESET)
--	WX8404 = AND(WX7820, RESET)
--	WX8406 = AND(WX7834, RESET)
--	WX8408 = AND(WX7848, RESET)
--	WX8410 = AND(WX7862, RESET)
--	WX8412 = AND(WX7876, RESET)
--	WX8414 = AND(WX7890, RESET)
--	WX8416 = AND(WX7904, RESET)
--	WX8418 = AND(WX7918, RESET)
--	WX8420 = AND(WX7932, RESET)
--	WX8422 = AND(WX7946, RESET)
--	WX8424 = AND(WX7960, RESET)
--	WX8426 = AND(WX7974, RESET)
--	WX8428 = AND(WX7988, RESET)
--	WX8430 = AND(WX8002, RESET)
--	WX8432 = AND(WX8016, RESET)
--	WX8434 = AND(WX8030, RESET)
--	WX8436 = AND(WX8044, RESET)
--	WX8438 = AND(WX8058, RESET)
--	WX8440 = AND(WX8072, RESET)
--	WX8442 = AND(WX8086, RESET)
--	WX8444 = AND(WX8100, RESET)
--	WX8446 = AND(WX8114, RESET)
--	WX8448 = AND(WX8128, RESET)
--	WX8450 = AND(WX8142, RESET)
--	WX8452 = AND(WX8156, RESET)
--	WX8454 = AND(WX8170, RESET)
--	WX8456 = AND(WX8184, RESET)
--	WX8458 = AND(WX8198, RESET)
--	WX8460 = AND(WX8212, RESET)
--	WX8462 = AND(WX8226, RESET)
--	WX8464 = AND(WX8240, RESET)
--	WX8466 = AND(WX8403, RESET)
--	WX8468 = AND(WX8405, RESET)
--	WX8470 = AND(WX8407, RESET)
--	WX8472 = AND(WX8409, RESET)
--	WX8474 = AND(WX8411, RESET)
--	WX8476 = AND(WX8413, RESET)
--	WX8478 = AND(WX8415, RESET)
--	WX8480 = AND(WX8417, RESET)
--	WX8482 = AND(WX8419, RESET)
--	WX8484 = AND(WX8421, RESET)
--	WX8486 = AND(WX8423, RESET)
--	WX8488 = AND(WX8425, RESET)
--	WX8490 = AND(WX8427, RESET)
--	WX8492 = AND(WX8429, RESET)
--	WX8494 = AND(WX8431, RESET)
--	WX8496 = AND(WX8433, RESET)
--	WX8498 = AND(WX8435, RESET)
--	WX8500 = AND(WX8437, RESET)
--	WX8502 = AND(WX8439, RESET)
--	WX8504 = AND(WX8441, RESET)
--	WX8506 = AND(WX8443, RESET)
--	WX8508 = AND(WX8445, RESET)
--	WX8510 = AND(WX8447, RESET)
--	WX8512 = AND(WX8449, RESET)
--	WX8514 = AND(WX8451, RESET)
--	WX8516 = AND(WX8453, RESET)
--	WX8518 = AND(WX8455, RESET)
--	WX8520 = AND(WX8457, RESET)
--	WX8522 = AND(WX8459, RESET)
--	WX8524 = AND(WX8461, RESET)
--	WX8526 = AND(WX8463, RESET)
--	WX8528 = AND(WX8465, RESET)
--	WX8530 = AND(WX8467, RESET)
--	WX8532 = AND(WX8469, RESET)
--	WX8534 = AND(WX8471, RESET)
--	WX8536 = AND(WX8473, RESET)
--	WX8538 = AND(WX8475, RESET)
--	WX8540 = AND(WX8477, RESET)
--	WX8542 = AND(WX8479, RESET)
--	WX8544 = AND(WX8481, RESET)
--	WX8546 = AND(WX8483, RESET)
--	WX8548 = AND(WX8485, RESET)
--	WX8550 = AND(WX8487, RESET)
--	WX8552 = AND(WX8489, RESET)
--	WX8554 = AND(WX8491, RESET)
--	WX8556 = AND(WX8493, RESET)
--	WX8558 = AND(WX8495, RESET)
--	WX8560 = AND(WX8497, RESET)
--	WX8562 = AND(WX8499, RESET)
--	WX8564 = AND(WX8501, RESET)
--	WX8566 = AND(WX8503, RESET)
--	WX8568 = AND(WX8505, RESET)
--	WX8570 = AND(WX8507, RESET)
--	WX8572 = AND(WX8509, RESET)
--	WX8574 = AND(WX8511, RESET)
--	WX8576 = AND(WX8513, RESET)
--	WX8578 = AND(WX8515, RESET)
--	WX8580 = AND(WX8517, RESET)
--	WX8582 = AND(WX8519, RESET)
--	WX8584 = AND(WX8521, RESET)
--	WX8586 = AND(WX8523, RESET)
--	WX8588 = AND(WX8525, RESET)
--	WX8590 = AND(WX8527, RESET)
--	WX8592 = AND(WX8529, RESET)
--	WX8594 = AND(WX8531, RESET)
--	WX8596 = AND(WX8533, RESET)
--	WX8598 = AND(WX8535, RESET)
--	WX8600 = AND(WX8537, RESET)
--	WX8602 = AND(WX8539, RESET)
--	WX8604 = AND(WX8541, RESET)
--	WX8606 = AND(WX8543, RESET)
--	WX8608 = AND(WX8545, RESET)
--	WX8610 = AND(WX8547, RESET)
--	WX8612 = AND(WX8549, RESET)
--	WX8614 = AND(WX8551, RESET)
--	WX8616 = AND(WX8553, RESET)
--	WX8618 = AND(WX8555, RESET)
--	WX8620 = AND(WX8557, RESET)
--	WX8622 = AND(WX8559, RESET)
--	WX8624 = AND(WX8561, RESET)
--	WX8626 = AND(WX8563, RESET)
--	WX8628 = AND(WX8565, RESET)
--	WX8630 = AND(WX8567, RESET)
--	WX8632 = AND(WX8569, RESET)
--	WX8634 = AND(WX8571, RESET)
--	WX8636 = AND(WX8573, RESET)
--	WX8638 = AND(WX8575, RESET)
--	WX8640 = AND(WX8577, RESET)
--	WX8642 = AND(WX8579, RESET)
--	WX8644 = AND(WX8581, RESET)
--	WX8646 = AND(WX8583, RESET)
--	WX8648 = AND(WX8585, RESET)
--	WX8650 = AND(WX8587, RESET)
--	WX8652 = AND(WX8589, RESET)
--	WX8654 = AND(WX8591, RESET)
--	WX8656 = AND(WX8593, RESET)
--	WX8765 = AND(WX8764, WX8763)
--	WX8766 = AND(WX8338, WX8767)
--	WX8772 = AND(WX8771, WX8763)
--	WX8773 = AND(WX8339, WX8774)
--	WX8779 = AND(WX8778, WX8763)
--	WX8780 = AND(WX8340, WX8781)
--	WX8786 = AND(WX8785, WX8763)
--	WX8787 = AND(WX8341, WX8788)
--	WX8793 = AND(WX8792, WX8763)
--	WX8794 = AND(WX8342, WX8795)
--	WX8800 = AND(WX8799, WX8763)
--	WX8801 = AND(WX8343, WX8802)
--	WX8807 = AND(WX8806, WX8763)
--	WX8808 = AND(WX8344, WX8809)
--	WX8814 = AND(WX8813, WX8763)
--	WX8815 = AND(WX8345, WX8816)
--	WX8821 = AND(WX8820, WX8763)
--	WX8822 = AND(WX8346, WX8823)
--	WX8828 = AND(WX8827, WX8763)
--	WX8829 = AND(WX8347, WX8830)
--	WX8835 = AND(WX8834, WX8763)
--	WX8836 = AND(WX8348, WX8837)
--	WX8842 = AND(WX8841, WX8763)
--	WX8843 = AND(WX8349, WX8844)
--	WX8849 = AND(WX8848, WX8763)
--	WX8850 = AND(WX8350, WX8851)
--	WX8856 = AND(WX8855, WX8763)
--	WX8857 = AND(WX8351, WX8858)
--	WX8863 = AND(WX8862, WX8763)
--	WX8864 = AND(WX8352, WX8865)
--	WX8870 = AND(WX8869, WX8763)
--	WX8871 = AND(WX8353, WX8872)
--	WX8877 = AND(WX8876, WX8763)
--	WX8878 = AND(WX8354, WX8879)
--	WX8884 = AND(WX8883, WX8763)
--	WX8885 = AND(WX8355, WX8886)
--	WX8891 = AND(WX8890, WX8763)
--	WX8892 = AND(WX8356, WX8893)
--	WX8898 = AND(WX8897, WX8763)
--	WX8899 = AND(WX8357, WX8900)
--	WX8905 = AND(WX8904, WX8763)
--	WX8906 = AND(WX8358, WX8907)
--	WX8912 = AND(WX8911, WX8763)
--	WX8913 = AND(WX8359, WX8914)
--	WX8919 = AND(WX8918, WX8763)
--	WX8920 = AND(WX8360, WX8921)
--	WX8926 = AND(WX8925, WX8763)
--	WX8927 = AND(WX8361, WX8928)
--	WX8933 = AND(WX8932, WX8763)
--	WX8934 = AND(WX8362, WX8935)
--	WX8940 = AND(WX8939, WX8763)
--	WX8941 = AND(WX8363, WX8942)
--	WX8947 = AND(WX8946, WX8763)
--	WX8948 = AND(WX8364, WX8949)
--	WX8954 = AND(WX8953, WX8763)
--	WX8955 = AND(WX8365, WX8956)
--	WX8961 = AND(WX8960, WX8763)
--	WX8962 = AND(WX8366, WX8963)
--	WX8968 = AND(WX8967, WX8763)
--	WX8969 = AND(WX8367, WX8970)
--	WX8975 = AND(WX8974, WX8763)
--	WX8976 = AND(WX8368, WX8977)
--	WX8982 = AND(WX8981, WX8763)
--	WX8983 = AND(WX8369, WX8984)
--	WX9022 = AND(WX8992, WX9021)
--	WX9024 = AND(WX9020, WX9021)
--	WX9026 = AND(WX9019, WX9021)
--	WX9028 = AND(WX9018, WX9021)
--	WX9030 = AND(WX8991, WX9021)
--	WX9032 = AND(WX9017, WX9021)
--	WX9034 = AND(WX9016, WX9021)
--	WX9036 = AND(WX9015, WX9021)
--	WX9038 = AND(WX9014, WX9021)
--	WX9040 = AND(WX9013, WX9021)
--	WX9042 = AND(WX9012, WX9021)
--	WX9044 = AND(WX8990, WX9021)
--	WX9046 = AND(WX9011, WX9021)
--	WX9048 = AND(WX9010, WX9021)
--	WX9050 = AND(WX9009, WX9021)
--	WX9052 = AND(WX9008, WX9021)
--	WX9054 = AND(WX8989, WX9021)
--	WX9056 = AND(WX9007, WX9021)
--	WX9058 = AND(WX9006, WX9021)
--	WX9060 = AND(WX9005, WX9021)
--	WX9062 = AND(WX9004, WX9021)
--	WX9064 = AND(WX9003, WX9021)
--	WX9066 = AND(WX9002, WX9021)
--	WX9068 = AND(WX9001, WX9021)
--	WX9070 = AND(WX9000, WX9021)
--	WX9072 = AND(WX8999, WX9021)
--	WX9074 = AND(WX8998, WX9021)
--	WX9076 = AND(WX8997, WX9021)
--	WX9078 = AND(WX8996, WX9021)
--	WX9080 = AND(WX8995, WX9021)
--	WX9082 = AND(WX8994, WX9021)
--	WX9084 = AND(WX8993, WX9021)
--	WX9086 = AND(WX9097, WX10054)
--	WX9087 = AND(WX9093, WX9088)
--	WX9090 = AND(CRC_OUT_2_31, WX10055)
--	WX9091 = AND(WX11356, WX9092)
--	WX9094 = AND(WX9536, WX10055)
--	WX9095 = AND(WX10063, WX9096)
--	WX9100 = AND(WX9111, WX10054)
--	WX9101 = AND(WX9107, WX9102)
--	WX9104 = AND(CRC_OUT_2_30, WX10055)
--	WX9105 = AND(WX11363, WX9106)
--	WX9108 = AND(WX9538, WX10055)
--	WX9109 = AND(WX10070, WX9110)
--	WX9114 = AND(WX9125, WX10054)
--	WX9115 = AND(WX9121, WX9116)
--	WX9118 = AND(CRC_OUT_2_29, WX10055)
--	WX9119 = AND(WX11370, WX9120)
--	WX9122 = AND(WX9540, WX10055)
--	WX9123 = AND(WX10077, WX9124)
--	WX9128 = AND(WX9139, WX10054)
--	WX9129 = AND(WX9135, WX9130)
--	WX9132 = AND(CRC_OUT_2_28, WX10055)
--	WX9133 = AND(WX11377, WX9134)
--	WX9136 = AND(WX9542, WX10055)
--	WX9137 = AND(WX10084, WX9138)
--	WX9142 = AND(WX9153, WX10054)
--	WX9143 = AND(WX9149, WX9144)
--	WX9146 = AND(CRC_OUT_2_27, WX10055)
--	WX9147 = AND(WX11384, WX9148)
--	WX9150 = AND(WX9544, WX10055)
--	WX9151 = AND(WX10091, WX9152)
--	WX9156 = AND(WX9167, WX10054)
--	WX9157 = AND(WX9163, WX9158)
--	WX9160 = AND(CRC_OUT_2_26, WX10055)
--	WX9161 = AND(WX11391, WX9162)
--	WX9164 = AND(WX9546, WX10055)
--	WX9165 = AND(WX10098, WX9166)
--	WX9170 = AND(WX9181, WX10054)
--	WX9171 = AND(WX9177, WX9172)
--	WX9174 = AND(CRC_OUT_2_25, WX10055)
--	WX9175 = AND(WX11398, WX9176)
--	WX9178 = AND(WX9548, WX10055)
--	WX9179 = AND(WX10105, WX9180)
--	WX9184 = AND(WX9195, WX10054)
--	WX9185 = AND(WX9191, WX9186)
--	WX9188 = AND(CRC_OUT_2_24, WX10055)
--	WX9189 = AND(WX11405, WX9190)
--	WX9192 = AND(WX9550, WX10055)
--	WX9193 = AND(WX10112, WX9194)
--	WX9198 = AND(WX9209, WX10054)
--	WX9199 = AND(WX9205, WX9200)
--	WX9202 = AND(CRC_OUT_2_23, WX10055)
--	WX9203 = AND(WX11412, WX9204)
--	WX9206 = AND(WX9552, WX10055)
--	WX9207 = AND(WX10119, WX9208)
--	WX9212 = AND(WX9223, WX10054)
--	WX9213 = AND(WX9219, WX9214)
--	WX9216 = AND(CRC_OUT_2_22, WX10055)
--	WX9217 = AND(WX11419, WX9218)
--	WX9220 = AND(WX9554, WX10055)
--	WX9221 = AND(WX10126, WX9222)
--	WX9226 = AND(WX9237, WX10054)
--	WX9227 = AND(WX9233, WX9228)
--	WX9230 = AND(CRC_OUT_2_21, WX10055)
--	WX9231 = AND(WX11426, WX9232)
--	WX9234 = AND(WX9556, WX10055)
--	WX9235 = AND(WX10133, WX9236)
--	WX9240 = AND(WX9251, WX10054)
--	WX9241 = AND(WX9247, WX9242)
--	WX9244 = AND(CRC_OUT_2_20, WX10055)
--	WX9245 = AND(WX11433, WX9246)
--	WX9248 = AND(WX9558, WX10055)
--	WX9249 = AND(WX10140, WX9250)
--	WX9254 = AND(WX9265, WX10054)
--	WX9255 = AND(WX9261, WX9256)
--	WX9258 = AND(CRC_OUT_2_19, WX10055)
--	WX9259 = AND(WX11440, WX9260)
--	WX9262 = AND(WX9560, WX10055)
--	WX9263 = AND(WX10147, WX9264)
--	WX9268 = AND(WX9279, WX10054)
--	WX9269 = AND(WX9275, WX9270)
--	WX9272 = AND(CRC_OUT_2_18, WX10055)
--	WX9273 = AND(WX11447, WX9274)
--	WX9276 = AND(WX9562, WX10055)
--	WX9277 = AND(WX10154, WX9278)
--	WX9282 = AND(WX9293, WX10054)
--	WX9283 = AND(WX9289, WX9284)
--	WX9286 = AND(CRC_OUT_2_17, WX10055)
--	WX9287 = AND(WX11454, WX9288)
--	WX9290 = AND(WX9564, WX10055)
--	WX9291 = AND(WX10161, WX9292)
--	WX9296 = AND(WX9307, WX10054)
--	WX9297 = AND(WX9303, WX9298)
--	WX9300 = AND(CRC_OUT_2_16, WX10055)
--	WX9301 = AND(WX11461, WX9302)
--	WX9304 = AND(WX9566, WX10055)
--	WX9305 = AND(WX10168, WX9306)
--	WX9310 = AND(WX9321, WX10054)
--	WX9311 = AND(WX9317, WX9312)
--	WX9314 = AND(CRC_OUT_2_15, WX10055)
--	WX9315 = AND(WX11468, WX9316)
--	WX9318 = AND(WX9568, WX10055)
--	WX9319 = AND(WX10175, WX9320)
--	WX9324 = AND(WX9335, WX10054)
--	WX9325 = AND(WX9331, WX9326)
--	WX9328 = AND(CRC_OUT_2_14, WX10055)
--	WX9329 = AND(WX11475, WX9330)
--	WX9332 = AND(WX9570, WX10055)
--	WX9333 = AND(WX10182, WX9334)
--	WX9338 = AND(WX9349, WX10054)
--	WX9339 = AND(WX9345, WX9340)
--	WX9342 = AND(CRC_OUT_2_13, WX10055)
--	WX9343 = AND(WX11482, WX9344)
--	WX9346 = AND(WX9572, WX10055)
--	WX9347 = AND(WX10189, WX9348)
--	WX9352 = AND(WX9363, WX10054)
--	WX9353 = AND(WX9359, WX9354)
--	WX9356 = AND(CRC_OUT_2_12, WX10055)
--	WX9357 = AND(WX11489, WX9358)
--	WX9360 = AND(WX9574, WX10055)
--	WX9361 = AND(WX10196, WX9362)
--	WX9366 = AND(WX9377, WX10054)
--	WX9367 = AND(WX9373, WX9368)
--	WX9370 = AND(CRC_OUT_2_11, WX10055)
--	WX9371 = AND(WX11496, WX9372)
--	WX9374 = AND(WX9576, WX10055)
--	WX9375 = AND(WX10203, WX9376)
--	WX9380 = AND(WX9391, WX10054)
--	WX9381 = AND(WX9387, WX9382)
--	WX9384 = AND(CRC_OUT_2_10, WX10055)
--	WX9385 = AND(WX11503, WX9386)
--	WX9388 = AND(WX9578, WX10055)
--	WX9389 = AND(WX10210, WX9390)
--	WX9394 = AND(WX9405, WX10054)
--	WX9395 = AND(WX9401, WX9396)
--	WX9398 = AND(CRC_OUT_2_9, WX10055)
--	WX9399 = AND(WX11510, WX9400)
--	WX9402 = AND(WX9580, WX10055)
--	WX9403 = AND(WX10217, WX9404)
--	WX9408 = AND(WX9419, WX10054)
--	WX9409 = AND(WX9415, WX9410)
--	WX9412 = AND(CRC_OUT_2_8, WX10055)
--	WX9413 = AND(WX11517, WX9414)
--	WX9416 = AND(WX9582, WX10055)
--	WX9417 = AND(WX10224, WX9418)
--	WX9422 = AND(WX9433, WX10054)
--	WX9423 = AND(WX9429, WX9424)
--	WX9426 = AND(CRC_OUT_2_7, WX10055)
--	WX9427 = AND(WX11524, WX9428)
--	WX9430 = AND(WX9584, WX10055)
--	WX9431 = AND(WX10231, WX9432)
--	WX9436 = AND(WX9447, WX10054)
--	WX9437 = AND(WX9443, WX9438)
--	WX9440 = AND(CRC_OUT_2_6, WX10055)
--	WX9441 = AND(WX11531, WX9442)
--	WX9444 = AND(WX9586, WX10055)
--	WX9445 = AND(WX10238, WX9446)
--	WX9450 = AND(WX9461, WX10054)
--	WX9451 = AND(WX9457, WX9452)
--	WX9454 = AND(CRC_OUT_2_5, WX10055)
--	WX9455 = AND(WX11538, WX9456)
--	WX9458 = AND(WX9588, WX10055)
--	WX9459 = AND(WX10245, WX9460)
--	WX9464 = AND(WX9475, WX10054)
--	WX9465 = AND(WX9471, WX9466)
--	WX9468 = AND(CRC_OUT_2_4, WX10055)
--	WX9469 = AND(WX11545, WX9470)
--	WX9472 = AND(WX9590, WX10055)
--	WX9473 = AND(WX10252, WX9474)
--	WX9478 = AND(WX9489, WX10054)
--	WX9479 = AND(WX9485, WX9480)
--	WX9482 = AND(CRC_OUT_2_3, WX10055)
--	WX9483 = AND(WX11552, WX9484)
--	WX9486 = AND(WX9592, WX10055)
--	WX9487 = AND(WX10259, WX9488)
--	WX9492 = AND(WX9503, WX10054)
--	WX9493 = AND(WX9499, WX9494)
--	WX9496 = AND(CRC_OUT_2_2, WX10055)
--	WX9497 = AND(WX11559, WX9498)
--	WX9500 = AND(WX9594, WX10055)
--	WX9501 = AND(WX10266, WX9502)
--	WX9506 = AND(WX9517, WX10054)
--	WX9507 = AND(WX9513, WX9508)
--	WX9510 = AND(CRC_OUT_2_1, WX10055)
--	WX9511 = AND(WX11566, WX9512)
--	WX9514 = AND(WX9596, WX10055)
--	WX9515 = AND(WX10273, WX9516)
--	WX9520 = AND(WX9531, WX10054)
--	WX9521 = AND(WX9527, WX9522)
--	WX9524 = AND(CRC_OUT_2_0, WX10055)
--	WX9525 = AND(WX11573, WX9526)
--	WX9528 = AND(WX9598, WX10055)
--	WX9529 = AND(WX10280, WX9530)
--	WX9535 = AND(WX9538, RESET)
--	WX9537 = AND(WX9540, RESET)
--	WX9539 = AND(WX9542, RESET)
--	WX9541 = AND(WX9544, RESET)
--	WX9543 = AND(WX9546, RESET)
--	WX9545 = AND(WX9548, RESET)
--	WX9547 = AND(WX9550, RESET)
--	WX9549 = AND(WX9552, RESET)
--	WX9551 = AND(WX9554, RESET)
--	WX9553 = AND(WX9556, RESET)
--	WX9555 = AND(WX9558, RESET)
--	WX9557 = AND(WX9560, RESET)
--	WX9559 = AND(WX9562, RESET)
--	WX9561 = AND(WX9564, RESET)
--	WX9563 = AND(WX9566, RESET)
--	WX9565 = AND(WX9568, RESET)
--	WX9567 = AND(WX9570, RESET)
--	WX9569 = AND(WX9572, RESET)
--	WX9571 = AND(WX9574, RESET)
--	WX9573 = AND(WX9576, RESET)
--	WX9575 = AND(WX9578, RESET)
--	WX9577 = AND(WX9580, RESET)
--	WX9579 = AND(WX9582, RESET)
--	WX9581 = AND(WX9584, RESET)
--	WX9583 = AND(WX9586, RESET)
--	WX9585 = AND(WX9588, RESET)
--	WX9587 = AND(WX9590, RESET)
--	WX9589 = AND(WX9592, RESET)
--	WX9591 = AND(WX9594, RESET)
--	WX9593 = AND(WX9596, RESET)
--	WX9595 = AND(WX9598, RESET)
--	WX9597 = AND(WX9534, RESET)
--	WX9695 = AND(WX9099, RESET)
--	WX9697 = AND(WX9113, RESET)
--	WX9699 = AND(WX9127, RESET)
--	WX9701 = AND(WX9141, RESET)
--	WX9703 = AND(WX9155, RESET)
--	WX9705 = AND(WX9169, RESET)
--	WX9707 = AND(WX9183, RESET)
--	WX9709 = AND(WX9197, RESET)
--	WX9711 = AND(WX9211, RESET)
--	WX9713 = AND(WX9225, RESET)
--	WX9715 = AND(WX9239, RESET)
--	WX9717 = AND(WX9253, RESET)
--	WX9719 = AND(WX9267, RESET)
--	WX9721 = AND(WX9281, RESET)
--	WX9723 = AND(WX9295, RESET)
--	WX9725 = AND(WX9309, RESET)
--	WX9727 = AND(WX9323, RESET)
--	WX9729 = AND(WX9337, RESET)
--	WX9731 = AND(WX9351, RESET)
--	WX9733 = AND(WX9365, RESET)
--	WX9735 = AND(WX9379, RESET)
--	WX9737 = AND(WX9393, RESET)
--	WX9739 = AND(WX9407, RESET)
--	WX9741 = AND(WX9421, RESET)
--	WX9743 = AND(WX9435, RESET)
--	WX9745 = AND(WX9449, RESET)
--	WX9747 = AND(WX9463, RESET)
--	WX9749 = AND(WX9477, RESET)
--	WX9751 = AND(WX9491, RESET)
--	WX9753 = AND(WX9505, RESET)
--	WX9755 = AND(WX9519, RESET)
--	WX9757 = AND(WX9533, RESET)
--	WX9759 = AND(WX9696, RESET)
--	WX9761 = AND(WX9698, RESET)
--	WX9763 = AND(WX9700, RESET)
--	WX9765 = AND(WX9702, RESET)
--	WX9767 = AND(WX9704, RESET)
--	WX9769 = AND(WX9706, RESET)
--	WX9771 = AND(WX9708, RESET)
--	WX9773 = AND(WX9710, RESET)
--	WX9775 = AND(WX9712, RESET)
--	WX9777 = AND(WX9714, RESET)
--	WX9779 = AND(WX9716, RESET)
--	WX9781 = AND(WX9718, RESET)
--	WX9783 = AND(WX9720, RESET)
--	WX9785 = AND(WX9722, RESET)
--	WX9787 = AND(WX9724, RESET)
--	WX9789 = AND(WX9726, RESET)
--	WX9791 = AND(WX9728, RESET)
--	WX9793 = AND(WX9730, RESET)
--	WX9795 = AND(WX9732, RESET)
--	WX9797 = AND(WX9734, RESET)
--	WX9799 = AND(WX9736, RESET)
--	WX9801 = AND(WX9738, RESET)
--	WX9803 = AND(WX9740, RESET)
--	WX9805 = AND(WX9742, RESET)
--	WX9807 = AND(WX9744, RESET)
--	WX9809 = AND(WX9746, RESET)
--	WX9811 = AND(WX9748, RESET)
--	WX9813 = AND(WX9750, RESET)
--	WX9815 = AND(WX9752, RESET)
--	WX9817 = AND(WX9754, RESET)
--	WX9819 = AND(WX9756, RESET)
--	WX9821 = AND(WX9758, RESET)
--	WX9823 = AND(WX9760, RESET)
--	WX9825 = AND(WX9762, RESET)
--	WX9827 = AND(WX9764, RESET)
--	WX9829 = AND(WX9766, RESET)
--	WX9831 = AND(WX9768, RESET)
--	WX9833 = AND(WX9770, RESET)
--	WX9835 = AND(WX9772, RESET)
--	WX9837 = AND(WX9774, RESET)
--	WX9839 = AND(WX9776, RESET)
--	WX9841 = AND(WX9778, RESET)
--	WX9843 = AND(WX9780, RESET)
--	WX9845 = AND(WX9782, RESET)
--	WX9847 = AND(WX9784, RESET)
--	WX9849 = AND(WX9786, RESET)
--	WX9851 = AND(WX9788, RESET)
--	WX9853 = AND(WX9790, RESET)
--	WX9855 = AND(WX9792, RESET)
--	WX9857 = AND(WX9794, RESET)
--	WX9859 = AND(WX9796, RESET)
--	WX9861 = AND(WX9798, RESET)
--	WX9863 = AND(WX9800, RESET)
--	WX9865 = AND(WX9802, RESET)
--	WX9867 = AND(WX9804, RESET)
--	WX9869 = AND(WX9806, RESET)
--	WX9871 = AND(WX9808, RESET)
--	WX9873 = AND(WX9810, RESET)
--	WX9875 = AND(WX9812, RESET)
--	WX9877 = AND(WX9814, RESET)
--	WX9879 = AND(WX9816, RESET)
--	WX9881 = AND(WX9818, RESET)
--	WX9883 = AND(WX9820, RESET)
--	WX9885 = AND(WX9822, RESET)
--	WX9887 = AND(WX9824, RESET)
--	WX9889 = AND(WX9826, RESET)
--	WX9891 = AND(WX9828, RESET)
--	WX9893 = AND(WX9830, RESET)
--	WX9895 = AND(WX9832, RESET)
--	WX9897 = AND(WX9834, RESET)
--	WX9899 = AND(WX9836, RESET)
--	WX9901 = AND(WX9838, RESET)
--	WX9903 = AND(WX9840, RESET)
--	WX9905 = AND(WX9842, RESET)
--	WX9907 = AND(WX9844, RESET)
--	WX9909 = AND(WX9846, RESET)
--	WX9911 = AND(WX9848, RESET)
--	WX9913 = AND(WX9850, RESET)
--	WX9915 = AND(WX9852, RESET)
--	WX9917 = AND(WX9854, RESET)
--	WX9919 = AND(WX9856, RESET)
--	WX9921 = AND(WX9858, RESET)
--	WX9923 = AND(WX9860, RESET)
--	WX9925 = AND(WX9862, RESET)
--	WX9927 = AND(WX9864, RESET)
--	WX9929 = AND(WX9866, RESET)
--	WX9931 = AND(WX9868, RESET)
--	WX9933 = AND(WX9870, RESET)
--	WX9935 = AND(WX9872, RESET)
--	WX9937 = AND(WX9874, RESET)
--	WX9939 = AND(WX9876, RESET)
--	WX9941 = AND(WX9878, RESET)
--	WX9943 = AND(WX9880, RESET)
--	WX9945 = AND(WX9882, RESET)
--	WX9947 = AND(WX9884, RESET)
--	WX9949 = AND(WX9886, RESET)
--	WX10058 = AND(WX10057, WX10056)
--	WX10059 = AND(WX9631, WX10060)
--	WX10065 = AND(WX10064, WX10056)
--	WX10066 = AND(WX9632, WX10067)
--	WX10072 = AND(WX10071, WX10056)
--	WX10073 = AND(WX9633, WX10074)
--	WX10079 = AND(WX10078, WX10056)
--	WX10080 = AND(WX9634, WX10081)
--	WX10086 = AND(WX10085, WX10056)
--	WX10087 = AND(WX9635, WX10088)
--	WX10093 = AND(WX10092, WX10056)
--	WX10094 = AND(WX9636, WX10095)
--	WX10100 = AND(WX10099, WX10056)
--	WX10101 = AND(WX9637, WX10102)
--	WX10107 = AND(WX10106, WX10056)
--	WX10108 = AND(WX9638, WX10109)
--	WX10114 = AND(WX10113, WX10056)
--	WX10115 = AND(WX9639, WX10116)
--	WX10121 = AND(WX10120, WX10056)
--	WX10122 = AND(WX9640, WX10123)
--	WX10128 = AND(WX10127, WX10056)
--	WX10129 = AND(WX9641, WX10130)
--	WX10135 = AND(WX10134, WX10056)
--	WX10136 = AND(WX9642, WX10137)
--	WX10142 = AND(WX10141, WX10056)
--	WX10143 = AND(WX9643, WX10144)
--	WX10149 = AND(WX10148, WX10056)
--	WX10150 = AND(WX9644, WX10151)
--	WX10156 = AND(WX10155, WX10056)
--	WX10157 = AND(WX9645, WX10158)
--	WX10163 = AND(WX10162, WX10056)
--	WX10164 = AND(WX9646, WX10165)
--	WX10170 = AND(WX10169, WX10056)
--	WX10171 = AND(WX9647, WX10172)
--	WX10177 = AND(WX10176, WX10056)
--	WX10178 = AND(WX9648, WX10179)
--	WX10184 = AND(WX10183, WX10056)
--	WX10185 = AND(WX9649, WX10186)
--	WX10191 = AND(WX10190, WX10056)
--	WX10192 = AND(WX9650, WX10193)
--	WX10198 = AND(WX10197, WX10056)
--	WX10199 = AND(WX9651, WX10200)
--	WX10205 = AND(WX10204, WX10056)
--	WX10206 = AND(WX9652, WX10207)
--	WX10212 = AND(WX10211, WX10056)
--	WX10213 = AND(WX9653, WX10214)
--	WX10219 = AND(WX10218, WX10056)
--	WX10220 = AND(WX9654, WX10221)
--	WX10226 = AND(WX10225, WX10056)
--	WX10227 = AND(WX9655, WX10228)
--	WX10233 = AND(WX10232, WX10056)
--	WX10234 = AND(WX9656, WX10235)
--	WX10240 = AND(WX10239, WX10056)
--	WX10241 = AND(WX9657, WX10242)
--	WX10247 = AND(WX10246, WX10056)
--	WX10248 = AND(WX9658, WX10249)
--	WX10254 = AND(WX10253, WX10056)
--	WX10255 = AND(WX9659, WX10256)
--	WX10261 = AND(WX10260, WX10056)
--	WX10262 = AND(WX9660, WX10263)
--	WX10268 = AND(WX10267, WX10056)
--	WX10269 = AND(WX9661, WX10270)
--	WX10275 = AND(WX10274, WX10056)
--	WX10276 = AND(WX9662, WX10277)
--	WX10315 = AND(WX10285, WX10314)
--	WX10317 = AND(WX10313, WX10314)
--	WX10319 = AND(WX10312, WX10314)
--	WX10321 = AND(WX10311, WX10314)
--	WX10323 = AND(WX10284, WX10314)
--	WX10325 = AND(WX10310, WX10314)
--	WX10327 = AND(WX10309, WX10314)
--	WX10329 = AND(WX10308, WX10314)
--	WX10331 = AND(WX10307, WX10314)
--	WX10333 = AND(WX10306, WX10314)
--	WX10335 = AND(WX10305, WX10314)
--	WX10337 = AND(WX10283, WX10314)
--	WX10339 = AND(WX10304, WX10314)
--	WX10341 = AND(WX10303, WX10314)
--	WX10343 = AND(WX10302, WX10314)
--	WX10345 = AND(WX10301, WX10314)
--	WX10347 = AND(WX10282, WX10314)
--	WX10349 = AND(WX10300, WX10314)
--	WX10351 = AND(WX10299, WX10314)
--	WX10353 = AND(WX10298, WX10314)
--	WX10355 = AND(WX10297, WX10314)
--	WX10357 = AND(WX10296, WX10314)
--	WX10359 = AND(WX10295, WX10314)
--	WX10361 = AND(WX10294, WX10314)
--	WX10363 = AND(WX10293, WX10314)
--	WX10365 = AND(WX10292, WX10314)
--	WX10367 = AND(WX10291, WX10314)
--	WX10369 = AND(WX10290, WX10314)
--	WX10371 = AND(WX10289, WX10314)
--	WX10373 = AND(WX10288, WX10314)
--	WX10375 = AND(WX10287, WX10314)
--	WX10377 = AND(WX10286, WX10314)
--	WX10379 = AND(WX10390, WX11347)
--	WX10380 = AND(WX10386, WX10381)
--	WX10383 = AND(CRC_OUT_1_31, WX11348)
--	WX10384 = AND(DATA_0_31, WX10385)
--	WX10387 = AND(WX10829, WX11348)
--	WX10388 = AND(WX11356, WX10389)
--	WX10393 = AND(WX10404, WX11347)
--	WX10394 = AND(WX10400, WX10395)
--	WX10397 = AND(CRC_OUT_1_30, WX11348)
--	WX10398 = AND(DATA_0_30, WX10399)
--	WX10401 = AND(WX10831, WX11348)
--	WX10402 = AND(WX11363, WX10403)
--	WX10407 = AND(WX10418, WX11347)
--	WX10408 = AND(WX10414, WX10409)
--	WX10411 = AND(CRC_OUT_1_29, WX11348)
--	WX10412 = AND(DATA_0_29, WX10413)
--	WX10415 = AND(WX10833, WX11348)
--	WX10416 = AND(WX11370, WX10417)
--	WX10421 = AND(WX10432, WX11347)
--	WX10422 = AND(WX10428, WX10423)
--	WX10425 = AND(CRC_OUT_1_28, WX11348)
--	WX10426 = AND(DATA_0_28, WX10427)
--	WX10429 = AND(WX10835, WX11348)
--	WX10430 = AND(WX11377, WX10431)
--	WX10435 = AND(WX10446, WX11347)
--	WX10436 = AND(WX10442, WX10437)
--	WX10439 = AND(CRC_OUT_1_27, WX11348)
--	WX10440 = AND(DATA_0_27, WX10441)
--	WX10443 = AND(WX10837, WX11348)
--	WX10444 = AND(WX11384, WX10445)
--	WX10449 = AND(WX10460, WX11347)
--	WX10450 = AND(WX10456, WX10451)
--	WX10453 = AND(CRC_OUT_1_26, WX11348)
--	WX10454 = AND(DATA_0_26, WX10455)
--	WX10457 = AND(WX10839, WX11348)
--	WX10458 = AND(WX11391, WX10459)
--	WX10463 = AND(WX10474, WX11347)
--	WX10464 = AND(WX10470, WX10465)
--	WX10467 = AND(CRC_OUT_1_25, WX11348)
--	WX10468 = AND(DATA_0_25, WX10469)
--	WX10471 = AND(WX10841, WX11348)
--	WX10472 = AND(WX11398, WX10473)
--	WX10477 = AND(WX10488, WX11347)
--	WX10478 = AND(WX10484, WX10479)
--	WX10481 = AND(CRC_OUT_1_24, WX11348)
--	WX10482 = AND(DATA_0_24, WX10483)
--	WX10485 = AND(WX10843, WX11348)
--	WX10486 = AND(WX11405, WX10487)
--	WX10491 = AND(WX10502, WX11347)
--	WX10492 = AND(WX10498, WX10493)
--	WX10495 = AND(CRC_OUT_1_23, WX11348)
--	WX10496 = AND(DATA_0_23, WX10497)
--	WX10499 = AND(WX10845, WX11348)
--	WX10500 = AND(WX11412, WX10501)
--	WX10505 = AND(WX10516, WX11347)
--	WX10506 = AND(WX10512, WX10507)
--	WX10509 = AND(CRC_OUT_1_22, WX11348)
--	WX10510 = AND(DATA_0_22, WX10511)
--	WX10513 = AND(WX10847, WX11348)
--	WX10514 = AND(WX11419, WX10515)
--	WX10519 = AND(WX10530, WX11347)
--	WX10520 = AND(WX10526, WX10521)
--	WX10523 = AND(CRC_OUT_1_21, WX11348)
--	WX10524 = AND(DATA_0_21, WX10525)
--	WX10527 = AND(WX10849, WX11348)
--	WX10528 = AND(WX11426, WX10529)
--	WX10533 = AND(WX10544, WX11347)
--	WX10534 = AND(WX10540, WX10535)
--	WX10537 = AND(CRC_OUT_1_20, WX11348)
--	WX10538 = AND(DATA_0_20, WX10539)
--	WX10541 = AND(WX10851, WX11348)
--	WX10542 = AND(WX11433, WX10543)
--	WX10547 = AND(WX10558, WX11347)
--	WX10548 = AND(WX10554, WX10549)
--	WX10551 = AND(CRC_OUT_1_19, WX11348)
--	WX10552 = AND(DATA_0_19, WX10553)
--	WX10555 = AND(WX10853, WX11348)
--	WX10556 = AND(WX11440, WX10557)
--	WX10561 = AND(WX10572, WX11347)
--	WX10562 = AND(WX10568, WX10563)
--	WX10565 = AND(CRC_OUT_1_18, WX11348)
--	WX10566 = AND(DATA_0_18, WX10567)
--	WX10569 = AND(WX10855, WX11348)
--	WX10570 = AND(WX11447, WX10571)
--	WX10575 = AND(WX10586, WX11347)
--	WX10576 = AND(WX10582, WX10577)
--	WX10579 = AND(CRC_OUT_1_17, WX11348)
--	WX10580 = AND(DATA_0_17, WX10581)
--	WX10583 = AND(WX10857, WX11348)
--	WX10584 = AND(WX11454, WX10585)
--	WX10589 = AND(WX10600, WX11347)
--	WX10590 = AND(WX10596, WX10591)
--	WX10593 = AND(CRC_OUT_1_16, WX11348)
--	WX10594 = AND(DATA_0_16, WX10595)
--	WX10597 = AND(WX10859, WX11348)
--	WX10598 = AND(WX11461, WX10599)
--	WX10603 = AND(WX10614, WX11347)
--	WX10604 = AND(WX10610, WX10605)
--	WX10607 = AND(CRC_OUT_1_15, WX11348)
--	WX10608 = AND(DATA_0_15, WX10609)
--	WX10611 = AND(WX10861, WX11348)
--	WX10612 = AND(WX11468, WX10613)
--	WX10617 = AND(WX10628, WX11347)
--	WX10618 = AND(WX10624, WX10619)
--	WX10621 = AND(CRC_OUT_1_14, WX11348)
--	WX10622 = AND(DATA_0_14, WX10623)
--	WX10625 = AND(WX10863, WX11348)
--	WX10626 = AND(WX11475, WX10627)
--	WX10631 = AND(WX10642, WX11347)
--	WX10632 = AND(WX10638, WX10633)
--	WX10635 = AND(CRC_OUT_1_13, WX11348)
--	WX10636 = AND(DATA_0_13, WX10637)
--	WX10639 = AND(WX10865, WX11348)
--	WX10640 = AND(WX11482, WX10641)
--	WX10645 = AND(WX10656, WX11347)
--	WX10646 = AND(WX10652, WX10647)
--	WX10649 = AND(CRC_OUT_1_12, WX11348)
--	WX10650 = AND(DATA_0_12, WX10651)
--	WX10653 = AND(WX10867, WX11348)
--	WX10654 = AND(WX11489, WX10655)
--	WX10659 = AND(WX10670, WX11347)
--	WX10660 = AND(WX10666, WX10661)
--	WX10663 = AND(CRC_OUT_1_11, WX11348)
--	WX10664 = AND(DATA_0_11, WX10665)
--	WX10667 = AND(WX10869, WX11348)
--	WX10668 = AND(WX11496, WX10669)
--	WX10673 = AND(WX10684, WX11347)
--	WX10674 = AND(WX10680, WX10675)
--	WX10677 = AND(CRC_OUT_1_10, WX11348)
--	WX10678 = AND(DATA_0_10, WX10679)
--	WX10681 = AND(WX10871, WX11348)
--	WX10682 = AND(WX11503, WX10683)
--	WX10687 = AND(WX10698, WX11347)
--	WX10688 = AND(WX10694, WX10689)
--	WX10691 = AND(CRC_OUT_1_9, WX11348)
--	WX10692 = AND(DATA_0_9, WX10693)
--	WX10695 = AND(WX10873, WX11348)
--	WX10696 = AND(WX11510, WX10697)
--	WX10701 = AND(WX10712, WX11347)
--	WX10702 = AND(WX10708, WX10703)
--	WX10705 = AND(CRC_OUT_1_8, WX11348)
--	WX10706 = AND(DATA_0_8, WX10707)
--	WX10709 = AND(WX10875, WX11348)
--	WX10710 = AND(WX11517, WX10711)
--	WX10715 = AND(WX10726, WX11347)
--	WX10716 = AND(WX10722, WX10717)
--	WX10719 = AND(CRC_OUT_1_7, WX11348)
--	WX10720 = AND(DATA_0_7, WX10721)
--	WX10723 = AND(WX10877, WX11348)
--	WX10724 = AND(WX11524, WX10725)
--	WX10729 = AND(WX10740, WX11347)
--	WX10730 = AND(WX10736, WX10731)
--	WX10733 = AND(CRC_OUT_1_6, WX11348)
--	WX10734 = AND(DATA_0_6, WX10735)
--	WX10737 = AND(WX10879, WX11348)
--	WX10738 = AND(WX11531, WX10739)
--	WX10743 = AND(WX10754, WX11347)
--	WX10744 = AND(WX10750, WX10745)
--	WX10747 = AND(CRC_OUT_1_5, WX11348)
--	WX10748 = AND(DATA_0_5, WX10749)
--	WX10751 = AND(WX10881, WX11348)
--	WX10752 = AND(WX11538, WX10753)
--	WX10757 = AND(WX10768, WX11347)
--	WX10758 = AND(WX10764, WX10759)
--	WX10761 = AND(CRC_OUT_1_4, WX11348)
--	WX10762 = AND(DATA_0_4, WX10763)
--	WX10765 = AND(WX10883, WX11348)
--	WX10766 = AND(WX11545, WX10767)
--	WX10771 = AND(WX10782, WX11347)
--	WX10772 = AND(WX10778, WX10773)
--	WX10775 = AND(CRC_OUT_1_3, WX11348)
--	WX10776 = AND(DATA_0_3, WX10777)
--	WX10779 = AND(WX10885, WX11348)
--	WX10780 = AND(WX11552, WX10781)
--	WX10785 = AND(WX10796, WX11347)
--	WX10786 = AND(WX10792, WX10787)
--	WX10789 = AND(CRC_OUT_1_2, WX11348)
--	WX10790 = AND(DATA_0_2, WX10791)
--	WX10793 = AND(WX10887, WX11348)
--	WX10794 = AND(WX11559, WX10795)
--	WX10799 = AND(WX10810, WX11347)
--	WX10800 = AND(WX10806, WX10801)
--	WX10803 = AND(CRC_OUT_1_1, WX11348)
--	WX10804 = AND(DATA_0_1, WX10805)
--	WX10807 = AND(WX10889, WX11348)
--	WX10808 = AND(WX11566, WX10809)
--	WX10813 = AND(WX10824, WX11347)
--	WX10814 = AND(WX10820, WX10815)
--	WX10817 = AND(CRC_OUT_1_0, WX11348)
--	WX10818 = AND(DATA_0_0, WX10819)
--	WX10821 = AND(WX10891, WX11348)
--	WX10822 = AND(WX11573, WX10823)
--	WX10828 = AND(WX10831, RESET)
--	WX10830 = AND(WX10833, RESET)
--	WX10832 = AND(WX10835, RESET)
--	WX10834 = AND(WX10837, RESET)
--	WX10836 = AND(WX10839, RESET)
--	WX10838 = AND(WX10841, RESET)
--	WX10840 = AND(WX10843, RESET)
--	WX10842 = AND(WX10845, RESET)
--	WX10844 = AND(WX10847, RESET)
--	WX10846 = AND(WX10849, RESET)
--	WX10848 = AND(WX10851, RESET)
--	WX10850 = AND(WX10853, RESET)
--	WX10852 = AND(WX10855, RESET)
--	WX10854 = AND(WX10857, RESET)
--	WX10856 = AND(WX10859, RESET)
--	WX10858 = AND(WX10861, RESET)
--	WX10860 = AND(WX10863, RESET)
--	WX10862 = AND(WX10865, RESET)
--	WX10864 = AND(WX10867, RESET)
--	WX10866 = AND(WX10869, RESET)
--	WX10868 = AND(WX10871, RESET)
--	WX10870 = AND(WX10873, RESET)
--	WX10872 = AND(WX10875, RESET)
--	WX10874 = AND(WX10877, RESET)
--	WX10876 = AND(WX10879, RESET)
--	WX10878 = AND(WX10881, RESET)
--	WX10880 = AND(WX10883, RESET)
--	WX10882 = AND(WX10885, RESET)
--	WX10884 = AND(WX10887, RESET)
--	WX10886 = AND(WX10889, RESET)
--	WX10888 = AND(WX10891, RESET)
--	WX10890 = AND(WX10827, RESET)
--	WX10988 = AND(WX10392, RESET)
--	WX10990 = AND(WX10406, RESET)
--	WX10992 = AND(WX10420, RESET)
--	WX10994 = AND(WX10434, RESET)
--	WX10996 = AND(WX10448, RESET)
--	WX10998 = AND(WX10462, RESET)
--	WX11000 = AND(WX10476, RESET)
--	WX11002 = AND(WX10490, RESET)
--	WX11004 = AND(WX10504, RESET)
--	WX11006 = AND(WX10518, RESET)
--	WX11008 = AND(WX10532, RESET)
--	WX11010 = AND(WX10546, RESET)
--	WX11012 = AND(WX10560, RESET)
--	WX11014 = AND(WX10574, RESET)
--	WX11016 = AND(WX10588, RESET)
--	WX11018 = AND(WX10602, RESET)
--	WX11020 = AND(WX10616, RESET)
--	WX11022 = AND(WX10630, RESET)
--	WX11024 = AND(WX10644, RESET)
--	WX11026 = AND(WX10658, RESET)
--	WX11028 = AND(WX10672, RESET)
--	WX11030 = AND(WX10686, RESET)
--	WX11032 = AND(WX10700, RESET)
--	WX11034 = AND(WX10714, RESET)
--	WX11036 = AND(WX10728, RESET)
--	WX11038 = AND(WX10742, RESET)
--	WX11040 = AND(WX10756, RESET)
--	WX11042 = AND(WX10770, RESET)
--	WX11044 = AND(WX10784, RESET)
--	WX11046 = AND(WX10798, RESET)
--	WX11048 = AND(WX10812, RESET)
--	WX11050 = AND(WX10826, RESET)
--	WX11052 = AND(WX10989, RESET)
--	WX11054 = AND(WX10991, RESET)
--	WX11056 = AND(WX10993, RESET)
--	WX11058 = AND(WX10995, RESET)
--	WX11060 = AND(WX10997, RESET)
--	WX11062 = AND(WX10999, RESET)
--	WX11064 = AND(WX11001, RESET)
--	WX11066 = AND(WX11003, RESET)
--	WX11068 = AND(WX11005, RESET)
--	WX11070 = AND(WX11007, RESET)
--	WX11072 = AND(WX11009, RESET)
--	WX11074 = AND(WX11011, RESET)
--	WX11076 = AND(WX11013, RESET)
--	WX11078 = AND(WX11015, RESET)
--	WX11080 = AND(WX11017, RESET)
--	WX11082 = AND(WX11019, RESET)
--	WX11084 = AND(WX11021, RESET)
--	WX11086 = AND(WX11023, RESET)
--	WX11088 = AND(WX11025, RESET)
--	WX11090 = AND(WX11027, RESET)
--	WX11092 = AND(WX11029, RESET)
--	WX11094 = AND(WX11031, RESET)
--	WX11096 = AND(WX11033, RESET)
--	WX11098 = AND(WX11035, RESET)
--	WX11100 = AND(WX11037, RESET)
--	WX11102 = AND(WX11039, RESET)
--	WX11104 = AND(WX11041, RESET)
--	WX11106 = AND(WX11043, RESET)
--	WX11108 = AND(WX11045, RESET)
--	WX11110 = AND(WX11047, RESET)
--	WX11112 = AND(WX11049, RESET)
--	WX11114 = AND(WX11051, RESET)
--	WX11116 = AND(WX11053, RESET)
--	WX11118 = AND(WX11055, RESET)
--	WX11120 = AND(WX11057, RESET)
--	WX11122 = AND(WX11059, RESET)
--	WX11124 = AND(WX11061, RESET)
--	WX11126 = AND(WX11063, RESET)
--	WX11128 = AND(WX11065, RESET)
--	WX11130 = AND(WX11067, RESET)
--	WX11132 = AND(WX11069, RESET)
--	WX11134 = AND(WX11071, RESET)
--	WX11136 = AND(WX11073, RESET)
--	WX11138 = AND(WX11075, RESET)
--	WX11140 = AND(WX11077, RESET)
--	WX11142 = AND(WX11079, RESET)
--	WX11144 = AND(WX11081, RESET)
--	WX11146 = AND(WX11083, RESET)
--	WX11148 = AND(WX11085, RESET)
--	WX11150 = AND(WX11087, RESET)
--	WX11152 = AND(WX11089, RESET)
--	WX11154 = AND(WX11091, RESET)
--	WX11156 = AND(WX11093, RESET)
--	WX11158 = AND(WX11095, RESET)
--	WX11160 = AND(WX11097, RESET)
--	WX11162 = AND(WX11099, RESET)
--	WX11164 = AND(WX11101, RESET)
--	WX11166 = AND(WX11103, RESET)
--	WX11168 = AND(WX11105, RESET)
--	WX11170 = AND(WX11107, RESET)
--	WX11172 = AND(WX11109, RESET)
--	WX11174 = AND(WX11111, RESET)
--	WX11176 = AND(WX11113, RESET)
--	WX11178 = AND(WX11115, RESET)
--	WX11180 = AND(WX11117, RESET)
--	WX11182 = AND(WX11119, RESET)
--	WX11184 = AND(WX11121, RESET)
--	WX11186 = AND(WX11123, RESET)
--	WX11188 = AND(WX11125, RESET)
--	WX11190 = AND(WX11127, RESET)
--	WX11192 = AND(WX11129, RESET)
--	WX11194 = AND(WX11131, RESET)
--	WX11196 = AND(WX11133, RESET)
--	WX11198 = AND(WX11135, RESET)
--	WX11200 = AND(WX11137, RESET)
--	WX11202 = AND(WX11139, RESET)
--	WX11204 = AND(WX11141, RESET)
--	WX11206 = AND(WX11143, RESET)
--	WX11208 = AND(WX11145, RESET)
--	WX11210 = AND(WX11147, RESET)
--	WX11212 = AND(WX11149, RESET)
--	WX11214 = AND(WX11151, RESET)
--	WX11216 = AND(WX11153, RESET)
--	WX11218 = AND(WX11155, RESET)
--	WX11220 = AND(WX11157, RESET)
--	WX11222 = AND(WX11159, RESET)
--	WX11224 = AND(WX11161, RESET)
--	WX11226 = AND(WX11163, RESET)
--	WX11228 = AND(WX11165, RESET)
--	WX11230 = AND(WX11167, RESET)
--	WX11232 = AND(WX11169, RESET)
--	WX11234 = AND(WX11171, RESET)
--	WX11236 = AND(WX11173, RESET)
--	WX11238 = AND(WX11175, RESET)
--	WX11240 = AND(WX11177, RESET)
--	WX11242 = AND(WX11179, RESET)
--	WX11351 = AND(WX11350, WX11349)
--	WX11352 = AND(WX10924, WX11353)
--	WX11358 = AND(WX11357, WX11349)
--	WX11359 = AND(WX10925, WX11360)
--	WX11365 = AND(WX11364, WX11349)
--	WX11366 = AND(WX10926, WX11367)
--	WX11372 = AND(WX11371, WX11349)
--	WX11373 = AND(WX10927, WX11374)
--	WX11379 = AND(WX11378, WX11349)
--	WX11380 = AND(WX10928, WX11381)
--	WX11386 = AND(WX11385, WX11349)
--	WX11387 = AND(WX10929, WX11388)
--	WX11393 = AND(WX11392, WX11349)
--	WX11394 = AND(WX10930, WX11395)
--	WX11400 = AND(WX11399, WX11349)
--	WX11401 = AND(WX10931, WX11402)
--	WX11407 = AND(WX11406, WX11349)
--	WX11408 = AND(WX10932, WX11409)
--	WX11414 = AND(WX11413, WX11349)
--	WX11415 = AND(WX10933, WX11416)
--	WX11421 = AND(WX11420, WX11349)
--	WX11422 = AND(WX10934, WX11423)
--	WX11428 = AND(WX11427, WX11349)
--	WX11429 = AND(WX10935, WX11430)
--	WX11435 = AND(WX11434, WX11349)
--	WX11436 = AND(WX10936, WX11437)
--	WX11442 = AND(WX11441, WX11349)
--	WX11443 = AND(WX10937, WX11444)
--	WX11449 = AND(WX11448, WX11349)
--	WX11450 = AND(WX10938, WX11451)
--	WX11456 = AND(WX11455, WX11349)
--	WX11457 = AND(WX10939, WX11458)
--	WX11463 = AND(WX11462, WX11349)
--	WX11464 = AND(WX10940, WX11465)
--	WX11470 = AND(WX11469, WX11349)
--	WX11471 = AND(WX10941, WX11472)
--	WX11477 = AND(WX11476, WX11349)
--	WX11478 = AND(WX10942, WX11479)
--	WX11484 = AND(WX11483, WX11349)
--	WX11485 = AND(WX10943, WX11486)
--	WX11491 = AND(WX11490, WX11349)
--	WX11492 = AND(WX10944, WX11493)
--	WX11498 = AND(WX11497, WX11349)
--	WX11499 = AND(WX10945, WX11500)
--	WX11505 = AND(WX11504, WX11349)
--	WX11506 = AND(WX10946, WX11507)
--	WX11512 = AND(WX11511, WX11349)
--	WX11513 = AND(WX10947, WX11514)
--	WX11519 = AND(WX11518, WX11349)
--	WX11520 = AND(WX10948, WX11521)
--	WX11526 = AND(WX11525, WX11349)
--	WX11527 = AND(WX10949, WX11528)
--	WX11533 = AND(WX11532, WX11349)
--	WX11534 = AND(WX10950, WX11535)
--	WX11540 = AND(WX11539, WX11349)
--	WX11541 = AND(WX10951, WX11542)
--	WX11547 = AND(WX11546, WX11349)
--	WX11548 = AND(WX10952, WX11549)
--	WX11554 = AND(WX11553, WX11349)
--	WX11555 = AND(WX10953, WX11556)
--	WX11561 = AND(WX11560, WX11349)
--	WX11562 = AND(WX10954, WX11563)
--	WX11568 = AND(WX11567, WX11349)
--	WX11569 = AND(WX10955, WX11570)
--	WX11608 = AND(WX11578, WX11607)
--	WX11610 = AND(WX11606, WX11607)
--	WX11612 = AND(WX11605, WX11607)
--	WX11614 = AND(WX11604, WX11607)
--	WX11616 = AND(WX11577, WX11607)
--	WX11618 = AND(WX11603, WX11607)
--	WX11620 = AND(WX11602, WX11607)
--	WX11622 = AND(WX11601, WX11607)
--	WX11624 = AND(WX11600, WX11607)
--	WX11626 = AND(WX11599, WX11607)
--	WX11628 = AND(WX11598, WX11607)
--	WX11630 = AND(WX11576, WX11607)
--	WX11632 = AND(WX11597, WX11607)
--	WX11634 = AND(WX11596, WX11607)
--	WX11636 = AND(WX11595, WX11607)
--	WX11638 = AND(WX11594, WX11607)
--	WX11640 = AND(WX11575, WX11607)
--	WX11642 = AND(WX11593, WX11607)
--	WX11644 = AND(WX11592, WX11607)
--	WX11646 = AND(WX11591, WX11607)
--	WX11648 = AND(WX11590, WX11607)
--	WX11650 = AND(WX11589, WX11607)
--	WX11652 = AND(WX11588, WX11607)
--	WX11654 = AND(WX11587, WX11607)
--	WX11656 = AND(WX11586, WX11607)
--	WX11658 = AND(WX11585, WX11607)
--	WX11660 = AND(WX11584, WX11607)
--	WX11662 = AND(WX11583, WX11607)
--	WX11664 = AND(WX11582, WX11607)
--	WX11666 = AND(WX11581, WX11607)
--	WX11668 = AND(WX11580, WX11607)
--	WX11670 = AND(WX11579, WX11607)
--	
--	WX38 = OR(WX36, WX35)
--	WX42 = OR(WX40, WX39)
--	WX46 = OR(WX44, WX43)
--	WX52 = OR(WX50, WX49)
--	WX56 = OR(WX54, WX53)
--	WX60 = OR(WX58, WX57)
--	WX66 = OR(WX64, WX63)
--	WX70 = OR(WX68, WX67)
--	WX74 = OR(WX72, WX71)
--	WX80 = OR(WX78, WX77)
--	WX84 = OR(WX82, WX81)
--	WX88 = OR(WX86, WX85)
--	WX94 = OR(WX92, WX91)
--	WX98 = OR(WX96, WX95)
--	WX102 = OR(WX100, WX99)
--	WX108 = OR(WX106, WX105)
--	WX112 = OR(WX110, WX109)
--	WX116 = OR(WX114, WX113)
--	WX122 = OR(WX120, WX119)
--	WX126 = OR(WX124, WX123)
--	WX130 = OR(WX128, WX127)
--	WX136 = OR(WX134, WX133)
--	WX140 = OR(WX138, WX137)
--	WX144 = OR(WX142, WX141)
--	WX150 = OR(WX148, WX147)
--	WX154 = OR(WX152, WX151)
--	WX158 = OR(WX156, WX155)
--	WX164 = OR(WX162, WX161)
--	WX168 = OR(WX166, WX165)
--	WX172 = OR(WX170, WX169)
--	WX178 = OR(WX176, WX175)
--	WX182 = OR(WX180, WX179)
--	WX186 = OR(WX184, WX183)
--	WX192 = OR(WX190, WX189)
--	WX196 = OR(WX194, WX193)
--	WX200 = OR(WX198, WX197)
--	WX206 = OR(WX204, WX203)
--	WX210 = OR(WX208, WX207)
--	WX214 = OR(WX212, WX211)
--	WX220 = OR(WX218, WX217)
--	WX224 = OR(WX222, WX221)
--	WX228 = OR(WX226, WX225)
--	WX234 = OR(WX232, WX231)
--	WX238 = OR(WX236, WX235)
--	WX242 = OR(WX240, WX239)
--	WX248 = OR(WX246, WX245)
--	WX252 = OR(WX250, WX249)
--	WX256 = OR(WX254, WX253)
--	WX262 = OR(WX260, WX259)
--	WX266 = OR(WX264, WX263)
--	WX270 = OR(WX268, WX267)
--	WX276 = OR(WX274, WX273)
--	WX280 = OR(WX278, WX277)
--	WX284 = OR(WX282, WX281)
--	WX290 = OR(WX288, WX287)
--	WX294 = OR(WX292, WX291)
--	WX298 = OR(WX296, WX295)
--	WX304 = OR(WX302, WX301)
--	WX308 = OR(WX306, WX305)
--	WX312 = OR(WX310, WX309)
--	WX318 = OR(WX316, WX315)
--	WX322 = OR(WX320, WX319)
--	WX326 = OR(WX324, WX323)
--	WX332 = OR(WX330, WX329)
--	WX336 = OR(WX334, WX333)
--	WX340 = OR(WX338, WX337)
--	WX346 = OR(WX344, WX343)
--	WX350 = OR(WX348, WX347)
--	WX354 = OR(WX352, WX351)
--	WX360 = OR(WX358, WX357)
--	WX364 = OR(WX362, WX361)
--	WX368 = OR(WX366, WX365)
--	WX374 = OR(WX372, WX371)
--	WX378 = OR(WX376, WX375)
--	WX382 = OR(WX380, WX379)
--	WX388 = OR(WX386, WX385)
--	WX392 = OR(WX390, WX389)
--	WX396 = OR(WX394, WX393)
--	WX402 = OR(WX400, WX399)
--	WX406 = OR(WX404, WX403)
--	WX410 = OR(WX408, WX407)
--	WX416 = OR(WX414, WX413)
--	WX420 = OR(WX418, WX417)
--	WX424 = OR(WX422, WX421)
--	WX430 = OR(WX428, WX427)
--	WX434 = OR(WX432, WX431)
--	WX438 = OR(WX436, WX435)
--	WX444 = OR(WX442, WX441)
--	WX448 = OR(WX446, WX445)
--	WX452 = OR(WX450, WX449)
--	WX458 = OR(WX456, WX455)
--	WX462 = OR(WX460, WX459)
--	WX466 = OR(WX464, WX463)
--	WX472 = OR(WX470, WX469)
--	WX476 = OR(WX474, WX473)
--	WX480 = OR(WX478, WX477)
--	WX1010 = OR(WX1008, WX1007)
--	WX1017 = OR(WX1015, WX1014)
--	WX1024 = OR(WX1022, WX1021)
--	WX1031 = OR(WX1029, WX1028)
--	WX1038 = OR(WX1036, WX1035)
--	WX1045 = OR(WX1043, WX1042)
--	WX1052 = OR(WX1050, WX1049)
--	WX1059 = OR(WX1057, WX1056)
--	WX1066 = OR(WX1064, WX1063)
--	WX1073 = OR(WX1071, WX1070)
--	WX1080 = OR(WX1078, WX1077)
--	WX1087 = OR(WX1085, WX1084)
--	WX1094 = OR(WX1092, WX1091)
--	WX1101 = OR(WX1099, WX1098)
--	WX1108 = OR(WX1106, WX1105)
--	WX1115 = OR(WX1113, WX1112)
--	WX1122 = OR(WX1120, WX1119)
--	WX1129 = OR(WX1127, WX1126)
--	WX1136 = OR(WX1134, WX1133)
--	WX1143 = OR(WX1141, WX1140)
--	WX1150 = OR(WX1148, WX1147)
--	WX1157 = OR(WX1155, WX1154)
--	WX1164 = OR(WX1162, WX1161)
--	WX1171 = OR(WX1169, WX1168)
--	WX1178 = OR(WX1176, WX1175)
--	WX1185 = OR(WX1183, WX1182)
--	WX1192 = OR(WX1190, WX1189)
--	WX1199 = OR(WX1197, WX1196)
--	WX1206 = OR(WX1204, WX1203)
--	WX1213 = OR(WX1211, WX1210)
--	WX1220 = OR(WX1218, WX1217)
--	WX1227 = OR(WX1225, WX1224)
--	WX1331 = OR(WX1329, WX1328)
--	WX1335 = OR(WX1333, WX1332)
--	WX1339 = OR(WX1337, WX1336)
--	WX1345 = OR(WX1343, WX1342)
--	WX1349 = OR(WX1347, WX1346)
--	WX1353 = OR(WX1351, WX1350)
--	WX1359 = OR(WX1357, WX1356)
--	WX1363 = OR(WX1361, WX1360)
--	WX1367 = OR(WX1365, WX1364)
--	WX1373 = OR(WX1371, WX1370)
--	WX1377 = OR(WX1375, WX1374)
--	WX1381 = OR(WX1379, WX1378)
--	WX1387 = OR(WX1385, WX1384)
--	WX1391 = OR(WX1389, WX1388)
--	WX1395 = OR(WX1393, WX1392)
--	WX1401 = OR(WX1399, WX1398)
--	WX1405 = OR(WX1403, WX1402)
--	WX1409 = OR(WX1407, WX1406)
--	WX1415 = OR(WX1413, WX1412)
--	WX1419 = OR(WX1417, WX1416)
--	WX1423 = OR(WX1421, WX1420)
--	WX1429 = OR(WX1427, WX1426)
--	WX1433 = OR(WX1431, WX1430)
--	WX1437 = OR(WX1435, WX1434)
--	WX1443 = OR(WX1441, WX1440)
--	WX1447 = OR(WX1445, WX1444)
--	WX1451 = OR(WX1449, WX1448)
--	WX1457 = OR(WX1455, WX1454)
--	WX1461 = OR(WX1459, WX1458)
--	WX1465 = OR(WX1463, WX1462)
--	WX1471 = OR(WX1469, WX1468)
--	WX1475 = OR(WX1473, WX1472)
--	WX1479 = OR(WX1477, WX1476)
--	WX1485 = OR(WX1483, WX1482)
--	WX1489 = OR(WX1487, WX1486)
--	WX1493 = OR(WX1491, WX1490)
--	WX1499 = OR(WX1497, WX1496)
--	WX1503 = OR(WX1501, WX1500)
--	WX1507 = OR(WX1505, WX1504)
--	WX1513 = OR(WX1511, WX1510)
--	WX1517 = OR(WX1515, WX1514)
--	WX1521 = OR(WX1519, WX1518)
--	WX1527 = OR(WX1525, WX1524)
--	WX1531 = OR(WX1529, WX1528)
--	WX1535 = OR(WX1533, WX1532)
--	WX1541 = OR(WX1539, WX1538)
--	WX1545 = OR(WX1543, WX1542)
--	WX1549 = OR(WX1547, WX1546)
--	WX1555 = OR(WX1553, WX1552)
--	WX1559 = OR(WX1557, WX1556)
--	WX1563 = OR(WX1561, WX1560)
--	WX1569 = OR(WX1567, WX1566)
--	WX1573 = OR(WX1571, WX1570)
--	WX1577 = OR(WX1575, WX1574)
--	WX1583 = OR(WX1581, WX1580)
--	WX1587 = OR(WX1585, WX1584)
--	WX1591 = OR(WX1589, WX1588)
--	WX1597 = OR(WX1595, WX1594)
--	WX1601 = OR(WX1599, WX1598)
--	WX1605 = OR(WX1603, WX1602)
--	WX1611 = OR(WX1609, WX1608)
--	WX1615 = OR(WX1613, WX1612)
--	WX1619 = OR(WX1617, WX1616)
--	WX1625 = OR(WX1623, WX1622)
--	WX1629 = OR(WX1627, WX1626)
--	WX1633 = OR(WX1631, WX1630)
--	WX1639 = OR(WX1637, WX1636)
--	WX1643 = OR(WX1641, WX1640)
--	WX1647 = OR(WX1645, WX1644)
--	WX1653 = OR(WX1651, WX1650)
--	WX1657 = OR(WX1655, WX1654)
--	WX1661 = OR(WX1659, WX1658)
--	WX1667 = OR(WX1665, WX1664)
--	WX1671 = OR(WX1669, WX1668)
--	WX1675 = OR(WX1673, WX1672)
--	WX1681 = OR(WX1679, WX1678)
--	WX1685 = OR(WX1683, WX1682)
--	WX1689 = OR(WX1687, WX1686)
--	WX1695 = OR(WX1693, WX1692)
--	WX1699 = OR(WX1697, WX1696)
--	WX1703 = OR(WX1701, WX1700)
--	WX1709 = OR(WX1707, WX1706)
--	WX1713 = OR(WX1711, WX1710)
--	WX1717 = OR(WX1715, WX1714)
--	WX1723 = OR(WX1721, WX1720)
--	WX1727 = OR(WX1725, WX1724)
--	WX1731 = OR(WX1729, WX1728)
--	WX1737 = OR(WX1735, WX1734)
--	WX1741 = OR(WX1739, WX1738)
--	WX1745 = OR(WX1743, WX1742)
--	WX1751 = OR(WX1749, WX1748)
--	WX1755 = OR(WX1753, WX1752)
--	WX1759 = OR(WX1757, WX1756)
--	WX1765 = OR(WX1763, WX1762)
--	WX1769 = OR(WX1767, WX1766)
--	WX1773 = OR(WX1771, WX1770)
--	WX2303 = OR(WX2301, WX2300)
--	WX2310 = OR(WX2308, WX2307)
--	WX2317 = OR(WX2315, WX2314)
--	WX2324 = OR(WX2322, WX2321)
--	WX2331 = OR(WX2329, WX2328)
--	WX2338 = OR(WX2336, WX2335)
--	WX2345 = OR(WX2343, WX2342)
--	WX2352 = OR(WX2350, WX2349)
--	WX2359 = OR(WX2357, WX2356)
--	WX2366 = OR(WX2364, WX2363)
--	WX2373 = OR(WX2371, WX2370)
--	WX2380 = OR(WX2378, WX2377)
--	WX2387 = OR(WX2385, WX2384)
--	WX2394 = OR(WX2392, WX2391)
--	WX2401 = OR(WX2399, WX2398)
--	WX2408 = OR(WX2406, WX2405)
--	WX2415 = OR(WX2413, WX2412)
--	WX2422 = OR(WX2420, WX2419)
--	WX2429 = OR(WX2427, WX2426)
--	WX2436 = OR(WX2434, WX2433)
--	WX2443 = OR(WX2441, WX2440)
--	WX2450 = OR(WX2448, WX2447)
--	WX2457 = OR(WX2455, WX2454)
--	WX2464 = OR(WX2462, WX2461)
--	WX2471 = OR(WX2469, WX2468)
--	WX2478 = OR(WX2476, WX2475)
--	WX2485 = OR(WX2483, WX2482)
--	WX2492 = OR(WX2490, WX2489)
--	WX2499 = OR(WX2497, WX2496)
--	WX2506 = OR(WX2504, WX2503)
--	WX2513 = OR(WX2511, WX2510)
--	WX2520 = OR(WX2518, WX2517)
--	WX2624 = OR(WX2622, WX2621)
--	WX2628 = OR(WX2626, WX2625)
--	WX2632 = OR(WX2630, WX2629)
--	WX2638 = OR(WX2636, WX2635)
--	WX2642 = OR(WX2640, WX2639)
--	WX2646 = OR(WX2644, WX2643)
--	WX2652 = OR(WX2650, WX2649)
--	WX2656 = OR(WX2654, WX2653)
--	WX2660 = OR(WX2658, WX2657)
--	WX2666 = OR(WX2664, WX2663)
--	WX2670 = OR(WX2668, WX2667)
--	WX2674 = OR(WX2672, WX2671)
--	WX2680 = OR(WX2678, WX2677)
--	WX2684 = OR(WX2682, WX2681)
--	WX2688 = OR(WX2686, WX2685)
--	WX2694 = OR(WX2692, WX2691)
--	WX2698 = OR(WX2696, WX2695)
--	WX2702 = OR(WX2700, WX2699)
--	WX2708 = OR(WX2706, WX2705)
--	WX2712 = OR(WX2710, WX2709)
--	WX2716 = OR(WX2714, WX2713)
--	WX2722 = OR(WX2720, WX2719)
--	WX2726 = OR(WX2724, WX2723)
--	WX2730 = OR(WX2728, WX2727)
--	WX2736 = OR(WX2734, WX2733)
--	WX2740 = OR(WX2738, WX2737)
--	WX2744 = OR(WX2742, WX2741)
--	WX2750 = OR(WX2748, WX2747)
--	WX2754 = OR(WX2752, WX2751)
--	WX2758 = OR(WX2756, WX2755)
--	WX2764 = OR(WX2762, WX2761)
--	WX2768 = OR(WX2766, WX2765)
--	WX2772 = OR(WX2770, WX2769)
--	WX2778 = OR(WX2776, WX2775)
--	WX2782 = OR(WX2780, WX2779)
--	WX2786 = OR(WX2784, WX2783)
--	WX2792 = OR(WX2790, WX2789)
--	WX2796 = OR(WX2794, WX2793)
--	WX2800 = OR(WX2798, WX2797)
--	WX2806 = OR(WX2804, WX2803)
--	WX2810 = OR(WX2808, WX2807)
--	WX2814 = OR(WX2812, WX2811)
--	WX2820 = OR(WX2818, WX2817)
--	WX2824 = OR(WX2822, WX2821)
--	WX2828 = OR(WX2826, WX2825)
--	WX2834 = OR(WX2832, WX2831)
--	WX2838 = OR(WX2836, WX2835)
--	WX2842 = OR(WX2840, WX2839)
--	WX2848 = OR(WX2846, WX2845)
--	WX2852 = OR(WX2850, WX2849)
--	WX2856 = OR(WX2854, WX2853)
--	WX2862 = OR(WX2860, WX2859)
--	WX2866 = OR(WX2864, WX2863)
--	WX2870 = OR(WX2868, WX2867)
--	WX2876 = OR(WX2874, WX2873)
--	WX2880 = OR(WX2878, WX2877)
--	WX2884 = OR(WX2882, WX2881)
--	WX2890 = OR(WX2888, WX2887)
--	WX2894 = OR(WX2892, WX2891)
--	WX2898 = OR(WX2896, WX2895)
--	WX2904 = OR(WX2902, WX2901)
--	WX2908 = OR(WX2906, WX2905)
--	WX2912 = OR(WX2910, WX2909)
--	WX2918 = OR(WX2916, WX2915)
--	WX2922 = OR(WX2920, WX2919)
--	WX2926 = OR(WX2924, WX2923)
--	WX2932 = OR(WX2930, WX2929)
--	WX2936 = OR(WX2934, WX2933)
--	WX2940 = OR(WX2938, WX2937)
--	WX2946 = OR(WX2944, WX2943)
--	WX2950 = OR(WX2948, WX2947)
--	WX2954 = OR(WX2952, WX2951)
--	WX2960 = OR(WX2958, WX2957)
--	WX2964 = OR(WX2962, WX2961)
--	WX2968 = OR(WX2966, WX2965)
--	WX2974 = OR(WX2972, WX2971)
--	WX2978 = OR(WX2976, WX2975)
--	WX2982 = OR(WX2980, WX2979)
--	WX2988 = OR(WX2986, WX2985)
--	WX2992 = OR(WX2990, WX2989)
--	WX2996 = OR(WX2994, WX2993)
--	WX3002 = OR(WX3000, WX2999)
--	WX3006 = OR(WX3004, WX3003)
--	WX3010 = OR(WX3008, WX3007)
--	WX3016 = OR(WX3014, WX3013)
--	WX3020 = OR(WX3018, WX3017)
--	WX3024 = OR(WX3022, WX3021)
--	WX3030 = OR(WX3028, WX3027)
--	WX3034 = OR(WX3032, WX3031)
--	WX3038 = OR(WX3036, WX3035)
--	WX3044 = OR(WX3042, WX3041)
--	WX3048 = OR(WX3046, WX3045)
--	WX3052 = OR(WX3050, WX3049)
--	WX3058 = OR(WX3056, WX3055)
--	WX3062 = OR(WX3060, WX3059)
--	WX3066 = OR(WX3064, WX3063)
--	WX3596 = OR(WX3594, WX3593)
--	WX3603 = OR(WX3601, WX3600)
--	WX3610 = OR(WX3608, WX3607)
--	WX3617 = OR(WX3615, WX3614)
--	WX3624 = OR(WX3622, WX3621)
--	WX3631 = OR(WX3629, WX3628)
--	WX3638 = OR(WX3636, WX3635)
--	WX3645 = OR(WX3643, WX3642)
--	WX3652 = OR(WX3650, WX3649)
--	WX3659 = OR(WX3657, WX3656)
--	WX3666 = OR(WX3664, WX3663)
--	WX3673 = OR(WX3671, WX3670)
--	WX3680 = OR(WX3678, WX3677)
--	WX3687 = OR(WX3685, WX3684)
--	WX3694 = OR(WX3692, WX3691)
--	WX3701 = OR(WX3699, WX3698)
--	WX3708 = OR(WX3706, WX3705)
--	WX3715 = OR(WX3713, WX3712)
--	WX3722 = OR(WX3720, WX3719)
--	WX3729 = OR(WX3727, WX3726)
--	WX3736 = OR(WX3734, WX3733)
--	WX3743 = OR(WX3741, WX3740)
--	WX3750 = OR(WX3748, WX3747)
--	WX3757 = OR(WX3755, WX3754)
--	WX3764 = OR(WX3762, WX3761)
--	WX3771 = OR(WX3769, WX3768)
--	WX3778 = OR(WX3776, WX3775)
--	WX3785 = OR(WX3783, WX3782)
--	WX3792 = OR(WX3790, WX3789)
--	WX3799 = OR(WX3797, WX3796)
--	WX3806 = OR(WX3804, WX3803)
--	WX3813 = OR(WX3811, WX3810)
--	WX3917 = OR(WX3915, WX3914)
--	WX3921 = OR(WX3919, WX3918)
--	WX3925 = OR(WX3923, WX3922)
--	WX3931 = OR(WX3929, WX3928)
--	WX3935 = OR(WX3933, WX3932)
--	WX3939 = OR(WX3937, WX3936)
--	WX3945 = OR(WX3943, WX3942)
--	WX3949 = OR(WX3947, WX3946)
--	WX3953 = OR(WX3951, WX3950)
--	WX3959 = OR(WX3957, WX3956)
--	WX3963 = OR(WX3961, WX3960)
--	WX3967 = OR(WX3965, WX3964)
--	WX3973 = OR(WX3971, WX3970)
--	WX3977 = OR(WX3975, WX3974)
--	WX3981 = OR(WX3979, WX3978)
--	WX3987 = OR(WX3985, WX3984)
--	WX3991 = OR(WX3989, WX3988)
--	WX3995 = OR(WX3993, WX3992)
--	WX4001 = OR(WX3999, WX3998)
--	WX4005 = OR(WX4003, WX4002)
--	WX4009 = OR(WX4007, WX4006)
--	WX4015 = OR(WX4013, WX4012)
--	WX4019 = OR(WX4017, WX4016)
--	WX4023 = OR(WX4021, WX4020)
--	WX4029 = OR(WX4027, WX4026)
--	WX4033 = OR(WX4031, WX4030)
--	WX4037 = OR(WX4035, WX4034)
--	WX4043 = OR(WX4041, WX4040)
--	WX4047 = OR(WX4045, WX4044)
--	WX4051 = OR(WX4049, WX4048)
--	WX4057 = OR(WX4055, WX4054)
--	WX4061 = OR(WX4059, WX4058)
--	WX4065 = OR(WX4063, WX4062)
--	WX4071 = OR(WX4069, WX4068)
--	WX4075 = OR(WX4073, WX4072)
--	WX4079 = OR(WX4077, WX4076)
--	WX4085 = OR(WX4083, WX4082)
--	WX4089 = OR(WX4087, WX4086)
--	WX4093 = OR(WX4091, WX4090)
--	WX4099 = OR(WX4097, WX4096)
--	WX4103 = OR(WX4101, WX4100)
--	WX4107 = OR(WX4105, WX4104)
--	WX4113 = OR(WX4111, WX4110)
--	WX4117 = OR(WX4115, WX4114)
--	WX4121 = OR(WX4119, WX4118)
--	WX4127 = OR(WX4125, WX4124)
--	WX4131 = OR(WX4129, WX4128)
--	WX4135 = OR(WX4133, WX4132)
--	WX4141 = OR(WX4139, WX4138)
--	WX4145 = OR(WX4143, WX4142)
--	WX4149 = OR(WX4147, WX4146)
--	WX4155 = OR(WX4153, WX4152)
--	WX4159 = OR(WX4157, WX4156)
--	WX4163 = OR(WX4161, WX4160)
--	WX4169 = OR(WX4167, WX4166)
--	WX4173 = OR(WX4171, WX4170)
--	WX4177 = OR(WX4175, WX4174)
--	WX4183 = OR(WX4181, WX4180)
--	WX4187 = OR(WX4185, WX4184)
--	WX4191 = OR(WX4189, WX4188)
--	WX4197 = OR(WX4195, WX4194)
--	WX4201 = OR(WX4199, WX4198)
--	WX4205 = OR(WX4203, WX4202)
--	WX4211 = OR(WX4209, WX4208)
--	WX4215 = OR(WX4213, WX4212)
--	WX4219 = OR(WX4217, WX4216)
--	WX4225 = OR(WX4223, WX4222)
--	WX4229 = OR(WX4227, WX4226)
--	WX4233 = OR(WX4231, WX4230)
--	WX4239 = OR(WX4237, WX4236)
--	WX4243 = OR(WX4241, WX4240)
--	WX4247 = OR(WX4245, WX4244)
--	WX4253 = OR(WX4251, WX4250)
--	WX4257 = OR(WX4255, WX4254)
--	WX4261 = OR(WX4259, WX4258)
--	WX4267 = OR(WX4265, WX4264)
--	WX4271 = OR(WX4269, WX4268)
--	WX4275 = OR(WX4273, WX4272)
--	WX4281 = OR(WX4279, WX4278)
--	WX4285 = OR(WX4283, WX4282)
--	WX4289 = OR(WX4287, WX4286)
--	WX4295 = OR(WX4293, WX4292)
--	WX4299 = OR(WX4297, WX4296)
--	WX4303 = OR(WX4301, WX4300)
--	WX4309 = OR(WX4307, WX4306)
--	WX4313 = OR(WX4311, WX4310)
--	WX4317 = OR(WX4315, WX4314)
--	WX4323 = OR(WX4321, WX4320)
--	WX4327 = OR(WX4325, WX4324)
--	WX4331 = OR(WX4329, WX4328)
--	WX4337 = OR(WX4335, WX4334)
--	WX4341 = OR(WX4339, WX4338)
--	WX4345 = OR(WX4343, WX4342)
--	WX4351 = OR(WX4349, WX4348)
--	WX4355 = OR(WX4353, WX4352)
--	WX4359 = OR(WX4357, WX4356)
--	WX4889 = OR(WX4887, WX4886)
--	WX4896 = OR(WX4894, WX4893)
--	WX4903 = OR(WX4901, WX4900)
--	WX4910 = OR(WX4908, WX4907)
--	WX4917 = OR(WX4915, WX4914)
--	WX4924 = OR(WX4922, WX4921)
--	WX4931 = OR(WX4929, WX4928)
--	WX4938 = OR(WX4936, WX4935)
--	WX4945 = OR(WX4943, WX4942)
--	WX4952 = OR(WX4950, WX4949)
--	WX4959 = OR(WX4957, WX4956)
--	WX4966 = OR(WX4964, WX4963)
--	WX4973 = OR(WX4971, WX4970)
--	WX4980 = OR(WX4978, WX4977)
--	WX4987 = OR(WX4985, WX4984)
--	WX4994 = OR(WX4992, WX4991)
--	WX5001 = OR(WX4999, WX4998)
--	WX5008 = OR(WX5006, WX5005)
--	WX5015 = OR(WX5013, WX5012)
--	WX5022 = OR(WX5020, WX5019)
--	WX5029 = OR(WX5027, WX5026)
--	WX5036 = OR(WX5034, WX5033)
--	WX5043 = OR(WX5041, WX5040)
--	WX5050 = OR(WX5048, WX5047)
--	WX5057 = OR(WX5055, WX5054)
--	WX5064 = OR(WX5062, WX5061)
--	WX5071 = OR(WX5069, WX5068)
--	WX5078 = OR(WX5076, WX5075)
--	WX5085 = OR(WX5083, WX5082)
--	WX5092 = OR(WX5090, WX5089)
--	WX5099 = OR(WX5097, WX5096)
--	WX5106 = OR(WX5104, WX5103)
--	WX5210 = OR(WX5208, WX5207)
--	WX5214 = OR(WX5212, WX5211)
--	WX5218 = OR(WX5216, WX5215)
--	WX5224 = OR(WX5222, WX5221)
--	WX5228 = OR(WX5226, WX5225)
--	WX5232 = OR(WX5230, WX5229)
--	WX5238 = OR(WX5236, WX5235)
--	WX5242 = OR(WX5240, WX5239)
--	WX5246 = OR(WX5244, WX5243)
--	WX5252 = OR(WX5250, WX5249)
--	WX5256 = OR(WX5254, WX5253)
--	WX5260 = OR(WX5258, WX5257)
--	WX5266 = OR(WX5264, WX5263)
--	WX5270 = OR(WX5268, WX5267)
--	WX5274 = OR(WX5272, WX5271)
--	WX5280 = OR(WX5278, WX5277)
--	WX5284 = OR(WX5282, WX5281)
--	WX5288 = OR(WX5286, WX5285)
--	WX5294 = OR(WX5292, WX5291)
--	WX5298 = OR(WX5296, WX5295)
--	WX5302 = OR(WX5300, WX5299)
--	WX5308 = OR(WX5306, WX5305)
--	WX5312 = OR(WX5310, WX5309)
--	WX5316 = OR(WX5314, WX5313)
--	WX5322 = OR(WX5320, WX5319)
--	WX5326 = OR(WX5324, WX5323)
--	WX5330 = OR(WX5328, WX5327)
--	WX5336 = OR(WX5334, WX5333)
--	WX5340 = OR(WX5338, WX5337)
--	WX5344 = OR(WX5342, WX5341)
--	WX5350 = OR(WX5348, WX5347)
--	WX5354 = OR(WX5352, WX5351)
--	WX5358 = OR(WX5356, WX5355)
--	WX5364 = OR(WX5362, WX5361)
--	WX5368 = OR(WX5366, WX5365)
--	WX5372 = OR(WX5370, WX5369)
--	WX5378 = OR(WX5376, WX5375)
--	WX5382 = OR(WX5380, WX5379)
--	WX5386 = OR(WX5384, WX5383)
--	WX5392 = OR(WX5390, WX5389)
--	WX5396 = OR(WX5394, WX5393)
--	WX5400 = OR(WX5398, WX5397)
--	WX5406 = OR(WX5404, WX5403)
--	WX5410 = OR(WX5408, WX5407)
--	WX5414 = OR(WX5412, WX5411)
--	WX5420 = OR(WX5418, WX5417)
--	WX5424 = OR(WX5422, WX5421)
--	WX5428 = OR(WX5426, WX5425)
--	WX5434 = OR(WX5432, WX5431)
--	WX5438 = OR(WX5436, WX5435)
--	WX5442 = OR(WX5440, WX5439)
--	WX5448 = OR(WX5446, WX5445)
--	WX5452 = OR(WX5450, WX5449)
--	WX5456 = OR(WX5454, WX5453)
--	WX5462 = OR(WX5460, WX5459)
--	WX5466 = OR(WX5464, WX5463)
--	WX5470 = OR(WX5468, WX5467)
--	WX5476 = OR(WX5474, WX5473)
--	WX5480 = OR(WX5478, WX5477)
--	WX5484 = OR(WX5482, WX5481)
--	WX5490 = OR(WX5488, WX5487)
--	WX5494 = OR(WX5492, WX5491)
--	WX5498 = OR(WX5496, WX5495)
--	WX5504 = OR(WX5502, WX5501)
--	WX5508 = OR(WX5506, WX5505)
--	WX5512 = OR(WX5510, WX5509)
--	WX5518 = OR(WX5516, WX5515)
--	WX5522 = OR(WX5520, WX5519)
--	WX5526 = OR(WX5524, WX5523)
--	WX5532 = OR(WX5530, WX5529)
--	WX5536 = OR(WX5534, WX5533)
--	WX5540 = OR(WX5538, WX5537)
--	WX5546 = OR(WX5544, WX5543)
--	WX5550 = OR(WX5548, WX5547)
--	WX5554 = OR(WX5552, WX5551)
--	WX5560 = OR(WX5558, WX5557)
--	WX5564 = OR(WX5562, WX5561)
--	WX5568 = OR(WX5566, WX5565)
--	WX5574 = OR(WX5572, WX5571)
--	WX5578 = OR(WX5576, WX5575)
--	WX5582 = OR(WX5580, WX5579)
--	WX5588 = OR(WX5586, WX5585)
--	WX5592 = OR(WX5590, WX5589)
--	WX5596 = OR(WX5594, WX5593)
--	WX5602 = OR(WX5600, WX5599)
--	WX5606 = OR(WX5604, WX5603)
--	WX5610 = OR(WX5608, WX5607)
--	WX5616 = OR(WX5614, WX5613)
--	WX5620 = OR(WX5618, WX5617)
--	WX5624 = OR(WX5622, WX5621)
--	WX5630 = OR(WX5628, WX5627)
--	WX5634 = OR(WX5632, WX5631)
--	WX5638 = OR(WX5636, WX5635)
--	WX5644 = OR(WX5642, WX5641)
--	WX5648 = OR(WX5646, WX5645)
--	WX5652 = OR(WX5650, WX5649)
--	WX6182 = OR(WX6180, WX6179)
--	WX6189 = OR(WX6187, WX6186)
--	WX6196 = OR(WX6194, WX6193)
--	WX6203 = OR(WX6201, WX6200)
--	WX6210 = OR(WX6208, WX6207)
--	WX6217 = OR(WX6215, WX6214)
--	WX6224 = OR(WX6222, WX6221)
--	WX6231 = OR(WX6229, WX6228)
--	WX6238 = OR(WX6236, WX6235)
--	WX6245 = OR(WX6243, WX6242)
--	WX6252 = OR(WX6250, WX6249)
--	WX6259 = OR(WX6257, WX6256)
--	WX6266 = OR(WX6264, WX6263)
--	WX6273 = OR(WX6271, WX6270)
--	WX6280 = OR(WX6278, WX6277)
--	WX6287 = OR(WX6285, WX6284)
--	WX6294 = OR(WX6292, WX6291)
--	WX6301 = OR(WX6299, WX6298)
--	WX6308 = OR(WX6306, WX6305)
--	WX6315 = OR(WX6313, WX6312)
--	WX6322 = OR(WX6320, WX6319)
--	WX6329 = OR(WX6327, WX6326)
--	WX6336 = OR(WX6334, WX6333)
--	WX6343 = OR(WX6341, WX6340)
--	WX6350 = OR(WX6348, WX6347)
--	WX6357 = OR(WX6355, WX6354)
--	WX6364 = OR(WX6362, WX6361)
--	WX6371 = OR(WX6369, WX6368)
--	WX6378 = OR(WX6376, WX6375)
--	WX6385 = OR(WX6383, WX6382)
--	WX6392 = OR(WX6390, WX6389)
--	WX6399 = OR(WX6397, WX6396)
--	WX6503 = OR(WX6501, WX6500)
--	WX6507 = OR(WX6505, WX6504)
--	WX6511 = OR(WX6509, WX6508)
--	WX6517 = OR(WX6515, WX6514)
--	WX6521 = OR(WX6519, WX6518)
--	WX6525 = OR(WX6523, WX6522)
--	WX6531 = OR(WX6529, WX6528)
--	WX6535 = OR(WX6533, WX6532)
--	WX6539 = OR(WX6537, WX6536)
--	WX6545 = OR(WX6543, WX6542)
--	WX6549 = OR(WX6547, WX6546)
--	WX6553 = OR(WX6551, WX6550)
--	WX6559 = OR(WX6557, WX6556)
--	WX6563 = OR(WX6561, WX6560)
--	WX6567 = OR(WX6565, WX6564)
--	WX6573 = OR(WX6571, WX6570)
--	WX6577 = OR(WX6575, WX6574)
--	WX6581 = OR(WX6579, WX6578)
--	WX6587 = OR(WX6585, WX6584)
--	WX6591 = OR(WX6589, WX6588)
--	WX6595 = OR(WX6593, WX6592)
--	WX6601 = OR(WX6599, WX6598)
--	WX6605 = OR(WX6603, WX6602)
--	WX6609 = OR(WX6607, WX6606)
--	WX6615 = OR(WX6613, WX6612)
--	WX6619 = OR(WX6617, WX6616)
--	WX6623 = OR(WX6621, WX6620)
--	WX6629 = OR(WX6627, WX6626)
--	WX6633 = OR(WX6631, WX6630)
--	WX6637 = OR(WX6635, WX6634)
--	WX6643 = OR(WX6641, WX6640)
--	WX6647 = OR(WX6645, WX6644)
--	WX6651 = OR(WX6649, WX6648)
--	WX6657 = OR(WX6655, WX6654)
--	WX6661 = OR(WX6659, WX6658)
--	WX6665 = OR(WX6663, WX6662)
--	WX6671 = OR(WX6669, WX6668)
--	WX6675 = OR(WX6673, WX6672)
--	WX6679 = OR(WX6677, WX6676)
--	WX6685 = OR(WX6683, WX6682)
--	WX6689 = OR(WX6687, WX6686)
--	WX6693 = OR(WX6691, WX6690)
--	WX6699 = OR(WX6697, WX6696)
--	WX6703 = OR(WX6701, WX6700)
--	WX6707 = OR(WX6705, WX6704)
--	WX6713 = OR(WX6711, WX6710)
--	WX6717 = OR(WX6715, WX6714)
--	WX6721 = OR(WX6719, WX6718)
--	WX6727 = OR(WX6725, WX6724)
--	WX6731 = OR(WX6729, WX6728)
--	WX6735 = OR(WX6733, WX6732)
--	WX6741 = OR(WX6739, WX6738)
--	WX6745 = OR(WX6743, WX6742)
--	WX6749 = OR(WX6747, WX6746)
--	WX6755 = OR(WX6753, WX6752)
--	WX6759 = OR(WX6757, WX6756)
--	WX6763 = OR(WX6761, WX6760)
--	WX6769 = OR(WX6767, WX6766)
--	WX6773 = OR(WX6771, WX6770)
--	WX6777 = OR(WX6775, WX6774)
--	WX6783 = OR(WX6781, WX6780)
--	WX6787 = OR(WX6785, WX6784)
--	WX6791 = OR(WX6789, WX6788)
--	WX6797 = OR(WX6795, WX6794)
--	WX6801 = OR(WX6799, WX6798)
--	WX6805 = OR(WX6803, WX6802)
--	WX6811 = OR(WX6809, WX6808)
--	WX6815 = OR(WX6813, WX6812)
--	WX6819 = OR(WX6817, WX6816)
--	WX6825 = OR(WX6823, WX6822)
--	WX6829 = OR(WX6827, WX6826)
--	WX6833 = OR(WX6831, WX6830)
--	WX6839 = OR(WX6837, WX6836)
--	WX6843 = OR(WX6841, WX6840)
--	WX6847 = OR(WX6845, WX6844)
--	WX6853 = OR(WX6851, WX6850)
--	WX6857 = OR(WX6855, WX6854)
--	WX6861 = OR(WX6859, WX6858)
--	WX6867 = OR(WX6865, WX6864)
--	WX6871 = OR(WX6869, WX6868)
--	WX6875 = OR(WX6873, WX6872)
--	WX6881 = OR(WX6879, WX6878)
--	WX6885 = OR(WX6883, WX6882)
--	WX6889 = OR(WX6887, WX6886)
--	WX6895 = OR(WX6893, WX6892)
--	WX6899 = OR(WX6897, WX6896)
--	WX6903 = OR(WX6901, WX6900)
--	WX6909 = OR(WX6907, WX6906)
--	WX6913 = OR(WX6911, WX6910)
--	WX6917 = OR(WX6915, WX6914)
--	WX6923 = OR(WX6921, WX6920)
--	WX6927 = OR(WX6925, WX6924)
--	WX6931 = OR(WX6929, WX6928)
--	WX6937 = OR(WX6935, WX6934)
--	WX6941 = OR(WX6939, WX6938)
--	WX6945 = OR(WX6943, WX6942)
--	WX7475 = OR(WX7473, WX7472)
--	WX7482 = OR(WX7480, WX7479)
--	WX7489 = OR(WX7487, WX7486)
--	WX7496 = OR(WX7494, WX7493)
--	WX7503 = OR(WX7501, WX7500)
--	WX7510 = OR(WX7508, WX7507)
--	WX7517 = OR(WX7515, WX7514)
--	WX7524 = OR(WX7522, WX7521)
--	WX7531 = OR(WX7529, WX7528)
--	WX7538 = OR(WX7536, WX7535)
--	WX7545 = OR(WX7543, WX7542)
--	WX7552 = OR(WX7550, WX7549)
--	WX7559 = OR(WX7557, WX7556)
--	WX7566 = OR(WX7564, WX7563)
--	WX7573 = OR(WX7571, WX7570)
--	WX7580 = OR(WX7578, WX7577)
--	WX7587 = OR(WX7585, WX7584)
--	WX7594 = OR(WX7592, WX7591)
--	WX7601 = OR(WX7599, WX7598)
--	WX7608 = OR(WX7606, WX7605)
--	WX7615 = OR(WX7613, WX7612)
--	WX7622 = OR(WX7620, WX7619)
--	WX7629 = OR(WX7627, WX7626)
--	WX7636 = OR(WX7634, WX7633)
--	WX7643 = OR(WX7641, WX7640)
--	WX7650 = OR(WX7648, WX7647)
--	WX7657 = OR(WX7655, WX7654)
--	WX7664 = OR(WX7662, WX7661)
--	WX7671 = OR(WX7669, WX7668)
--	WX7678 = OR(WX7676, WX7675)
--	WX7685 = OR(WX7683, WX7682)
--	WX7692 = OR(WX7690, WX7689)
--	WX7796 = OR(WX7794, WX7793)
--	WX7800 = OR(WX7798, WX7797)
--	WX7804 = OR(WX7802, WX7801)
--	WX7810 = OR(WX7808, WX7807)
--	WX7814 = OR(WX7812, WX7811)
--	WX7818 = OR(WX7816, WX7815)
--	WX7824 = OR(WX7822, WX7821)
--	WX7828 = OR(WX7826, WX7825)
--	WX7832 = OR(WX7830, WX7829)
--	WX7838 = OR(WX7836, WX7835)
--	WX7842 = OR(WX7840, WX7839)
--	WX7846 = OR(WX7844, WX7843)
--	WX7852 = OR(WX7850, WX7849)
--	WX7856 = OR(WX7854, WX7853)
--	WX7860 = OR(WX7858, WX7857)
--	WX7866 = OR(WX7864, WX7863)
--	WX7870 = OR(WX7868, WX7867)
--	WX7874 = OR(WX7872, WX7871)
--	WX7880 = OR(WX7878, WX7877)
--	WX7884 = OR(WX7882, WX7881)
--	WX7888 = OR(WX7886, WX7885)
--	WX7894 = OR(WX7892, WX7891)
--	WX7898 = OR(WX7896, WX7895)
--	WX7902 = OR(WX7900, WX7899)
--	WX7908 = OR(WX7906, WX7905)
--	WX7912 = OR(WX7910, WX7909)
--	WX7916 = OR(WX7914, WX7913)
--	WX7922 = OR(WX7920, WX7919)
--	WX7926 = OR(WX7924, WX7923)
--	WX7930 = OR(WX7928, WX7927)
--	WX7936 = OR(WX7934, WX7933)
--	WX7940 = OR(WX7938, WX7937)
--	WX7944 = OR(WX7942, WX7941)
--	WX7950 = OR(WX7948, WX7947)
--	WX7954 = OR(WX7952, WX7951)
--	WX7958 = OR(WX7956, WX7955)
--	WX7964 = OR(WX7962, WX7961)
--	WX7968 = OR(WX7966, WX7965)
--	WX7972 = OR(WX7970, WX7969)
--	WX7978 = OR(WX7976, WX7975)
--	WX7982 = OR(WX7980, WX7979)
--	WX7986 = OR(WX7984, WX7983)
--	WX7992 = OR(WX7990, WX7989)
--	WX7996 = OR(WX7994, WX7993)
--	WX8000 = OR(WX7998, WX7997)
--	WX8006 = OR(WX8004, WX8003)
--	WX8010 = OR(WX8008, WX8007)
--	WX8014 = OR(WX8012, WX8011)
--	WX8020 = OR(WX8018, WX8017)
--	WX8024 = OR(WX8022, WX8021)
--	WX8028 = OR(WX8026, WX8025)
--	WX8034 = OR(WX8032, WX8031)
--	WX8038 = OR(WX8036, WX8035)
--	WX8042 = OR(WX8040, WX8039)
--	WX8048 = OR(WX8046, WX8045)
--	WX8052 = OR(WX8050, WX8049)
--	WX8056 = OR(WX8054, WX8053)
--	WX8062 = OR(WX8060, WX8059)
--	WX8066 = OR(WX8064, WX8063)
--	WX8070 = OR(WX8068, WX8067)
--	WX8076 = OR(WX8074, WX8073)
--	WX8080 = OR(WX8078, WX8077)
--	WX8084 = OR(WX8082, WX8081)
--	WX8090 = OR(WX8088, WX8087)
--	WX8094 = OR(WX8092, WX8091)
--	WX8098 = OR(WX8096, WX8095)
--	WX8104 = OR(WX8102, WX8101)
--	WX8108 = OR(WX8106, WX8105)
--	WX8112 = OR(WX8110, WX8109)
--	WX8118 = OR(WX8116, WX8115)
--	WX8122 = OR(WX8120, WX8119)
--	WX8126 = OR(WX8124, WX8123)
--	WX8132 = OR(WX8130, WX8129)
--	WX8136 = OR(WX8134, WX8133)
--	WX8140 = OR(WX8138, WX8137)
--	WX8146 = OR(WX8144, WX8143)
--	WX8150 = OR(WX8148, WX8147)
--	WX8154 = OR(WX8152, WX8151)
--	WX8160 = OR(WX8158, WX8157)
--	WX8164 = OR(WX8162, WX8161)
--	WX8168 = OR(WX8166, WX8165)
--	WX8174 = OR(WX8172, WX8171)
--	WX8178 = OR(WX8176, WX8175)
--	WX8182 = OR(WX8180, WX8179)
--	WX8188 = OR(WX8186, WX8185)
--	WX8192 = OR(WX8190, WX8189)
--	WX8196 = OR(WX8194, WX8193)
--	WX8202 = OR(WX8200, WX8199)
--	WX8206 = OR(WX8204, WX8203)
--	WX8210 = OR(WX8208, WX8207)
--	WX8216 = OR(WX8214, WX8213)
--	WX8220 = OR(WX8218, WX8217)
--	WX8224 = OR(WX8222, WX8221)
--	WX8230 = OR(WX8228, WX8227)
--	WX8234 = OR(WX8232, WX8231)
--	WX8238 = OR(WX8236, WX8235)
--	WX8768 = OR(WX8766, WX8765)
--	WX8775 = OR(WX8773, WX8772)
--	WX8782 = OR(WX8780, WX8779)
--	WX8789 = OR(WX8787, WX8786)
--	WX8796 = OR(WX8794, WX8793)
--	WX8803 = OR(WX8801, WX8800)
--	WX8810 = OR(WX8808, WX8807)
--	WX8817 = OR(WX8815, WX8814)
--	WX8824 = OR(WX8822, WX8821)
--	WX8831 = OR(WX8829, WX8828)
--	WX8838 = OR(WX8836, WX8835)
--	WX8845 = OR(WX8843, WX8842)
--	WX8852 = OR(WX8850, WX8849)
--	WX8859 = OR(WX8857, WX8856)
--	WX8866 = OR(WX8864, WX8863)
--	WX8873 = OR(WX8871, WX8870)
--	WX8880 = OR(WX8878, WX8877)
--	WX8887 = OR(WX8885, WX8884)
--	WX8894 = OR(WX8892, WX8891)
--	WX8901 = OR(WX8899, WX8898)
--	WX8908 = OR(WX8906, WX8905)
--	WX8915 = OR(WX8913, WX8912)
--	WX8922 = OR(WX8920, WX8919)
--	WX8929 = OR(WX8927, WX8926)
--	WX8936 = OR(WX8934, WX8933)
--	WX8943 = OR(WX8941, WX8940)
--	WX8950 = OR(WX8948, WX8947)
--	WX8957 = OR(WX8955, WX8954)
--	WX8964 = OR(WX8962, WX8961)
--	WX8971 = OR(WX8969, WX8968)
--	WX8978 = OR(WX8976, WX8975)
--	WX8985 = OR(WX8983, WX8982)
--	WX9089 = OR(WX9087, WX9086)
--	WX9093 = OR(WX9091, WX9090)
--	WX9097 = OR(WX9095, WX9094)
--	WX9103 = OR(WX9101, WX9100)
--	WX9107 = OR(WX9105, WX9104)
--	WX9111 = OR(WX9109, WX9108)
--	WX9117 = OR(WX9115, WX9114)
--	WX9121 = OR(WX9119, WX9118)
--	WX9125 = OR(WX9123, WX9122)
--	WX9131 = OR(WX9129, WX9128)
--	WX9135 = OR(WX9133, WX9132)
--	WX9139 = OR(WX9137, WX9136)
--	WX9145 = OR(WX9143, WX9142)
--	WX9149 = OR(WX9147, WX9146)
--	WX9153 = OR(WX9151, WX9150)
--	WX9159 = OR(WX9157, WX9156)
--	WX9163 = OR(WX9161, WX9160)
--	WX9167 = OR(WX9165, WX9164)
--	WX9173 = OR(WX9171, WX9170)
--	WX9177 = OR(WX9175, WX9174)
--	WX9181 = OR(WX9179, WX9178)
--	WX9187 = OR(WX9185, WX9184)
--	WX9191 = OR(WX9189, WX9188)
--	WX9195 = OR(WX9193, WX9192)
--	WX9201 = OR(WX9199, WX9198)
--	WX9205 = OR(WX9203, WX9202)
--	WX9209 = OR(WX9207, WX9206)
--	WX9215 = OR(WX9213, WX9212)
--	WX9219 = OR(WX9217, WX9216)
--	WX9223 = OR(WX9221, WX9220)
--	WX9229 = OR(WX9227, WX9226)
--	WX9233 = OR(WX9231, WX9230)
--	WX9237 = OR(WX9235, WX9234)
--	WX9243 = OR(WX9241, WX9240)
--	WX9247 = OR(WX9245, WX9244)
--	WX9251 = OR(WX9249, WX9248)
--	WX9257 = OR(WX9255, WX9254)
--	WX9261 = OR(WX9259, WX9258)
--	WX9265 = OR(WX9263, WX9262)
--	WX9271 = OR(WX9269, WX9268)
--	WX9275 = OR(WX9273, WX9272)
--	WX9279 = OR(WX9277, WX9276)
--	WX9285 = OR(WX9283, WX9282)
--	WX9289 = OR(WX9287, WX9286)
--	WX9293 = OR(WX9291, WX9290)
--	WX9299 = OR(WX9297, WX9296)
--	WX9303 = OR(WX9301, WX9300)
--	WX9307 = OR(WX9305, WX9304)
--	WX9313 = OR(WX9311, WX9310)
--	WX9317 = OR(WX9315, WX9314)
--	WX9321 = OR(WX9319, WX9318)
--	WX9327 = OR(WX9325, WX9324)
--	WX9331 = OR(WX9329, WX9328)
--	WX9335 = OR(WX9333, WX9332)
--	WX9341 = OR(WX9339, WX9338)
--	WX9345 = OR(WX9343, WX9342)
--	WX9349 = OR(WX9347, WX9346)
--	WX9355 = OR(WX9353, WX9352)
--	WX9359 = OR(WX9357, WX9356)
--	WX9363 = OR(WX9361, WX9360)
--	WX9369 = OR(WX9367, WX9366)
--	WX9373 = OR(WX9371, WX9370)
--	WX9377 = OR(WX9375, WX9374)
--	WX9383 = OR(WX9381, WX9380)
--	WX9387 = OR(WX9385, WX9384)
--	WX9391 = OR(WX9389, WX9388)
--	WX9397 = OR(WX9395, WX9394)
--	WX9401 = OR(WX9399, WX9398)
--	WX9405 = OR(WX9403, WX9402)
--	WX9411 = OR(WX9409, WX9408)
--	WX9415 = OR(WX9413, WX9412)
--	WX9419 = OR(WX9417, WX9416)
--	WX9425 = OR(WX9423, WX9422)
--	WX9429 = OR(WX9427, WX9426)
--	WX9433 = OR(WX9431, WX9430)
--	WX9439 = OR(WX9437, WX9436)
--	WX9443 = OR(WX9441, WX9440)
--	WX9447 = OR(WX9445, WX9444)
--	WX9453 = OR(WX9451, WX9450)
--	WX9457 = OR(WX9455, WX9454)
--	WX9461 = OR(WX9459, WX9458)
--	WX9467 = OR(WX9465, WX9464)
--	WX9471 = OR(WX9469, WX9468)
--	WX9475 = OR(WX9473, WX9472)
--	WX9481 = OR(WX9479, WX9478)
--	WX9485 = OR(WX9483, WX9482)
--	WX9489 = OR(WX9487, WX9486)
--	WX9495 = OR(WX9493, WX9492)
--	WX9499 = OR(WX9497, WX9496)
--	WX9503 = OR(WX9501, WX9500)
--	WX9509 = OR(WX9507, WX9506)
--	WX9513 = OR(WX9511, WX9510)
--	WX9517 = OR(WX9515, WX9514)
--	WX9523 = OR(WX9521, WX9520)
--	WX9527 = OR(WX9525, WX9524)
--	WX9531 = OR(WX9529, WX9528)
--	WX10061 = OR(WX10059, WX10058)
--	WX10068 = OR(WX10066, WX10065)
--	WX10075 = OR(WX10073, WX10072)
--	WX10082 = OR(WX10080, WX10079)
--	WX10089 = OR(WX10087, WX10086)
--	WX10096 = OR(WX10094, WX10093)
--	WX10103 = OR(WX10101, WX10100)
--	WX10110 = OR(WX10108, WX10107)
--	WX10117 = OR(WX10115, WX10114)
--	WX10124 = OR(WX10122, WX10121)
--	WX10131 = OR(WX10129, WX10128)
--	WX10138 = OR(WX10136, WX10135)
--	WX10145 = OR(WX10143, WX10142)
--	WX10152 = OR(WX10150, WX10149)
--	WX10159 = OR(WX10157, WX10156)
--	WX10166 = OR(WX10164, WX10163)
--	WX10173 = OR(WX10171, WX10170)
--	WX10180 = OR(WX10178, WX10177)
--	WX10187 = OR(WX10185, WX10184)
--	WX10194 = OR(WX10192, WX10191)
--	WX10201 = OR(WX10199, WX10198)
--	WX10208 = OR(WX10206, WX10205)
--	WX10215 = OR(WX10213, WX10212)
--	WX10222 = OR(WX10220, WX10219)
--	WX10229 = OR(WX10227, WX10226)
--	WX10236 = OR(WX10234, WX10233)
--	WX10243 = OR(WX10241, WX10240)
--	WX10250 = OR(WX10248, WX10247)
--	WX10257 = OR(WX10255, WX10254)
--	WX10264 = OR(WX10262, WX10261)
--	WX10271 = OR(WX10269, WX10268)
--	WX10278 = OR(WX10276, WX10275)
--	WX10382 = OR(WX10380, WX10379)
--	WX10386 = OR(WX10384, WX10383)
--	WX10390 = OR(WX10388, WX10387)
--	WX10396 = OR(WX10394, WX10393)
--	WX10400 = OR(WX10398, WX10397)
--	WX10404 = OR(WX10402, WX10401)
--	WX10410 = OR(WX10408, WX10407)
--	WX10414 = OR(WX10412, WX10411)
--	WX10418 = OR(WX10416, WX10415)
--	WX10424 = OR(WX10422, WX10421)
--	WX10428 = OR(WX10426, WX10425)
--	WX10432 = OR(WX10430, WX10429)
--	WX10438 = OR(WX10436, WX10435)
--	WX10442 = OR(WX10440, WX10439)
--	WX10446 = OR(WX10444, WX10443)
--	WX10452 = OR(WX10450, WX10449)
--	WX10456 = OR(WX10454, WX10453)
--	WX10460 = OR(WX10458, WX10457)
--	WX10466 = OR(WX10464, WX10463)
--	WX10470 = OR(WX10468, WX10467)
--	WX10474 = OR(WX10472, WX10471)
--	WX10480 = OR(WX10478, WX10477)
--	WX10484 = OR(WX10482, WX10481)
--	WX10488 = OR(WX10486, WX10485)
--	WX10494 = OR(WX10492, WX10491)
--	WX10498 = OR(WX10496, WX10495)
--	WX10502 = OR(WX10500, WX10499)
--	WX10508 = OR(WX10506, WX10505)
--	WX10512 = OR(WX10510, WX10509)
--	WX10516 = OR(WX10514, WX10513)
--	WX10522 = OR(WX10520, WX10519)
--	WX10526 = OR(WX10524, WX10523)
--	WX10530 = OR(WX10528, WX10527)
--	WX10536 = OR(WX10534, WX10533)
--	WX10540 = OR(WX10538, WX10537)
--	WX10544 = OR(WX10542, WX10541)
--	WX10550 = OR(WX10548, WX10547)
--	WX10554 = OR(WX10552, WX10551)
--	WX10558 = OR(WX10556, WX10555)
--	WX10564 = OR(WX10562, WX10561)
--	WX10568 = OR(WX10566, WX10565)
--	WX10572 = OR(WX10570, WX10569)
--	WX10578 = OR(WX10576, WX10575)
--	WX10582 = OR(WX10580, WX10579)
--	WX10586 = OR(WX10584, WX10583)
--	WX10592 = OR(WX10590, WX10589)
--	WX10596 = OR(WX10594, WX10593)
--	WX10600 = OR(WX10598, WX10597)
--	WX10606 = OR(WX10604, WX10603)
--	WX10610 = OR(WX10608, WX10607)
--	WX10614 = OR(WX10612, WX10611)
--	WX10620 = OR(WX10618, WX10617)
--	WX10624 = OR(WX10622, WX10621)
--	WX10628 = OR(WX10626, WX10625)
--	WX10634 = OR(WX10632, WX10631)
--	WX10638 = OR(WX10636, WX10635)
--	WX10642 = OR(WX10640, WX10639)
--	WX10648 = OR(WX10646, WX10645)
--	WX10652 = OR(WX10650, WX10649)
--	WX10656 = OR(WX10654, WX10653)
--	WX10662 = OR(WX10660, WX10659)
--	WX10666 = OR(WX10664, WX10663)
--	WX10670 = OR(WX10668, WX10667)
--	WX10676 = OR(WX10674, WX10673)
--	WX10680 = OR(WX10678, WX10677)
--	WX10684 = OR(WX10682, WX10681)
--	WX10690 = OR(WX10688, WX10687)
--	WX10694 = OR(WX10692, WX10691)
--	WX10698 = OR(WX10696, WX10695)
--	WX10704 = OR(WX10702, WX10701)
--	WX10708 = OR(WX10706, WX10705)
--	WX10712 = OR(WX10710, WX10709)
--	WX10718 = OR(WX10716, WX10715)
--	WX10722 = OR(WX10720, WX10719)
--	WX10726 = OR(WX10724, WX10723)
--	WX10732 = OR(WX10730, WX10729)
--	WX10736 = OR(WX10734, WX10733)
--	WX10740 = OR(WX10738, WX10737)
--	WX10746 = OR(WX10744, WX10743)
--	WX10750 = OR(WX10748, WX10747)
--	WX10754 = OR(WX10752, WX10751)
--	WX10760 = OR(WX10758, WX10757)
--	WX10764 = OR(WX10762, WX10761)
--	WX10768 = OR(WX10766, WX10765)
--	WX10774 = OR(WX10772, WX10771)
--	WX10778 = OR(WX10776, WX10775)
--	WX10782 = OR(WX10780, WX10779)
--	WX10788 = OR(WX10786, WX10785)
--	WX10792 = OR(WX10790, WX10789)
--	WX10796 = OR(WX10794, WX10793)
--	WX10802 = OR(WX10800, WX10799)
--	WX10806 = OR(WX10804, WX10803)
--	WX10810 = OR(WX10808, WX10807)
--	WX10816 = OR(WX10814, WX10813)
--	WX10820 = OR(WX10818, WX10817)
--	WX10824 = OR(WX10822, WX10821)
--	WX11354 = OR(WX11352, WX11351)
--	WX11361 = OR(WX11359, WX11358)
--	WX11368 = OR(WX11366, WX11365)
--	WX11375 = OR(WX11373, WX11372)
--	WX11382 = OR(WX11380, WX11379)
--	WX11389 = OR(WX11387, WX11386)
--	WX11396 = OR(WX11394, WX11393)
--	WX11403 = OR(WX11401, WX11400)
--	WX11410 = OR(WX11408, WX11407)
--	WX11417 = OR(WX11415, WX11414)
--	WX11424 = OR(WX11422, WX11421)
--	WX11431 = OR(WX11429, WX11428)
--	WX11438 = OR(WX11436, WX11435)
--	WX11445 = OR(WX11443, WX11442)
--	WX11452 = OR(WX11450, WX11449)
--	WX11459 = OR(WX11457, WX11456)
--	WX11466 = OR(WX11464, WX11463)
--	WX11473 = OR(WX11471, WX11470)
--	WX11480 = OR(WX11478, WX11477)
--	WX11487 = OR(WX11485, WX11484)
--	WX11494 = OR(WX11492, WX11491)
--	WX11501 = OR(WX11499, WX11498)
--	WX11508 = OR(WX11506, WX11505)
--	WX11515 = OR(WX11513, WX11512)
--	WX11522 = OR(WX11520, WX11519)
--	WX11529 = OR(WX11527, WX11526)
--	WX11536 = OR(WX11534, WX11533)
--	WX11543 = OR(WX11541, WX11540)
--	WX11550 = OR(WX11548, WX11547)
--	WX11557 = OR(WX11555, WX11554)
--	WX11564 = OR(WX11562, WX11561)
--	WX11571 = OR(WX11569, WX11568)
--	
--	I1988 = NAND(WX1001, WX645)
--	I1989 = NAND(WX1001, I1988)
--	I1990 = NAND(WX645, I1988)
--	I1987 = NAND(I1989, I1990)
--	I1995 = NAND(WX709, I1987)
--	I1996 = NAND(WX709, I1995)
--	I1997 = NAND(I1987, I1995)
--	I1986 = NAND(I1996, I1997)
--	I2003 = NAND(WX773, WX837)
--	I2004 = NAND(WX773, I2003)
--	I2005 = NAND(WX837, I2003)
--	I2002 = NAND(I2004, I2005)
--	I2010 = NAND(I1986, I2002)
--	I2011 = NAND(I1986, I2010)
--	I2012 = NAND(I2002, I2010)
--	WX900 = NAND(I2011, I2012)
--	I2019 = NAND(WX1001, WX647)
--	I2020 = NAND(WX1001, I2019)
--	I2021 = NAND(WX647, I2019)
--	I2018 = NAND(I2020, I2021)
--	I2026 = NAND(WX711, I2018)
--	I2027 = NAND(WX711, I2026)
--	I2028 = NAND(I2018, I2026)
--	I2017 = NAND(I2027, I2028)
--	I2034 = NAND(WX775, WX839)
--	I2035 = NAND(WX775, I2034)
--	I2036 = NAND(WX839, I2034)
--	I2033 = NAND(I2035, I2036)
--	I2041 = NAND(I2017, I2033)
--	I2042 = NAND(I2017, I2041)
--	I2043 = NAND(I2033, I2041)
--	WX901 = NAND(I2042, I2043)
--	I2050 = NAND(WX1001, WX649)
--	I2051 = NAND(WX1001, I2050)
--	I2052 = NAND(WX649, I2050)
--	I2049 = NAND(I2051, I2052)
--	I2057 = NAND(WX713, I2049)
--	I2058 = NAND(WX713, I2057)
--	I2059 = NAND(I2049, I2057)
--	I2048 = NAND(I2058, I2059)
--	I2065 = NAND(WX777, WX841)
--	I2066 = NAND(WX777, I2065)
--	I2067 = NAND(WX841, I2065)
--	I2064 = NAND(I2066, I2067)
--	I2072 = NAND(I2048, I2064)
--	I2073 = NAND(I2048, I2072)
--	I2074 = NAND(I2064, I2072)
--	WX902 = NAND(I2073, I2074)
--	I2081 = NAND(WX1001, WX651)
--	I2082 = NAND(WX1001, I2081)
--	I2083 = NAND(WX651, I2081)
--	I2080 = NAND(I2082, I2083)
--	I2088 = NAND(WX715, I2080)
--	I2089 = NAND(WX715, I2088)
--	I2090 = NAND(I2080, I2088)
--	I2079 = NAND(I2089, I2090)
--	I2096 = NAND(WX779, WX843)
--	I2097 = NAND(WX779, I2096)
--	I2098 = NAND(WX843, I2096)
--	I2095 = NAND(I2097, I2098)
--	I2103 = NAND(I2079, I2095)
--	I2104 = NAND(I2079, I2103)
--	I2105 = NAND(I2095, I2103)
--	WX903 = NAND(I2104, I2105)
--	I2112 = NAND(WX1001, WX653)
--	I2113 = NAND(WX1001, I2112)
--	I2114 = NAND(WX653, I2112)
--	I2111 = NAND(I2113, I2114)
--	I2119 = NAND(WX717, I2111)
--	I2120 = NAND(WX717, I2119)
--	I2121 = NAND(I2111, I2119)
--	I2110 = NAND(I2120, I2121)
--	I2127 = NAND(WX781, WX845)
--	I2128 = NAND(WX781, I2127)
--	I2129 = NAND(WX845, I2127)
--	I2126 = NAND(I2128, I2129)
--	I2134 = NAND(I2110, I2126)
--	I2135 = NAND(I2110, I2134)
--	I2136 = NAND(I2126, I2134)
--	WX904 = NAND(I2135, I2136)
--	I2143 = NAND(WX1001, WX655)
--	I2144 = NAND(WX1001, I2143)
--	I2145 = NAND(WX655, I2143)
--	I2142 = NAND(I2144, I2145)
--	I2150 = NAND(WX719, I2142)
--	I2151 = NAND(WX719, I2150)
--	I2152 = NAND(I2142, I2150)
--	I2141 = NAND(I2151, I2152)
--	I2158 = NAND(WX783, WX847)
--	I2159 = NAND(WX783, I2158)
--	I2160 = NAND(WX847, I2158)
--	I2157 = NAND(I2159, I2160)
--	I2165 = NAND(I2141, I2157)
--	I2166 = NAND(I2141, I2165)
--	I2167 = NAND(I2157, I2165)
--	WX905 = NAND(I2166, I2167)
--	I2174 = NAND(WX1001, WX657)
--	I2175 = NAND(WX1001, I2174)
--	I2176 = NAND(WX657, I2174)
--	I2173 = NAND(I2175, I2176)
--	I2181 = NAND(WX721, I2173)
--	I2182 = NAND(WX721, I2181)
--	I2183 = NAND(I2173, I2181)
--	I2172 = NAND(I2182, I2183)
--	I2189 = NAND(WX785, WX849)
--	I2190 = NAND(WX785, I2189)
--	I2191 = NAND(WX849, I2189)
--	I2188 = NAND(I2190, I2191)
--	I2196 = NAND(I2172, I2188)
--	I2197 = NAND(I2172, I2196)
--	I2198 = NAND(I2188, I2196)
--	WX906 = NAND(I2197, I2198)
--	I2205 = NAND(WX1001, WX659)
--	I2206 = NAND(WX1001, I2205)
--	I2207 = NAND(WX659, I2205)
--	I2204 = NAND(I2206, I2207)
--	I2212 = NAND(WX723, I2204)
--	I2213 = NAND(WX723, I2212)
--	I2214 = NAND(I2204, I2212)
--	I2203 = NAND(I2213, I2214)
--	I2220 = NAND(WX787, WX851)
--	I2221 = NAND(WX787, I2220)
--	I2222 = NAND(WX851, I2220)
--	I2219 = NAND(I2221, I2222)
--	I2227 = NAND(I2203, I2219)
--	I2228 = NAND(I2203, I2227)
--	I2229 = NAND(I2219, I2227)
--	WX907 = NAND(I2228, I2229)
--	I2236 = NAND(WX1001, WX661)
--	I2237 = NAND(WX1001, I2236)
--	I2238 = NAND(WX661, I2236)
--	I2235 = NAND(I2237, I2238)
--	I2243 = NAND(WX725, I2235)
--	I2244 = NAND(WX725, I2243)
--	I2245 = NAND(I2235, I2243)
--	I2234 = NAND(I2244, I2245)
--	I2251 = NAND(WX789, WX853)
--	I2252 = NAND(WX789, I2251)
--	I2253 = NAND(WX853, I2251)
--	I2250 = NAND(I2252, I2253)
--	I2258 = NAND(I2234, I2250)
--	I2259 = NAND(I2234, I2258)
--	I2260 = NAND(I2250, I2258)
--	WX908 = NAND(I2259, I2260)
--	I2267 = NAND(WX1001, WX663)
--	I2268 = NAND(WX1001, I2267)
--	I2269 = NAND(WX663, I2267)
--	I2266 = NAND(I2268, I2269)
--	I2274 = NAND(WX727, I2266)
--	I2275 = NAND(WX727, I2274)
--	I2276 = NAND(I2266, I2274)
--	I2265 = NAND(I2275, I2276)
--	I2282 = NAND(WX791, WX855)
--	I2283 = NAND(WX791, I2282)
--	I2284 = NAND(WX855, I2282)
--	I2281 = NAND(I2283, I2284)
--	I2289 = NAND(I2265, I2281)
--	I2290 = NAND(I2265, I2289)
--	I2291 = NAND(I2281, I2289)
--	WX909 = NAND(I2290, I2291)
--	I2298 = NAND(WX1001, WX665)
--	I2299 = NAND(WX1001, I2298)
--	I2300 = NAND(WX665, I2298)
--	I2297 = NAND(I2299, I2300)
--	I2305 = NAND(WX729, I2297)
--	I2306 = NAND(WX729, I2305)
--	I2307 = NAND(I2297, I2305)
--	I2296 = NAND(I2306, I2307)
--	I2313 = NAND(WX793, WX857)
--	I2314 = NAND(WX793, I2313)
--	I2315 = NAND(WX857, I2313)
--	I2312 = NAND(I2314, I2315)
--	I2320 = NAND(I2296, I2312)
--	I2321 = NAND(I2296, I2320)
--	I2322 = NAND(I2312, I2320)
--	WX910 = NAND(I2321, I2322)
--	I2329 = NAND(WX1001, WX667)
--	I2330 = NAND(WX1001, I2329)
--	I2331 = NAND(WX667, I2329)
--	I2328 = NAND(I2330, I2331)
--	I2336 = NAND(WX731, I2328)
--	I2337 = NAND(WX731, I2336)
--	I2338 = NAND(I2328, I2336)
--	I2327 = NAND(I2337, I2338)
--	I2344 = NAND(WX795, WX859)
--	I2345 = NAND(WX795, I2344)
--	I2346 = NAND(WX859, I2344)
--	I2343 = NAND(I2345, I2346)
--	I2351 = NAND(I2327, I2343)
--	I2352 = NAND(I2327, I2351)
--	I2353 = NAND(I2343, I2351)
--	WX911 = NAND(I2352, I2353)
--	I2360 = NAND(WX1001, WX669)
--	I2361 = NAND(WX1001, I2360)
--	I2362 = NAND(WX669, I2360)
--	I2359 = NAND(I2361, I2362)
--	I2367 = NAND(WX733, I2359)
--	I2368 = NAND(WX733, I2367)
--	I2369 = NAND(I2359, I2367)
--	I2358 = NAND(I2368, I2369)
--	I2375 = NAND(WX797, WX861)
--	I2376 = NAND(WX797, I2375)
--	I2377 = NAND(WX861, I2375)
--	I2374 = NAND(I2376, I2377)
--	I2382 = NAND(I2358, I2374)
--	I2383 = NAND(I2358, I2382)
--	I2384 = NAND(I2374, I2382)
--	WX912 = NAND(I2383, I2384)
--	I2391 = NAND(WX1001, WX671)
--	I2392 = NAND(WX1001, I2391)
--	I2393 = NAND(WX671, I2391)
--	I2390 = NAND(I2392, I2393)
--	I2398 = NAND(WX735, I2390)
--	I2399 = NAND(WX735, I2398)
--	I2400 = NAND(I2390, I2398)
--	I2389 = NAND(I2399, I2400)
--	I2406 = NAND(WX799, WX863)
--	I2407 = NAND(WX799, I2406)
--	I2408 = NAND(WX863, I2406)
--	I2405 = NAND(I2407, I2408)
--	I2413 = NAND(I2389, I2405)
--	I2414 = NAND(I2389, I2413)
--	I2415 = NAND(I2405, I2413)
--	WX913 = NAND(I2414, I2415)
--	I2422 = NAND(WX1001, WX673)
--	I2423 = NAND(WX1001, I2422)
--	I2424 = NAND(WX673, I2422)
--	I2421 = NAND(I2423, I2424)
--	I2429 = NAND(WX737, I2421)
--	I2430 = NAND(WX737, I2429)
--	I2431 = NAND(I2421, I2429)
--	I2420 = NAND(I2430, I2431)
--	I2437 = NAND(WX801, WX865)
--	I2438 = NAND(WX801, I2437)
--	I2439 = NAND(WX865, I2437)
--	I2436 = NAND(I2438, I2439)
--	I2444 = NAND(I2420, I2436)
--	I2445 = NAND(I2420, I2444)
--	I2446 = NAND(I2436, I2444)
--	WX914 = NAND(I2445, I2446)
--	I2453 = NAND(WX1001, WX675)
--	I2454 = NAND(WX1001, I2453)
--	I2455 = NAND(WX675, I2453)
--	I2452 = NAND(I2454, I2455)
--	I2460 = NAND(WX739, I2452)
--	I2461 = NAND(WX739, I2460)
--	I2462 = NAND(I2452, I2460)
--	I2451 = NAND(I2461, I2462)
--	I2468 = NAND(WX803, WX867)
--	I2469 = NAND(WX803, I2468)
--	I2470 = NAND(WX867, I2468)
--	I2467 = NAND(I2469, I2470)
--	I2475 = NAND(I2451, I2467)
--	I2476 = NAND(I2451, I2475)
--	I2477 = NAND(I2467, I2475)
--	WX915 = NAND(I2476, I2477)
--	I2484 = NAND(WX1002, WX677)
--	I2485 = NAND(WX1002, I2484)
--	I2486 = NAND(WX677, I2484)
--	I2483 = NAND(I2485, I2486)
--	I2491 = NAND(WX741, I2483)
--	I2492 = NAND(WX741, I2491)
--	I2493 = NAND(I2483, I2491)
--	I2482 = NAND(I2492, I2493)
--	I2499 = NAND(WX805, WX869)
--	I2500 = NAND(WX805, I2499)
--	I2501 = NAND(WX869, I2499)
--	I2498 = NAND(I2500, I2501)
--	I2506 = NAND(I2482, I2498)
--	I2507 = NAND(I2482, I2506)
--	I2508 = NAND(I2498, I2506)
--	WX916 = NAND(I2507, I2508)
--	I2515 = NAND(WX1002, WX679)
--	I2516 = NAND(WX1002, I2515)
--	I2517 = NAND(WX679, I2515)
--	I2514 = NAND(I2516, I2517)
--	I2522 = NAND(WX743, I2514)
--	I2523 = NAND(WX743, I2522)
--	I2524 = NAND(I2514, I2522)
--	I2513 = NAND(I2523, I2524)
--	I2530 = NAND(WX807, WX871)
--	I2531 = NAND(WX807, I2530)
--	I2532 = NAND(WX871, I2530)
--	I2529 = NAND(I2531, I2532)
--	I2537 = NAND(I2513, I2529)
--	I2538 = NAND(I2513, I2537)
--	I2539 = NAND(I2529, I2537)
--	WX917 = NAND(I2538, I2539)
--	I2546 = NAND(WX1002, WX681)
--	I2547 = NAND(WX1002, I2546)
--	I2548 = NAND(WX681, I2546)
--	I2545 = NAND(I2547, I2548)
--	I2553 = NAND(WX745, I2545)
--	I2554 = NAND(WX745, I2553)
--	I2555 = NAND(I2545, I2553)
--	I2544 = NAND(I2554, I2555)
--	I2561 = NAND(WX809, WX873)
--	I2562 = NAND(WX809, I2561)
--	I2563 = NAND(WX873, I2561)
--	I2560 = NAND(I2562, I2563)
--	I2568 = NAND(I2544, I2560)
--	I2569 = NAND(I2544, I2568)
--	I2570 = NAND(I2560, I2568)
--	WX918 = NAND(I2569, I2570)
--	I2577 = NAND(WX1002, WX683)
--	I2578 = NAND(WX1002, I2577)
--	I2579 = NAND(WX683, I2577)
--	I2576 = NAND(I2578, I2579)
--	I2584 = NAND(WX747, I2576)
--	I2585 = NAND(WX747, I2584)
--	I2586 = NAND(I2576, I2584)
--	I2575 = NAND(I2585, I2586)
--	I2592 = NAND(WX811, WX875)
--	I2593 = NAND(WX811, I2592)
--	I2594 = NAND(WX875, I2592)
--	I2591 = NAND(I2593, I2594)
--	I2599 = NAND(I2575, I2591)
--	I2600 = NAND(I2575, I2599)
--	I2601 = NAND(I2591, I2599)
--	WX919 = NAND(I2600, I2601)
--	I2608 = NAND(WX1002, WX685)
--	I2609 = NAND(WX1002, I2608)
--	I2610 = NAND(WX685, I2608)
--	I2607 = NAND(I2609, I2610)
--	I2615 = NAND(WX749, I2607)
--	I2616 = NAND(WX749, I2615)
--	I2617 = NAND(I2607, I2615)
--	I2606 = NAND(I2616, I2617)
--	I2623 = NAND(WX813, WX877)
--	I2624 = NAND(WX813, I2623)
--	I2625 = NAND(WX877, I2623)
--	I2622 = NAND(I2624, I2625)
--	I2630 = NAND(I2606, I2622)
--	I2631 = NAND(I2606, I2630)
--	I2632 = NAND(I2622, I2630)
--	WX920 = NAND(I2631, I2632)
--	I2639 = NAND(WX1002, WX687)
--	I2640 = NAND(WX1002, I2639)
--	I2641 = NAND(WX687, I2639)
--	I2638 = NAND(I2640, I2641)
--	I2646 = NAND(WX751, I2638)
--	I2647 = NAND(WX751, I2646)
--	I2648 = NAND(I2638, I2646)
--	I2637 = NAND(I2647, I2648)
--	I2654 = NAND(WX815, WX879)
--	I2655 = NAND(WX815, I2654)
--	I2656 = NAND(WX879, I2654)
--	I2653 = NAND(I2655, I2656)
--	I2661 = NAND(I2637, I2653)
--	I2662 = NAND(I2637, I2661)
--	I2663 = NAND(I2653, I2661)
--	WX921 = NAND(I2662, I2663)
--	I2670 = NAND(WX1002, WX689)
--	I2671 = NAND(WX1002, I2670)
--	I2672 = NAND(WX689, I2670)
--	I2669 = NAND(I2671, I2672)
--	I2677 = NAND(WX753, I2669)
--	I2678 = NAND(WX753, I2677)
--	I2679 = NAND(I2669, I2677)
--	I2668 = NAND(I2678, I2679)
--	I2685 = NAND(WX817, WX881)
--	I2686 = NAND(WX817, I2685)
--	I2687 = NAND(WX881, I2685)
--	I2684 = NAND(I2686, I2687)
--	I2692 = NAND(I2668, I2684)
--	I2693 = NAND(I2668, I2692)
--	I2694 = NAND(I2684, I2692)
--	WX922 = NAND(I2693, I2694)
--	I2701 = NAND(WX1002, WX691)
--	I2702 = NAND(WX1002, I2701)
--	I2703 = NAND(WX691, I2701)
--	I2700 = NAND(I2702, I2703)
--	I2708 = NAND(WX755, I2700)
--	I2709 = NAND(WX755, I2708)
--	I2710 = NAND(I2700, I2708)
--	I2699 = NAND(I2709, I2710)
--	I2716 = NAND(WX819, WX883)
--	I2717 = NAND(WX819, I2716)
--	I2718 = NAND(WX883, I2716)
--	I2715 = NAND(I2717, I2718)
--	I2723 = NAND(I2699, I2715)
--	I2724 = NAND(I2699, I2723)
--	I2725 = NAND(I2715, I2723)
--	WX923 = NAND(I2724, I2725)
--	I2732 = NAND(WX1002, WX693)
--	I2733 = NAND(WX1002, I2732)
--	I2734 = NAND(WX693, I2732)
--	I2731 = NAND(I2733, I2734)
--	I2739 = NAND(WX757, I2731)
--	I2740 = NAND(WX757, I2739)
--	I2741 = NAND(I2731, I2739)
--	I2730 = NAND(I2740, I2741)
--	I2747 = NAND(WX821, WX885)
--	I2748 = NAND(WX821, I2747)
--	I2749 = NAND(WX885, I2747)
--	I2746 = NAND(I2748, I2749)
--	I2754 = NAND(I2730, I2746)
--	I2755 = NAND(I2730, I2754)
--	I2756 = NAND(I2746, I2754)
--	WX924 = NAND(I2755, I2756)
--	I2763 = NAND(WX1002, WX695)
--	I2764 = NAND(WX1002, I2763)
--	I2765 = NAND(WX695, I2763)
--	I2762 = NAND(I2764, I2765)
--	I2770 = NAND(WX759, I2762)
--	I2771 = NAND(WX759, I2770)
--	I2772 = NAND(I2762, I2770)
--	I2761 = NAND(I2771, I2772)
--	I2778 = NAND(WX823, WX887)
--	I2779 = NAND(WX823, I2778)
--	I2780 = NAND(WX887, I2778)
--	I2777 = NAND(I2779, I2780)
--	I2785 = NAND(I2761, I2777)
--	I2786 = NAND(I2761, I2785)
--	I2787 = NAND(I2777, I2785)
--	WX925 = NAND(I2786, I2787)
--	I2794 = NAND(WX1002, WX697)
--	I2795 = NAND(WX1002, I2794)
--	I2796 = NAND(WX697, I2794)
--	I2793 = NAND(I2795, I2796)
--	I2801 = NAND(WX761, I2793)
--	I2802 = NAND(WX761, I2801)
--	I2803 = NAND(I2793, I2801)
--	I2792 = NAND(I2802, I2803)
--	I2809 = NAND(WX825, WX889)
--	I2810 = NAND(WX825, I2809)
--	I2811 = NAND(WX889, I2809)
--	I2808 = NAND(I2810, I2811)
--	I2816 = NAND(I2792, I2808)
--	I2817 = NAND(I2792, I2816)
--	I2818 = NAND(I2808, I2816)
--	WX926 = NAND(I2817, I2818)
--	I2825 = NAND(WX1002, WX699)
--	I2826 = NAND(WX1002, I2825)
--	I2827 = NAND(WX699, I2825)
--	I2824 = NAND(I2826, I2827)
--	I2832 = NAND(WX763, I2824)
--	I2833 = NAND(WX763, I2832)
--	I2834 = NAND(I2824, I2832)
--	I2823 = NAND(I2833, I2834)
--	I2840 = NAND(WX827, WX891)
--	I2841 = NAND(WX827, I2840)
--	I2842 = NAND(WX891, I2840)
--	I2839 = NAND(I2841, I2842)
--	I2847 = NAND(I2823, I2839)
--	I2848 = NAND(I2823, I2847)
--	I2849 = NAND(I2839, I2847)
--	WX927 = NAND(I2848, I2849)
--	I2856 = NAND(WX1002, WX701)
--	I2857 = NAND(WX1002, I2856)
--	I2858 = NAND(WX701, I2856)
--	I2855 = NAND(I2857, I2858)
--	I2863 = NAND(WX765, I2855)
--	I2864 = NAND(WX765, I2863)
--	I2865 = NAND(I2855, I2863)
--	I2854 = NAND(I2864, I2865)
--	I2871 = NAND(WX829, WX893)
--	I2872 = NAND(WX829, I2871)
--	I2873 = NAND(WX893, I2871)
--	I2870 = NAND(I2872, I2873)
--	I2878 = NAND(I2854, I2870)
--	I2879 = NAND(I2854, I2878)
--	I2880 = NAND(I2870, I2878)
--	WX928 = NAND(I2879, I2880)
--	I2887 = NAND(WX1002, WX703)
--	I2888 = NAND(WX1002, I2887)
--	I2889 = NAND(WX703, I2887)
--	I2886 = NAND(I2888, I2889)
--	I2894 = NAND(WX767, I2886)
--	I2895 = NAND(WX767, I2894)
--	I2896 = NAND(I2886, I2894)
--	I2885 = NAND(I2895, I2896)
--	I2902 = NAND(WX831, WX895)
--	I2903 = NAND(WX831, I2902)
--	I2904 = NAND(WX895, I2902)
--	I2901 = NAND(I2903, I2904)
--	I2909 = NAND(I2885, I2901)
--	I2910 = NAND(I2885, I2909)
--	I2911 = NAND(I2901, I2909)
--	WX929 = NAND(I2910, I2911)
--	I2918 = NAND(WX1002, WX705)
--	I2919 = NAND(WX1002, I2918)
--	I2920 = NAND(WX705, I2918)
--	I2917 = NAND(I2919, I2920)
--	I2925 = NAND(WX769, I2917)
--	I2926 = NAND(WX769, I2925)
--	I2927 = NAND(I2917, I2925)
--	I2916 = NAND(I2926, I2927)
--	I2933 = NAND(WX833, WX897)
--	I2934 = NAND(WX833, I2933)
--	I2935 = NAND(WX897, I2933)
--	I2932 = NAND(I2934, I2935)
--	I2940 = NAND(I2916, I2932)
--	I2941 = NAND(I2916, I2940)
--	I2942 = NAND(I2932, I2940)
--	WX930 = NAND(I2941, I2942)
--	I2949 = NAND(WX1002, WX707)
--	I2950 = NAND(WX1002, I2949)
--	I2951 = NAND(WX707, I2949)
--	I2948 = NAND(I2950, I2951)
--	I2956 = NAND(WX771, I2948)
--	I2957 = NAND(WX771, I2956)
--	I2958 = NAND(I2948, I2956)
--	I2947 = NAND(I2957, I2958)
--	I2964 = NAND(WX835, WX899)
--	I2965 = NAND(WX835, I2964)
--	I2966 = NAND(WX899, I2964)
--	I2963 = NAND(I2965, I2966)
--	I2971 = NAND(I2947, I2963)
--	I2972 = NAND(I2947, I2971)
--	I2973 = NAND(I2963, I2971)
--	WX931 = NAND(I2972, I2973)
--	I3052 = NAND(WX580, WX485)
--	I3053 = NAND(WX580, I3052)
--	I3054 = NAND(WX485, I3052)
--	WX1006 = NAND(I3053, I3054)
--	I3065 = NAND(WX581, WX487)
--	I3066 = NAND(WX581, I3065)
--	I3067 = NAND(WX487, I3065)
--	WX1013 = NAND(I3066, I3067)
--	I3078 = NAND(WX582, WX489)
--	I3079 = NAND(WX582, I3078)
--	I3080 = NAND(WX489, I3078)
--	WX1020 = NAND(I3079, I3080)
--	I3091 = NAND(WX583, WX491)
--	I3092 = NAND(WX583, I3091)
--	I3093 = NAND(WX491, I3091)
--	WX1027 = NAND(I3092, I3093)
--	I3104 = NAND(WX584, WX493)
--	I3105 = NAND(WX584, I3104)
--	I3106 = NAND(WX493, I3104)
--	WX1034 = NAND(I3105, I3106)
--	I3117 = NAND(WX585, WX495)
--	I3118 = NAND(WX585, I3117)
--	I3119 = NAND(WX495, I3117)
--	WX1041 = NAND(I3118, I3119)
--	I3130 = NAND(WX586, WX497)
--	I3131 = NAND(WX586, I3130)
--	I3132 = NAND(WX497, I3130)
--	WX1048 = NAND(I3131, I3132)
--	I3143 = NAND(WX587, WX499)
--	I3144 = NAND(WX587, I3143)
--	I3145 = NAND(WX499, I3143)
--	WX1055 = NAND(I3144, I3145)
--	I3156 = NAND(WX588, WX501)
--	I3157 = NAND(WX588, I3156)
--	I3158 = NAND(WX501, I3156)
--	WX1062 = NAND(I3157, I3158)
--	I3169 = NAND(WX589, WX503)
--	I3170 = NAND(WX589, I3169)
--	I3171 = NAND(WX503, I3169)
--	WX1069 = NAND(I3170, I3171)
--	I3182 = NAND(WX590, WX505)
--	I3183 = NAND(WX590, I3182)
--	I3184 = NAND(WX505, I3182)
--	WX1076 = NAND(I3183, I3184)
--	I3195 = NAND(WX591, WX507)
--	I3196 = NAND(WX591, I3195)
--	I3197 = NAND(WX507, I3195)
--	WX1083 = NAND(I3196, I3197)
--	I3208 = NAND(WX592, WX509)
--	I3209 = NAND(WX592, I3208)
--	I3210 = NAND(WX509, I3208)
--	WX1090 = NAND(I3209, I3210)
--	I3221 = NAND(WX593, WX511)
--	I3222 = NAND(WX593, I3221)
--	I3223 = NAND(WX511, I3221)
--	WX1097 = NAND(I3222, I3223)
--	I3234 = NAND(WX594, WX513)
--	I3235 = NAND(WX594, I3234)
--	I3236 = NAND(WX513, I3234)
--	WX1104 = NAND(I3235, I3236)
--	I3247 = NAND(WX595, WX515)
--	I3248 = NAND(WX595, I3247)
--	I3249 = NAND(WX515, I3247)
--	WX1111 = NAND(I3248, I3249)
--	I3260 = NAND(WX596, WX517)
--	I3261 = NAND(WX596, I3260)
--	I3262 = NAND(WX517, I3260)
--	WX1118 = NAND(I3261, I3262)
--	I3273 = NAND(WX597, WX519)
--	I3274 = NAND(WX597, I3273)
--	I3275 = NAND(WX519, I3273)
--	WX1125 = NAND(I3274, I3275)
--	I3286 = NAND(WX598, WX521)
--	I3287 = NAND(WX598, I3286)
--	I3288 = NAND(WX521, I3286)
--	WX1132 = NAND(I3287, I3288)
--	I3299 = NAND(WX599, WX523)
--	I3300 = NAND(WX599, I3299)
--	I3301 = NAND(WX523, I3299)
--	WX1139 = NAND(I3300, I3301)
--	I3312 = NAND(WX600, WX525)
--	I3313 = NAND(WX600, I3312)
--	I3314 = NAND(WX525, I3312)
--	WX1146 = NAND(I3313, I3314)
--	I3325 = NAND(WX601, WX527)
--	I3326 = NAND(WX601, I3325)
--	I3327 = NAND(WX527, I3325)
--	WX1153 = NAND(I3326, I3327)
--	I3338 = NAND(WX602, WX529)
--	I3339 = NAND(WX602, I3338)
--	I3340 = NAND(WX529, I3338)
--	WX1160 = NAND(I3339, I3340)
--	I3351 = NAND(WX603, WX531)
--	I3352 = NAND(WX603, I3351)
--	I3353 = NAND(WX531, I3351)
--	WX1167 = NAND(I3352, I3353)
--	I3364 = NAND(WX604, WX533)
--	I3365 = NAND(WX604, I3364)
--	I3366 = NAND(WX533, I3364)
--	WX1174 = NAND(I3365, I3366)
--	I3377 = NAND(WX605, WX535)
--	I3378 = NAND(WX605, I3377)
--	I3379 = NAND(WX535, I3377)
--	WX1181 = NAND(I3378, I3379)
--	I3390 = NAND(WX606, WX537)
--	I3391 = NAND(WX606, I3390)
--	I3392 = NAND(WX537, I3390)
--	WX1188 = NAND(I3391, I3392)
--	I3403 = NAND(WX607, WX539)
--	I3404 = NAND(WX607, I3403)
--	I3405 = NAND(WX539, I3403)
--	WX1195 = NAND(I3404, I3405)
--	I3416 = NAND(WX608, WX541)
--	I3417 = NAND(WX608, I3416)
--	I3418 = NAND(WX541, I3416)
--	WX1202 = NAND(I3417, I3418)
--	I3429 = NAND(WX609, WX543)
--	I3430 = NAND(WX609, I3429)
--	I3431 = NAND(WX543, I3429)
--	WX1209 = NAND(I3430, I3431)
--	I3442 = NAND(WX610, WX545)
--	I3443 = NAND(WX610, I3442)
--	I3444 = NAND(WX545, I3442)
--	WX1216 = NAND(I3443, I3444)
--	I3455 = NAND(WX611, WX547)
--	I3456 = NAND(WX611, I3455)
--	I3457 = NAND(WX547, I3455)
--	WX1223 = NAND(I3456, I3457)
--	I3470 = NAND(WX627, CRC_OUT_9_31)
--	I3471 = NAND(WX627, I3470)
--	I3472 = NAND(CRC_OUT_9_31, I3470)
--	I3469 = NAND(I3471, I3472)
--	I3477 = NAND(CRC_OUT_9_15, I3469)
--	I3478 = NAND(CRC_OUT_9_15, I3477)
--	I3479 = NAND(I3469, I3477)
--	WX1231 = NAND(I3478, I3479)
--	I3485 = NAND(WX632, CRC_OUT_9_31)
--	I3486 = NAND(WX632, I3485)
--	I3487 = NAND(CRC_OUT_9_31, I3485)
--	I3484 = NAND(I3486, I3487)
--	I3492 = NAND(CRC_OUT_9_10, I3484)
--	I3493 = NAND(CRC_OUT_9_10, I3492)
--	I3494 = NAND(I3484, I3492)
--	WX1232 = NAND(I3493, I3494)
--	I3500 = NAND(WX639, CRC_OUT_9_31)
--	I3501 = NAND(WX639, I3500)
--	I3502 = NAND(CRC_OUT_9_31, I3500)
--	I3499 = NAND(I3501, I3502)
--	I3507 = NAND(CRC_OUT_9_3, I3499)
--	I3508 = NAND(CRC_OUT_9_3, I3507)
--	I3509 = NAND(I3499, I3507)
--	WX1233 = NAND(I3508, I3509)
--	I3514 = NAND(WX643, CRC_OUT_9_31)
--	I3515 = NAND(WX643, I3514)
--	I3516 = NAND(CRC_OUT_9_31, I3514)
--	WX1234 = NAND(I3515, I3516)
--	I3521 = NAND(WX612, CRC_OUT_9_30)
--	I3522 = NAND(WX612, I3521)
--	I3523 = NAND(CRC_OUT_9_30, I3521)
--	WX1235 = NAND(I3522, I3523)
--	I3528 = NAND(WX613, CRC_OUT_9_29)
--	I3529 = NAND(WX613, I3528)
--	I3530 = NAND(CRC_OUT_9_29, I3528)
--	WX1236 = NAND(I3529, I3530)
--	I3535 = NAND(WX614, CRC_OUT_9_28)
--	I3536 = NAND(WX614, I3535)
--	I3537 = NAND(CRC_OUT_9_28, I3535)
--	WX1237 = NAND(I3536, I3537)
--	I3542 = NAND(WX615, CRC_OUT_9_27)
--	I3543 = NAND(WX615, I3542)
--	I3544 = NAND(CRC_OUT_9_27, I3542)
--	WX1238 = NAND(I3543, I3544)
--	I3549 = NAND(WX616, CRC_OUT_9_26)
--	I3550 = NAND(WX616, I3549)
--	I3551 = NAND(CRC_OUT_9_26, I3549)
--	WX1239 = NAND(I3550, I3551)
--	I3556 = NAND(WX617, CRC_OUT_9_25)
--	I3557 = NAND(WX617, I3556)
--	I3558 = NAND(CRC_OUT_9_25, I3556)
--	WX1240 = NAND(I3557, I3558)
--	I3563 = NAND(WX618, CRC_OUT_9_24)
--	I3564 = NAND(WX618, I3563)
--	I3565 = NAND(CRC_OUT_9_24, I3563)
--	WX1241 = NAND(I3564, I3565)
--	I3570 = NAND(WX619, CRC_OUT_9_23)
--	I3571 = NAND(WX619, I3570)
--	I3572 = NAND(CRC_OUT_9_23, I3570)
--	WX1242 = NAND(I3571, I3572)
--	I3577 = NAND(WX620, CRC_OUT_9_22)
--	I3578 = NAND(WX620, I3577)
--	I3579 = NAND(CRC_OUT_9_22, I3577)
--	WX1243 = NAND(I3578, I3579)
--	I3584 = NAND(WX621, CRC_OUT_9_21)
--	I3585 = NAND(WX621, I3584)
--	I3586 = NAND(CRC_OUT_9_21, I3584)
--	WX1244 = NAND(I3585, I3586)
--	I3591 = NAND(WX622, CRC_OUT_9_20)
--	I3592 = NAND(WX622, I3591)
--	I3593 = NAND(CRC_OUT_9_20, I3591)
--	WX1245 = NAND(I3592, I3593)
--	I3598 = NAND(WX623, CRC_OUT_9_19)
--	I3599 = NAND(WX623, I3598)
--	I3600 = NAND(CRC_OUT_9_19, I3598)
--	WX1246 = NAND(I3599, I3600)
--	I3605 = NAND(WX624, CRC_OUT_9_18)
--	I3606 = NAND(WX624, I3605)
--	I3607 = NAND(CRC_OUT_9_18, I3605)
--	WX1247 = NAND(I3606, I3607)
--	I3612 = NAND(WX625, CRC_OUT_9_17)
--	I3613 = NAND(WX625, I3612)
--	I3614 = NAND(CRC_OUT_9_17, I3612)
--	WX1248 = NAND(I3613, I3614)
--	I3619 = NAND(WX626, CRC_OUT_9_16)
--	I3620 = NAND(WX626, I3619)
--	I3621 = NAND(CRC_OUT_9_16, I3619)
--	WX1249 = NAND(I3620, I3621)
--	I3626 = NAND(WX628, CRC_OUT_9_14)
--	I3627 = NAND(WX628, I3626)
--	I3628 = NAND(CRC_OUT_9_14, I3626)
--	WX1250 = NAND(I3627, I3628)
--	I3633 = NAND(WX629, CRC_OUT_9_13)
--	I3634 = NAND(WX629, I3633)
--	I3635 = NAND(CRC_OUT_9_13, I3633)
--	WX1251 = NAND(I3634, I3635)
--	I3640 = NAND(WX630, CRC_OUT_9_12)
--	I3641 = NAND(WX630, I3640)
--	I3642 = NAND(CRC_OUT_9_12, I3640)
--	WX1252 = NAND(I3641, I3642)
--	I3647 = NAND(WX631, CRC_OUT_9_11)
--	I3648 = NAND(WX631, I3647)
--	I3649 = NAND(CRC_OUT_9_11, I3647)
--	WX1253 = NAND(I3648, I3649)
--	I3654 = NAND(WX633, CRC_OUT_9_9)
--	I3655 = NAND(WX633, I3654)
--	I3656 = NAND(CRC_OUT_9_9, I3654)
--	WX1254 = NAND(I3655, I3656)
--	I3661 = NAND(WX634, CRC_OUT_9_8)
--	I3662 = NAND(WX634, I3661)
--	I3663 = NAND(CRC_OUT_9_8, I3661)
--	WX1255 = NAND(I3662, I3663)
--	I3668 = NAND(WX635, CRC_OUT_9_7)
--	I3669 = NAND(WX635, I3668)
--	I3670 = NAND(CRC_OUT_9_7, I3668)
--	WX1256 = NAND(I3669, I3670)
--	I3675 = NAND(WX636, CRC_OUT_9_6)
--	I3676 = NAND(WX636, I3675)
--	I3677 = NAND(CRC_OUT_9_6, I3675)
--	WX1257 = NAND(I3676, I3677)
--	I3682 = NAND(WX637, CRC_OUT_9_5)
--	I3683 = NAND(WX637, I3682)
--	I3684 = NAND(CRC_OUT_9_5, I3682)
--	WX1258 = NAND(I3683, I3684)
--	I3689 = NAND(WX638, CRC_OUT_9_4)
--	I3690 = NAND(WX638, I3689)
--	I3691 = NAND(CRC_OUT_9_4, I3689)
--	WX1259 = NAND(I3690, I3691)
--	I3696 = NAND(WX640, CRC_OUT_9_2)
--	I3697 = NAND(WX640, I3696)
--	I3698 = NAND(CRC_OUT_9_2, I3696)
--	WX1260 = NAND(I3697, I3698)
--	I3703 = NAND(WX641, CRC_OUT_9_1)
--	I3704 = NAND(WX641, I3703)
--	I3705 = NAND(CRC_OUT_9_1, I3703)
--	WX1261 = NAND(I3704, I3705)
--	I3710 = NAND(WX642, CRC_OUT_9_0)
--	I3711 = NAND(WX642, I3710)
--	I3712 = NAND(CRC_OUT_9_0, I3710)
--	WX1262 = NAND(I3711, I3712)
--	I5993 = NAND(WX2294, WX1938)
--	I5994 = NAND(WX2294, I5993)
--	I5995 = NAND(WX1938, I5993)
--	I5992 = NAND(I5994, I5995)
--	I6000 = NAND(WX2002, I5992)
--	I6001 = NAND(WX2002, I6000)
--	I6002 = NAND(I5992, I6000)
--	I5991 = NAND(I6001, I6002)
--	I6008 = NAND(WX2066, WX2130)
--	I6009 = NAND(WX2066, I6008)
--	I6010 = NAND(WX2130, I6008)
--	I6007 = NAND(I6009, I6010)
--	I6015 = NAND(I5991, I6007)
--	I6016 = NAND(I5991, I6015)
--	I6017 = NAND(I6007, I6015)
--	WX2193 = NAND(I6016, I6017)
--	I6024 = NAND(WX2294, WX1940)
--	I6025 = NAND(WX2294, I6024)
--	I6026 = NAND(WX1940, I6024)
--	I6023 = NAND(I6025, I6026)
--	I6031 = NAND(WX2004, I6023)
--	I6032 = NAND(WX2004, I6031)
--	I6033 = NAND(I6023, I6031)
--	I6022 = NAND(I6032, I6033)
--	I6039 = NAND(WX2068, WX2132)
--	I6040 = NAND(WX2068, I6039)
--	I6041 = NAND(WX2132, I6039)
--	I6038 = NAND(I6040, I6041)
--	I6046 = NAND(I6022, I6038)
--	I6047 = NAND(I6022, I6046)
--	I6048 = NAND(I6038, I6046)
--	WX2194 = NAND(I6047, I6048)
--	I6055 = NAND(WX2294, WX1942)
--	I6056 = NAND(WX2294, I6055)
--	I6057 = NAND(WX1942, I6055)
--	I6054 = NAND(I6056, I6057)
--	I6062 = NAND(WX2006, I6054)
--	I6063 = NAND(WX2006, I6062)
--	I6064 = NAND(I6054, I6062)
--	I6053 = NAND(I6063, I6064)
--	I6070 = NAND(WX2070, WX2134)
--	I6071 = NAND(WX2070, I6070)
--	I6072 = NAND(WX2134, I6070)
--	I6069 = NAND(I6071, I6072)
--	I6077 = NAND(I6053, I6069)
--	I6078 = NAND(I6053, I6077)
--	I6079 = NAND(I6069, I6077)
--	WX2195 = NAND(I6078, I6079)
--	I6086 = NAND(WX2294, WX1944)
--	I6087 = NAND(WX2294, I6086)
--	I6088 = NAND(WX1944, I6086)
--	I6085 = NAND(I6087, I6088)
--	I6093 = NAND(WX2008, I6085)
--	I6094 = NAND(WX2008, I6093)
--	I6095 = NAND(I6085, I6093)
--	I6084 = NAND(I6094, I6095)
--	I6101 = NAND(WX2072, WX2136)
--	I6102 = NAND(WX2072, I6101)
--	I6103 = NAND(WX2136, I6101)
--	I6100 = NAND(I6102, I6103)
--	I6108 = NAND(I6084, I6100)
--	I6109 = NAND(I6084, I6108)
--	I6110 = NAND(I6100, I6108)
--	WX2196 = NAND(I6109, I6110)
--	I6117 = NAND(WX2294, WX1946)
--	I6118 = NAND(WX2294, I6117)
--	I6119 = NAND(WX1946, I6117)
--	I6116 = NAND(I6118, I6119)
--	I6124 = NAND(WX2010, I6116)
--	I6125 = NAND(WX2010, I6124)
--	I6126 = NAND(I6116, I6124)
--	I6115 = NAND(I6125, I6126)
--	I6132 = NAND(WX2074, WX2138)
--	I6133 = NAND(WX2074, I6132)
--	I6134 = NAND(WX2138, I6132)
--	I6131 = NAND(I6133, I6134)
--	I6139 = NAND(I6115, I6131)
--	I6140 = NAND(I6115, I6139)
--	I6141 = NAND(I6131, I6139)
--	WX2197 = NAND(I6140, I6141)
--	I6148 = NAND(WX2294, WX1948)
--	I6149 = NAND(WX2294, I6148)
--	I6150 = NAND(WX1948, I6148)
--	I6147 = NAND(I6149, I6150)
--	I6155 = NAND(WX2012, I6147)
--	I6156 = NAND(WX2012, I6155)
--	I6157 = NAND(I6147, I6155)
--	I6146 = NAND(I6156, I6157)
--	I6163 = NAND(WX2076, WX2140)
--	I6164 = NAND(WX2076, I6163)
--	I6165 = NAND(WX2140, I6163)
--	I6162 = NAND(I6164, I6165)
--	I6170 = NAND(I6146, I6162)
--	I6171 = NAND(I6146, I6170)
--	I6172 = NAND(I6162, I6170)
--	WX2198 = NAND(I6171, I6172)
--	I6179 = NAND(WX2294, WX1950)
--	I6180 = NAND(WX2294, I6179)
--	I6181 = NAND(WX1950, I6179)
--	I6178 = NAND(I6180, I6181)
--	I6186 = NAND(WX2014, I6178)
--	I6187 = NAND(WX2014, I6186)
--	I6188 = NAND(I6178, I6186)
--	I6177 = NAND(I6187, I6188)
--	I6194 = NAND(WX2078, WX2142)
--	I6195 = NAND(WX2078, I6194)
--	I6196 = NAND(WX2142, I6194)
--	I6193 = NAND(I6195, I6196)
--	I6201 = NAND(I6177, I6193)
--	I6202 = NAND(I6177, I6201)
--	I6203 = NAND(I6193, I6201)
--	WX2199 = NAND(I6202, I6203)
--	I6210 = NAND(WX2294, WX1952)
--	I6211 = NAND(WX2294, I6210)
--	I6212 = NAND(WX1952, I6210)
--	I6209 = NAND(I6211, I6212)
--	I6217 = NAND(WX2016, I6209)
--	I6218 = NAND(WX2016, I6217)
--	I6219 = NAND(I6209, I6217)
--	I6208 = NAND(I6218, I6219)
--	I6225 = NAND(WX2080, WX2144)
--	I6226 = NAND(WX2080, I6225)
--	I6227 = NAND(WX2144, I6225)
--	I6224 = NAND(I6226, I6227)
--	I6232 = NAND(I6208, I6224)
--	I6233 = NAND(I6208, I6232)
--	I6234 = NAND(I6224, I6232)
--	WX2200 = NAND(I6233, I6234)
--	I6241 = NAND(WX2294, WX1954)
--	I6242 = NAND(WX2294, I6241)
--	I6243 = NAND(WX1954, I6241)
--	I6240 = NAND(I6242, I6243)
--	I6248 = NAND(WX2018, I6240)
--	I6249 = NAND(WX2018, I6248)
--	I6250 = NAND(I6240, I6248)
--	I6239 = NAND(I6249, I6250)
--	I6256 = NAND(WX2082, WX2146)
--	I6257 = NAND(WX2082, I6256)
--	I6258 = NAND(WX2146, I6256)
--	I6255 = NAND(I6257, I6258)
--	I6263 = NAND(I6239, I6255)
--	I6264 = NAND(I6239, I6263)
--	I6265 = NAND(I6255, I6263)
--	WX2201 = NAND(I6264, I6265)
--	I6272 = NAND(WX2294, WX1956)
--	I6273 = NAND(WX2294, I6272)
--	I6274 = NAND(WX1956, I6272)
--	I6271 = NAND(I6273, I6274)
--	I6279 = NAND(WX2020, I6271)
--	I6280 = NAND(WX2020, I6279)
--	I6281 = NAND(I6271, I6279)
--	I6270 = NAND(I6280, I6281)
--	I6287 = NAND(WX2084, WX2148)
--	I6288 = NAND(WX2084, I6287)
--	I6289 = NAND(WX2148, I6287)
--	I6286 = NAND(I6288, I6289)
--	I6294 = NAND(I6270, I6286)
--	I6295 = NAND(I6270, I6294)
--	I6296 = NAND(I6286, I6294)
--	WX2202 = NAND(I6295, I6296)
--	I6303 = NAND(WX2294, WX1958)
--	I6304 = NAND(WX2294, I6303)
--	I6305 = NAND(WX1958, I6303)
--	I6302 = NAND(I6304, I6305)
--	I6310 = NAND(WX2022, I6302)
--	I6311 = NAND(WX2022, I6310)
--	I6312 = NAND(I6302, I6310)
--	I6301 = NAND(I6311, I6312)
--	I6318 = NAND(WX2086, WX2150)
--	I6319 = NAND(WX2086, I6318)
--	I6320 = NAND(WX2150, I6318)
--	I6317 = NAND(I6319, I6320)
--	I6325 = NAND(I6301, I6317)
--	I6326 = NAND(I6301, I6325)
--	I6327 = NAND(I6317, I6325)
--	WX2203 = NAND(I6326, I6327)
--	I6334 = NAND(WX2294, WX1960)
--	I6335 = NAND(WX2294, I6334)
--	I6336 = NAND(WX1960, I6334)
--	I6333 = NAND(I6335, I6336)
--	I6341 = NAND(WX2024, I6333)
--	I6342 = NAND(WX2024, I6341)
--	I6343 = NAND(I6333, I6341)
--	I6332 = NAND(I6342, I6343)
--	I6349 = NAND(WX2088, WX2152)
--	I6350 = NAND(WX2088, I6349)
--	I6351 = NAND(WX2152, I6349)
--	I6348 = NAND(I6350, I6351)
--	I6356 = NAND(I6332, I6348)
--	I6357 = NAND(I6332, I6356)
--	I6358 = NAND(I6348, I6356)
--	WX2204 = NAND(I6357, I6358)
--	I6365 = NAND(WX2294, WX1962)
--	I6366 = NAND(WX2294, I6365)
--	I6367 = NAND(WX1962, I6365)
--	I6364 = NAND(I6366, I6367)
--	I6372 = NAND(WX2026, I6364)
--	I6373 = NAND(WX2026, I6372)
--	I6374 = NAND(I6364, I6372)
--	I6363 = NAND(I6373, I6374)
--	I6380 = NAND(WX2090, WX2154)
--	I6381 = NAND(WX2090, I6380)
--	I6382 = NAND(WX2154, I6380)
--	I6379 = NAND(I6381, I6382)
--	I6387 = NAND(I6363, I6379)
--	I6388 = NAND(I6363, I6387)
--	I6389 = NAND(I6379, I6387)
--	WX2205 = NAND(I6388, I6389)
--	I6396 = NAND(WX2294, WX1964)
--	I6397 = NAND(WX2294, I6396)
--	I6398 = NAND(WX1964, I6396)
--	I6395 = NAND(I6397, I6398)
--	I6403 = NAND(WX2028, I6395)
--	I6404 = NAND(WX2028, I6403)
--	I6405 = NAND(I6395, I6403)
--	I6394 = NAND(I6404, I6405)
--	I6411 = NAND(WX2092, WX2156)
--	I6412 = NAND(WX2092, I6411)
--	I6413 = NAND(WX2156, I6411)
--	I6410 = NAND(I6412, I6413)
--	I6418 = NAND(I6394, I6410)
--	I6419 = NAND(I6394, I6418)
--	I6420 = NAND(I6410, I6418)
--	WX2206 = NAND(I6419, I6420)
--	I6427 = NAND(WX2294, WX1966)
--	I6428 = NAND(WX2294, I6427)
--	I6429 = NAND(WX1966, I6427)
--	I6426 = NAND(I6428, I6429)
--	I6434 = NAND(WX2030, I6426)
--	I6435 = NAND(WX2030, I6434)
--	I6436 = NAND(I6426, I6434)
--	I6425 = NAND(I6435, I6436)
--	I6442 = NAND(WX2094, WX2158)
--	I6443 = NAND(WX2094, I6442)
--	I6444 = NAND(WX2158, I6442)
--	I6441 = NAND(I6443, I6444)
--	I6449 = NAND(I6425, I6441)
--	I6450 = NAND(I6425, I6449)
--	I6451 = NAND(I6441, I6449)
--	WX2207 = NAND(I6450, I6451)
--	I6458 = NAND(WX2294, WX1968)
--	I6459 = NAND(WX2294, I6458)
--	I6460 = NAND(WX1968, I6458)
--	I6457 = NAND(I6459, I6460)
--	I6465 = NAND(WX2032, I6457)
--	I6466 = NAND(WX2032, I6465)
--	I6467 = NAND(I6457, I6465)
--	I6456 = NAND(I6466, I6467)
--	I6473 = NAND(WX2096, WX2160)
--	I6474 = NAND(WX2096, I6473)
--	I6475 = NAND(WX2160, I6473)
--	I6472 = NAND(I6474, I6475)
--	I6480 = NAND(I6456, I6472)
--	I6481 = NAND(I6456, I6480)
--	I6482 = NAND(I6472, I6480)
--	WX2208 = NAND(I6481, I6482)
--	I6489 = NAND(WX2295, WX1970)
--	I6490 = NAND(WX2295, I6489)
--	I6491 = NAND(WX1970, I6489)
--	I6488 = NAND(I6490, I6491)
--	I6496 = NAND(WX2034, I6488)
--	I6497 = NAND(WX2034, I6496)
--	I6498 = NAND(I6488, I6496)
--	I6487 = NAND(I6497, I6498)
--	I6504 = NAND(WX2098, WX2162)
--	I6505 = NAND(WX2098, I6504)
--	I6506 = NAND(WX2162, I6504)
--	I6503 = NAND(I6505, I6506)
--	I6511 = NAND(I6487, I6503)
--	I6512 = NAND(I6487, I6511)
--	I6513 = NAND(I6503, I6511)
--	WX2209 = NAND(I6512, I6513)
--	I6520 = NAND(WX2295, WX1972)
--	I6521 = NAND(WX2295, I6520)
--	I6522 = NAND(WX1972, I6520)
--	I6519 = NAND(I6521, I6522)
--	I6527 = NAND(WX2036, I6519)
--	I6528 = NAND(WX2036, I6527)
--	I6529 = NAND(I6519, I6527)
--	I6518 = NAND(I6528, I6529)
--	I6535 = NAND(WX2100, WX2164)
--	I6536 = NAND(WX2100, I6535)
--	I6537 = NAND(WX2164, I6535)
--	I6534 = NAND(I6536, I6537)
--	I6542 = NAND(I6518, I6534)
--	I6543 = NAND(I6518, I6542)
--	I6544 = NAND(I6534, I6542)
--	WX2210 = NAND(I6543, I6544)
--	I6551 = NAND(WX2295, WX1974)
--	I6552 = NAND(WX2295, I6551)
--	I6553 = NAND(WX1974, I6551)
--	I6550 = NAND(I6552, I6553)
--	I6558 = NAND(WX2038, I6550)
--	I6559 = NAND(WX2038, I6558)
--	I6560 = NAND(I6550, I6558)
--	I6549 = NAND(I6559, I6560)
--	I6566 = NAND(WX2102, WX2166)
--	I6567 = NAND(WX2102, I6566)
--	I6568 = NAND(WX2166, I6566)
--	I6565 = NAND(I6567, I6568)
--	I6573 = NAND(I6549, I6565)
--	I6574 = NAND(I6549, I6573)
--	I6575 = NAND(I6565, I6573)
--	WX2211 = NAND(I6574, I6575)
--	I6582 = NAND(WX2295, WX1976)
--	I6583 = NAND(WX2295, I6582)
--	I6584 = NAND(WX1976, I6582)
--	I6581 = NAND(I6583, I6584)
--	I6589 = NAND(WX2040, I6581)
--	I6590 = NAND(WX2040, I6589)
--	I6591 = NAND(I6581, I6589)
--	I6580 = NAND(I6590, I6591)
--	I6597 = NAND(WX2104, WX2168)
--	I6598 = NAND(WX2104, I6597)
--	I6599 = NAND(WX2168, I6597)
--	I6596 = NAND(I6598, I6599)
--	I6604 = NAND(I6580, I6596)
--	I6605 = NAND(I6580, I6604)
--	I6606 = NAND(I6596, I6604)
--	WX2212 = NAND(I6605, I6606)
--	I6613 = NAND(WX2295, WX1978)
--	I6614 = NAND(WX2295, I6613)
--	I6615 = NAND(WX1978, I6613)
--	I6612 = NAND(I6614, I6615)
--	I6620 = NAND(WX2042, I6612)
--	I6621 = NAND(WX2042, I6620)
--	I6622 = NAND(I6612, I6620)
--	I6611 = NAND(I6621, I6622)
--	I6628 = NAND(WX2106, WX2170)
--	I6629 = NAND(WX2106, I6628)
--	I6630 = NAND(WX2170, I6628)
--	I6627 = NAND(I6629, I6630)
--	I6635 = NAND(I6611, I6627)
--	I6636 = NAND(I6611, I6635)
--	I6637 = NAND(I6627, I6635)
--	WX2213 = NAND(I6636, I6637)
--	I6644 = NAND(WX2295, WX1980)
--	I6645 = NAND(WX2295, I6644)
--	I6646 = NAND(WX1980, I6644)
--	I6643 = NAND(I6645, I6646)
--	I6651 = NAND(WX2044, I6643)
--	I6652 = NAND(WX2044, I6651)
--	I6653 = NAND(I6643, I6651)
--	I6642 = NAND(I6652, I6653)
--	I6659 = NAND(WX2108, WX2172)
--	I6660 = NAND(WX2108, I6659)
--	I6661 = NAND(WX2172, I6659)
--	I6658 = NAND(I6660, I6661)
--	I6666 = NAND(I6642, I6658)
--	I6667 = NAND(I6642, I6666)
--	I6668 = NAND(I6658, I6666)
--	WX2214 = NAND(I6667, I6668)
--	I6675 = NAND(WX2295, WX1982)
--	I6676 = NAND(WX2295, I6675)
--	I6677 = NAND(WX1982, I6675)
--	I6674 = NAND(I6676, I6677)
--	I6682 = NAND(WX2046, I6674)
--	I6683 = NAND(WX2046, I6682)
--	I6684 = NAND(I6674, I6682)
--	I6673 = NAND(I6683, I6684)
--	I6690 = NAND(WX2110, WX2174)
--	I6691 = NAND(WX2110, I6690)
--	I6692 = NAND(WX2174, I6690)
--	I6689 = NAND(I6691, I6692)
--	I6697 = NAND(I6673, I6689)
--	I6698 = NAND(I6673, I6697)
--	I6699 = NAND(I6689, I6697)
--	WX2215 = NAND(I6698, I6699)
--	I6706 = NAND(WX2295, WX1984)
--	I6707 = NAND(WX2295, I6706)
--	I6708 = NAND(WX1984, I6706)
--	I6705 = NAND(I6707, I6708)
--	I6713 = NAND(WX2048, I6705)
--	I6714 = NAND(WX2048, I6713)
--	I6715 = NAND(I6705, I6713)
--	I6704 = NAND(I6714, I6715)
--	I6721 = NAND(WX2112, WX2176)
--	I6722 = NAND(WX2112, I6721)
--	I6723 = NAND(WX2176, I6721)
--	I6720 = NAND(I6722, I6723)
--	I6728 = NAND(I6704, I6720)
--	I6729 = NAND(I6704, I6728)
--	I6730 = NAND(I6720, I6728)
--	WX2216 = NAND(I6729, I6730)
--	I6737 = NAND(WX2295, WX1986)
--	I6738 = NAND(WX2295, I6737)
--	I6739 = NAND(WX1986, I6737)
--	I6736 = NAND(I6738, I6739)
--	I6744 = NAND(WX2050, I6736)
--	I6745 = NAND(WX2050, I6744)
--	I6746 = NAND(I6736, I6744)
--	I6735 = NAND(I6745, I6746)
--	I6752 = NAND(WX2114, WX2178)
--	I6753 = NAND(WX2114, I6752)
--	I6754 = NAND(WX2178, I6752)
--	I6751 = NAND(I6753, I6754)
--	I6759 = NAND(I6735, I6751)
--	I6760 = NAND(I6735, I6759)
--	I6761 = NAND(I6751, I6759)
--	WX2217 = NAND(I6760, I6761)
--	I6768 = NAND(WX2295, WX1988)
--	I6769 = NAND(WX2295, I6768)
--	I6770 = NAND(WX1988, I6768)
--	I6767 = NAND(I6769, I6770)
--	I6775 = NAND(WX2052, I6767)
--	I6776 = NAND(WX2052, I6775)
--	I6777 = NAND(I6767, I6775)
--	I6766 = NAND(I6776, I6777)
--	I6783 = NAND(WX2116, WX2180)
--	I6784 = NAND(WX2116, I6783)
--	I6785 = NAND(WX2180, I6783)
--	I6782 = NAND(I6784, I6785)
--	I6790 = NAND(I6766, I6782)
--	I6791 = NAND(I6766, I6790)
--	I6792 = NAND(I6782, I6790)
--	WX2218 = NAND(I6791, I6792)
--	I6799 = NAND(WX2295, WX1990)
--	I6800 = NAND(WX2295, I6799)
--	I6801 = NAND(WX1990, I6799)
--	I6798 = NAND(I6800, I6801)
--	I6806 = NAND(WX2054, I6798)
--	I6807 = NAND(WX2054, I6806)
--	I6808 = NAND(I6798, I6806)
--	I6797 = NAND(I6807, I6808)
--	I6814 = NAND(WX2118, WX2182)
--	I6815 = NAND(WX2118, I6814)
--	I6816 = NAND(WX2182, I6814)
--	I6813 = NAND(I6815, I6816)
--	I6821 = NAND(I6797, I6813)
--	I6822 = NAND(I6797, I6821)
--	I6823 = NAND(I6813, I6821)
--	WX2219 = NAND(I6822, I6823)
--	I6830 = NAND(WX2295, WX1992)
--	I6831 = NAND(WX2295, I6830)
--	I6832 = NAND(WX1992, I6830)
--	I6829 = NAND(I6831, I6832)
--	I6837 = NAND(WX2056, I6829)
--	I6838 = NAND(WX2056, I6837)
--	I6839 = NAND(I6829, I6837)
--	I6828 = NAND(I6838, I6839)
--	I6845 = NAND(WX2120, WX2184)
--	I6846 = NAND(WX2120, I6845)
--	I6847 = NAND(WX2184, I6845)
--	I6844 = NAND(I6846, I6847)
--	I6852 = NAND(I6828, I6844)
--	I6853 = NAND(I6828, I6852)
--	I6854 = NAND(I6844, I6852)
--	WX2220 = NAND(I6853, I6854)
--	I6861 = NAND(WX2295, WX1994)
--	I6862 = NAND(WX2295, I6861)
--	I6863 = NAND(WX1994, I6861)
--	I6860 = NAND(I6862, I6863)
--	I6868 = NAND(WX2058, I6860)
--	I6869 = NAND(WX2058, I6868)
--	I6870 = NAND(I6860, I6868)
--	I6859 = NAND(I6869, I6870)
--	I6876 = NAND(WX2122, WX2186)
--	I6877 = NAND(WX2122, I6876)
--	I6878 = NAND(WX2186, I6876)
--	I6875 = NAND(I6877, I6878)
--	I6883 = NAND(I6859, I6875)
--	I6884 = NAND(I6859, I6883)
--	I6885 = NAND(I6875, I6883)
--	WX2221 = NAND(I6884, I6885)
--	I6892 = NAND(WX2295, WX1996)
--	I6893 = NAND(WX2295, I6892)
--	I6894 = NAND(WX1996, I6892)
--	I6891 = NAND(I6893, I6894)
--	I6899 = NAND(WX2060, I6891)
--	I6900 = NAND(WX2060, I6899)
--	I6901 = NAND(I6891, I6899)
--	I6890 = NAND(I6900, I6901)
--	I6907 = NAND(WX2124, WX2188)
--	I6908 = NAND(WX2124, I6907)
--	I6909 = NAND(WX2188, I6907)
--	I6906 = NAND(I6908, I6909)
--	I6914 = NAND(I6890, I6906)
--	I6915 = NAND(I6890, I6914)
--	I6916 = NAND(I6906, I6914)
--	WX2222 = NAND(I6915, I6916)
--	I6923 = NAND(WX2295, WX1998)
--	I6924 = NAND(WX2295, I6923)
--	I6925 = NAND(WX1998, I6923)
--	I6922 = NAND(I6924, I6925)
--	I6930 = NAND(WX2062, I6922)
--	I6931 = NAND(WX2062, I6930)
--	I6932 = NAND(I6922, I6930)
--	I6921 = NAND(I6931, I6932)
--	I6938 = NAND(WX2126, WX2190)
--	I6939 = NAND(WX2126, I6938)
--	I6940 = NAND(WX2190, I6938)
--	I6937 = NAND(I6939, I6940)
--	I6945 = NAND(I6921, I6937)
--	I6946 = NAND(I6921, I6945)
--	I6947 = NAND(I6937, I6945)
--	WX2223 = NAND(I6946, I6947)
--	I6954 = NAND(WX2295, WX2000)
--	I6955 = NAND(WX2295, I6954)
--	I6956 = NAND(WX2000, I6954)
--	I6953 = NAND(I6955, I6956)
--	I6961 = NAND(WX2064, I6953)
--	I6962 = NAND(WX2064, I6961)
--	I6963 = NAND(I6953, I6961)
--	I6952 = NAND(I6962, I6963)
--	I6969 = NAND(WX2128, WX2192)
--	I6970 = NAND(WX2128, I6969)
--	I6971 = NAND(WX2192, I6969)
--	I6968 = NAND(I6970, I6971)
--	I6976 = NAND(I6952, I6968)
--	I6977 = NAND(I6952, I6976)
--	I6978 = NAND(I6968, I6976)
--	WX2224 = NAND(I6977, I6978)
--	I7057 = NAND(WX1873, WX1778)
--	I7058 = NAND(WX1873, I7057)
--	I7059 = NAND(WX1778, I7057)
--	WX2299 = NAND(I7058, I7059)
--	I7070 = NAND(WX1874, WX1780)
--	I7071 = NAND(WX1874, I7070)
--	I7072 = NAND(WX1780, I7070)
--	WX2306 = NAND(I7071, I7072)
--	I7083 = NAND(WX1875, WX1782)
--	I7084 = NAND(WX1875, I7083)
--	I7085 = NAND(WX1782, I7083)
--	WX2313 = NAND(I7084, I7085)
--	I7096 = NAND(WX1876, WX1784)
--	I7097 = NAND(WX1876, I7096)
--	I7098 = NAND(WX1784, I7096)
--	WX2320 = NAND(I7097, I7098)
--	I7109 = NAND(WX1877, WX1786)
--	I7110 = NAND(WX1877, I7109)
--	I7111 = NAND(WX1786, I7109)
--	WX2327 = NAND(I7110, I7111)
--	I7122 = NAND(WX1878, WX1788)
--	I7123 = NAND(WX1878, I7122)
--	I7124 = NAND(WX1788, I7122)
--	WX2334 = NAND(I7123, I7124)
--	I7135 = NAND(WX1879, WX1790)
--	I7136 = NAND(WX1879, I7135)
--	I7137 = NAND(WX1790, I7135)
--	WX2341 = NAND(I7136, I7137)
--	I7148 = NAND(WX1880, WX1792)
--	I7149 = NAND(WX1880, I7148)
--	I7150 = NAND(WX1792, I7148)
--	WX2348 = NAND(I7149, I7150)
--	I7161 = NAND(WX1881, WX1794)
--	I7162 = NAND(WX1881, I7161)
--	I7163 = NAND(WX1794, I7161)
--	WX2355 = NAND(I7162, I7163)
--	I7174 = NAND(WX1882, WX1796)
--	I7175 = NAND(WX1882, I7174)
--	I7176 = NAND(WX1796, I7174)
--	WX2362 = NAND(I7175, I7176)
--	I7187 = NAND(WX1883, WX1798)
--	I7188 = NAND(WX1883, I7187)
--	I7189 = NAND(WX1798, I7187)
--	WX2369 = NAND(I7188, I7189)
--	I7200 = NAND(WX1884, WX1800)
--	I7201 = NAND(WX1884, I7200)
--	I7202 = NAND(WX1800, I7200)
--	WX2376 = NAND(I7201, I7202)
--	I7213 = NAND(WX1885, WX1802)
--	I7214 = NAND(WX1885, I7213)
--	I7215 = NAND(WX1802, I7213)
--	WX2383 = NAND(I7214, I7215)
--	I7226 = NAND(WX1886, WX1804)
--	I7227 = NAND(WX1886, I7226)
--	I7228 = NAND(WX1804, I7226)
--	WX2390 = NAND(I7227, I7228)
--	I7239 = NAND(WX1887, WX1806)
--	I7240 = NAND(WX1887, I7239)
--	I7241 = NAND(WX1806, I7239)
--	WX2397 = NAND(I7240, I7241)
--	I7252 = NAND(WX1888, WX1808)
--	I7253 = NAND(WX1888, I7252)
--	I7254 = NAND(WX1808, I7252)
--	WX2404 = NAND(I7253, I7254)
--	I7265 = NAND(WX1889, WX1810)
--	I7266 = NAND(WX1889, I7265)
--	I7267 = NAND(WX1810, I7265)
--	WX2411 = NAND(I7266, I7267)
--	I7278 = NAND(WX1890, WX1812)
--	I7279 = NAND(WX1890, I7278)
--	I7280 = NAND(WX1812, I7278)
--	WX2418 = NAND(I7279, I7280)
--	I7291 = NAND(WX1891, WX1814)
--	I7292 = NAND(WX1891, I7291)
--	I7293 = NAND(WX1814, I7291)
--	WX2425 = NAND(I7292, I7293)
--	I7304 = NAND(WX1892, WX1816)
--	I7305 = NAND(WX1892, I7304)
--	I7306 = NAND(WX1816, I7304)
--	WX2432 = NAND(I7305, I7306)
--	I7317 = NAND(WX1893, WX1818)
--	I7318 = NAND(WX1893, I7317)
--	I7319 = NAND(WX1818, I7317)
--	WX2439 = NAND(I7318, I7319)
--	I7330 = NAND(WX1894, WX1820)
--	I7331 = NAND(WX1894, I7330)
--	I7332 = NAND(WX1820, I7330)
--	WX2446 = NAND(I7331, I7332)
--	I7343 = NAND(WX1895, WX1822)
--	I7344 = NAND(WX1895, I7343)
--	I7345 = NAND(WX1822, I7343)
--	WX2453 = NAND(I7344, I7345)
--	I7356 = NAND(WX1896, WX1824)
--	I7357 = NAND(WX1896, I7356)
--	I7358 = NAND(WX1824, I7356)
--	WX2460 = NAND(I7357, I7358)
--	I7369 = NAND(WX1897, WX1826)
--	I7370 = NAND(WX1897, I7369)
--	I7371 = NAND(WX1826, I7369)
--	WX2467 = NAND(I7370, I7371)
--	I7382 = NAND(WX1898, WX1828)
--	I7383 = NAND(WX1898, I7382)
--	I7384 = NAND(WX1828, I7382)
--	WX2474 = NAND(I7383, I7384)
--	I7395 = NAND(WX1899, WX1830)
--	I7396 = NAND(WX1899, I7395)
--	I7397 = NAND(WX1830, I7395)
--	WX2481 = NAND(I7396, I7397)
--	I7408 = NAND(WX1900, WX1832)
--	I7409 = NAND(WX1900, I7408)
--	I7410 = NAND(WX1832, I7408)
--	WX2488 = NAND(I7409, I7410)
--	I7421 = NAND(WX1901, WX1834)
--	I7422 = NAND(WX1901, I7421)
--	I7423 = NAND(WX1834, I7421)
--	WX2495 = NAND(I7422, I7423)
--	I7434 = NAND(WX1902, WX1836)
--	I7435 = NAND(WX1902, I7434)
--	I7436 = NAND(WX1836, I7434)
--	WX2502 = NAND(I7435, I7436)
--	I7447 = NAND(WX1903, WX1838)
--	I7448 = NAND(WX1903, I7447)
--	I7449 = NAND(WX1838, I7447)
--	WX2509 = NAND(I7448, I7449)
--	I7460 = NAND(WX1904, WX1840)
--	I7461 = NAND(WX1904, I7460)
--	I7462 = NAND(WX1840, I7460)
--	WX2516 = NAND(I7461, I7462)
--	I7475 = NAND(WX1920, CRC_OUT_8_31)
--	I7476 = NAND(WX1920, I7475)
--	I7477 = NAND(CRC_OUT_8_31, I7475)
--	I7474 = NAND(I7476, I7477)
--	I7482 = NAND(CRC_OUT_8_15, I7474)
--	I7483 = NAND(CRC_OUT_8_15, I7482)
--	I7484 = NAND(I7474, I7482)
--	WX2524 = NAND(I7483, I7484)
--	I7490 = NAND(WX1925, CRC_OUT_8_31)
--	I7491 = NAND(WX1925, I7490)
--	I7492 = NAND(CRC_OUT_8_31, I7490)
--	I7489 = NAND(I7491, I7492)
--	I7497 = NAND(CRC_OUT_8_10, I7489)
--	I7498 = NAND(CRC_OUT_8_10, I7497)
--	I7499 = NAND(I7489, I7497)
--	WX2525 = NAND(I7498, I7499)
--	I7505 = NAND(WX1932, CRC_OUT_8_31)
--	I7506 = NAND(WX1932, I7505)
--	I7507 = NAND(CRC_OUT_8_31, I7505)
--	I7504 = NAND(I7506, I7507)
--	I7512 = NAND(CRC_OUT_8_3, I7504)
--	I7513 = NAND(CRC_OUT_8_3, I7512)
--	I7514 = NAND(I7504, I7512)
--	WX2526 = NAND(I7513, I7514)
--	I7519 = NAND(WX1936, CRC_OUT_8_31)
--	I7520 = NAND(WX1936, I7519)
--	I7521 = NAND(CRC_OUT_8_31, I7519)
--	WX2527 = NAND(I7520, I7521)
--	I7526 = NAND(WX1905, CRC_OUT_8_30)
--	I7527 = NAND(WX1905, I7526)
--	I7528 = NAND(CRC_OUT_8_30, I7526)
--	WX2528 = NAND(I7527, I7528)
--	I7533 = NAND(WX1906, CRC_OUT_8_29)
--	I7534 = NAND(WX1906, I7533)
--	I7535 = NAND(CRC_OUT_8_29, I7533)
--	WX2529 = NAND(I7534, I7535)
--	I7540 = NAND(WX1907, CRC_OUT_8_28)
--	I7541 = NAND(WX1907, I7540)
--	I7542 = NAND(CRC_OUT_8_28, I7540)
--	WX2530 = NAND(I7541, I7542)
--	I7547 = NAND(WX1908, CRC_OUT_8_27)
--	I7548 = NAND(WX1908, I7547)
--	I7549 = NAND(CRC_OUT_8_27, I7547)
--	WX2531 = NAND(I7548, I7549)
--	I7554 = NAND(WX1909, CRC_OUT_8_26)
--	I7555 = NAND(WX1909, I7554)
--	I7556 = NAND(CRC_OUT_8_26, I7554)
--	WX2532 = NAND(I7555, I7556)
--	I7561 = NAND(WX1910, CRC_OUT_8_25)
--	I7562 = NAND(WX1910, I7561)
--	I7563 = NAND(CRC_OUT_8_25, I7561)
--	WX2533 = NAND(I7562, I7563)
--	I7568 = NAND(WX1911, CRC_OUT_8_24)
--	I7569 = NAND(WX1911, I7568)
--	I7570 = NAND(CRC_OUT_8_24, I7568)
--	WX2534 = NAND(I7569, I7570)
--	I7575 = NAND(WX1912, CRC_OUT_8_23)
--	I7576 = NAND(WX1912, I7575)
--	I7577 = NAND(CRC_OUT_8_23, I7575)
--	WX2535 = NAND(I7576, I7577)
--	I7582 = NAND(WX1913, CRC_OUT_8_22)
--	I7583 = NAND(WX1913, I7582)
--	I7584 = NAND(CRC_OUT_8_22, I7582)
--	WX2536 = NAND(I7583, I7584)
--	I7589 = NAND(WX1914, CRC_OUT_8_21)
--	I7590 = NAND(WX1914, I7589)
--	I7591 = NAND(CRC_OUT_8_21, I7589)
--	WX2537 = NAND(I7590, I7591)
--	I7596 = NAND(WX1915, CRC_OUT_8_20)
--	I7597 = NAND(WX1915, I7596)
--	I7598 = NAND(CRC_OUT_8_20, I7596)
--	WX2538 = NAND(I7597, I7598)
--	I7603 = NAND(WX1916, CRC_OUT_8_19)
--	I7604 = NAND(WX1916, I7603)
--	I7605 = NAND(CRC_OUT_8_19, I7603)
--	WX2539 = NAND(I7604, I7605)
--	I7610 = NAND(WX1917, CRC_OUT_8_18)
--	I7611 = NAND(WX1917, I7610)
--	I7612 = NAND(CRC_OUT_8_18, I7610)
--	WX2540 = NAND(I7611, I7612)
--	I7617 = NAND(WX1918, CRC_OUT_8_17)
--	I7618 = NAND(WX1918, I7617)
--	I7619 = NAND(CRC_OUT_8_17, I7617)
--	WX2541 = NAND(I7618, I7619)
--	I7624 = NAND(WX1919, CRC_OUT_8_16)
--	I7625 = NAND(WX1919, I7624)
--	I7626 = NAND(CRC_OUT_8_16, I7624)
--	WX2542 = NAND(I7625, I7626)
--	I7631 = NAND(WX1921, CRC_OUT_8_14)
--	I7632 = NAND(WX1921, I7631)
--	I7633 = NAND(CRC_OUT_8_14, I7631)
--	WX2543 = NAND(I7632, I7633)
--	I7638 = NAND(WX1922, CRC_OUT_8_13)
--	I7639 = NAND(WX1922, I7638)
--	I7640 = NAND(CRC_OUT_8_13, I7638)
--	WX2544 = NAND(I7639, I7640)
--	I7645 = NAND(WX1923, CRC_OUT_8_12)
--	I7646 = NAND(WX1923, I7645)
--	I7647 = NAND(CRC_OUT_8_12, I7645)
--	WX2545 = NAND(I7646, I7647)
--	I7652 = NAND(WX1924, CRC_OUT_8_11)
--	I7653 = NAND(WX1924, I7652)
--	I7654 = NAND(CRC_OUT_8_11, I7652)
--	WX2546 = NAND(I7653, I7654)
--	I7659 = NAND(WX1926, CRC_OUT_8_9)
--	I7660 = NAND(WX1926, I7659)
--	I7661 = NAND(CRC_OUT_8_9, I7659)
--	WX2547 = NAND(I7660, I7661)
--	I7666 = NAND(WX1927, CRC_OUT_8_8)
--	I7667 = NAND(WX1927, I7666)
--	I7668 = NAND(CRC_OUT_8_8, I7666)
--	WX2548 = NAND(I7667, I7668)
--	I7673 = NAND(WX1928, CRC_OUT_8_7)
--	I7674 = NAND(WX1928, I7673)
--	I7675 = NAND(CRC_OUT_8_7, I7673)
--	WX2549 = NAND(I7674, I7675)
--	I7680 = NAND(WX1929, CRC_OUT_8_6)
--	I7681 = NAND(WX1929, I7680)
--	I7682 = NAND(CRC_OUT_8_6, I7680)
--	WX2550 = NAND(I7681, I7682)
--	I7687 = NAND(WX1930, CRC_OUT_8_5)
--	I7688 = NAND(WX1930, I7687)
--	I7689 = NAND(CRC_OUT_8_5, I7687)
--	WX2551 = NAND(I7688, I7689)
--	I7694 = NAND(WX1931, CRC_OUT_8_4)
--	I7695 = NAND(WX1931, I7694)
--	I7696 = NAND(CRC_OUT_8_4, I7694)
--	WX2552 = NAND(I7695, I7696)
--	I7701 = NAND(WX1933, CRC_OUT_8_2)
--	I7702 = NAND(WX1933, I7701)
--	I7703 = NAND(CRC_OUT_8_2, I7701)
--	WX2553 = NAND(I7702, I7703)
--	I7708 = NAND(WX1934, CRC_OUT_8_1)
--	I7709 = NAND(WX1934, I7708)
--	I7710 = NAND(CRC_OUT_8_1, I7708)
--	WX2554 = NAND(I7709, I7710)
--	I7715 = NAND(WX1935, CRC_OUT_8_0)
--	I7716 = NAND(WX1935, I7715)
--	I7717 = NAND(CRC_OUT_8_0, I7715)
--	WX2555 = NAND(I7716, I7717)
--	I9998 = NAND(WX3587, WX3231)
--	I9999 = NAND(WX3587, I9998)
--	I10000 = NAND(WX3231, I9998)
--	I9997 = NAND(I9999, I10000)
--	I10005 = NAND(WX3295, I9997)
--	I10006 = NAND(WX3295, I10005)
--	I10007 = NAND(I9997, I10005)
--	I9996 = NAND(I10006, I10007)
--	I10013 = NAND(WX3359, WX3423)
--	I10014 = NAND(WX3359, I10013)
--	I10015 = NAND(WX3423, I10013)
--	I10012 = NAND(I10014, I10015)
--	I10020 = NAND(I9996, I10012)
--	I10021 = NAND(I9996, I10020)
--	I10022 = NAND(I10012, I10020)
--	WX3486 = NAND(I10021, I10022)
--	I10029 = NAND(WX3587, WX3233)
--	I10030 = NAND(WX3587, I10029)
--	I10031 = NAND(WX3233, I10029)
--	I10028 = NAND(I10030, I10031)
--	I10036 = NAND(WX3297, I10028)
--	I10037 = NAND(WX3297, I10036)
--	I10038 = NAND(I10028, I10036)
--	I10027 = NAND(I10037, I10038)
--	I10044 = NAND(WX3361, WX3425)
--	I10045 = NAND(WX3361, I10044)
--	I10046 = NAND(WX3425, I10044)
--	I10043 = NAND(I10045, I10046)
--	I10051 = NAND(I10027, I10043)
--	I10052 = NAND(I10027, I10051)
--	I10053 = NAND(I10043, I10051)
--	WX3487 = NAND(I10052, I10053)
--	I10060 = NAND(WX3587, WX3235)
--	I10061 = NAND(WX3587, I10060)
--	I10062 = NAND(WX3235, I10060)
--	I10059 = NAND(I10061, I10062)
--	I10067 = NAND(WX3299, I10059)
--	I10068 = NAND(WX3299, I10067)
--	I10069 = NAND(I10059, I10067)
--	I10058 = NAND(I10068, I10069)
--	I10075 = NAND(WX3363, WX3427)
--	I10076 = NAND(WX3363, I10075)
--	I10077 = NAND(WX3427, I10075)
--	I10074 = NAND(I10076, I10077)
--	I10082 = NAND(I10058, I10074)
--	I10083 = NAND(I10058, I10082)
--	I10084 = NAND(I10074, I10082)
--	WX3488 = NAND(I10083, I10084)
--	I10091 = NAND(WX3587, WX3237)
--	I10092 = NAND(WX3587, I10091)
--	I10093 = NAND(WX3237, I10091)
--	I10090 = NAND(I10092, I10093)
--	I10098 = NAND(WX3301, I10090)
--	I10099 = NAND(WX3301, I10098)
--	I10100 = NAND(I10090, I10098)
--	I10089 = NAND(I10099, I10100)
--	I10106 = NAND(WX3365, WX3429)
--	I10107 = NAND(WX3365, I10106)
--	I10108 = NAND(WX3429, I10106)
--	I10105 = NAND(I10107, I10108)
--	I10113 = NAND(I10089, I10105)
--	I10114 = NAND(I10089, I10113)
--	I10115 = NAND(I10105, I10113)
--	WX3489 = NAND(I10114, I10115)
--	I10122 = NAND(WX3587, WX3239)
--	I10123 = NAND(WX3587, I10122)
--	I10124 = NAND(WX3239, I10122)
--	I10121 = NAND(I10123, I10124)
--	I10129 = NAND(WX3303, I10121)
--	I10130 = NAND(WX3303, I10129)
--	I10131 = NAND(I10121, I10129)
--	I10120 = NAND(I10130, I10131)
--	I10137 = NAND(WX3367, WX3431)
--	I10138 = NAND(WX3367, I10137)
--	I10139 = NAND(WX3431, I10137)
--	I10136 = NAND(I10138, I10139)
--	I10144 = NAND(I10120, I10136)
--	I10145 = NAND(I10120, I10144)
--	I10146 = NAND(I10136, I10144)
--	WX3490 = NAND(I10145, I10146)
--	I10153 = NAND(WX3587, WX3241)
--	I10154 = NAND(WX3587, I10153)
--	I10155 = NAND(WX3241, I10153)
--	I10152 = NAND(I10154, I10155)
--	I10160 = NAND(WX3305, I10152)
--	I10161 = NAND(WX3305, I10160)
--	I10162 = NAND(I10152, I10160)
--	I10151 = NAND(I10161, I10162)
--	I10168 = NAND(WX3369, WX3433)
--	I10169 = NAND(WX3369, I10168)
--	I10170 = NAND(WX3433, I10168)
--	I10167 = NAND(I10169, I10170)
--	I10175 = NAND(I10151, I10167)
--	I10176 = NAND(I10151, I10175)
--	I10177 = NAND(I10167, I10175)
--	WX3491 = NAND(I10176, I10177)
--	I10184 = NAND(WX3587, WX3243)
--	I10185 = NAND(WX3587, I10184)
--	I10186 = NAND(WX3243, I10184)
--	I10183 = NAND(I10185, I10186)
--	I10191 = NAND(WX3307, I10183)
--	I10192 = NAND(WX3307, I10191)
--	I10193 = NAND(I10183, I10191)
--	I10182 = NAND(I10192, I10193)
--	I10199 = NAND(WX3371, WX3435)
--	I10200 = NAND(WX3371, I10199)
--	I10201 = NAND(WX3435, I10199)
--	I10198 = NAND(I10200, I10201)
--	I10206 = NAND(I10182, I10198)
--	I10207 = NAND(I10182, I10206)
--	I10208 = NAND(I10198, I10206)
--	WX3492 = NAND(I10207, I10208)
--	I10215 = NAND(WX3587, WX3245)
--	I10216 = NAND(WX3587, I10215)
--	I10217 = NAND(WX3245, I10215)
--	I10214 = NAND(I10216, I10217)
--	I10222 = NAND(WX3309, I10214)
--	I10223 = NAND(WX3309, I10222)
--	I10224 = NAND(I10214, I10222)
--	I10213 = NAND(I10223, I10224)
--	I10230 = NAND(WX3373, WX3437)
--	I10231 = NAND(WX3373, I10230)
--	I10232 = NAND(WX3437, I10230)
--	I10229 = NAND(I10231, I10232)
--	I10237 = NAND(I10213, I10229)
--	I10238 = NAND(I10213, I10237)
--	I10239 = NAND(I10229, I10237)
--	WX3493 = NAND(I10238, I10239)
--	I10246 = NAND(WX3587, WX3247)
--	I10247 = NAND(WX3587, I10246)
--	I10248 = NAND(WX3247, I10246)
--	I10245 = NAND(I10247, I10248)
--	I10253 = NAND(WX3311, I10245)
--	I10254 = NAND(WX3311, I10253)
--	I10255 = NAND(I10245, I10253)
--	I10244 = NAND(I10254, I10255)
--	I10261 = NAND(WX3375, WX3439)
--	I10262 = NAND(WX3375, I10261)
--	I10263 = NAND(WX3439, I10261)
--	I10260 = NAND(I10262, I10263)
--	I10268 = NAND(I10244, I10260)
--	I10269 = NAND(I10244, I10268)
--	I10270 = NAND(I10260, I10268)
--	WX3494 = NAND(I10269, I10270)
--	I10277 = NAND(WX3587, WX3249)
--	I10278 = NAND(WX3587, I10277)
--	I10279 = NAND(WX3249, I10277)
--	I10276 = NAND(I10278, I10279)
--	I10284 = NAND(WX3313, I10276)
--	I10285 = NAND(WX3313, I10284)
--	I10286 = NAND(I10276, I10284)
--	I10275 = NAND(I10285, I10286)
--	I10292 = NAND(WX3377, WX3441)
--	I10293 = NAND(WX3377, I10292)
--	I10294 = NAND(WX3441, I10292)
--	I10291 = NAND(I10293, I10294)
--	I10299 = NAND(I10275, I10291)
--	I10300 = NAND(I10275, I10299)
--	I10301 = NAND(I10291, I10299)
--	WX3495 = NAND(I10300, I10301)
--	I10308 = NAND(WX3587, WX3251)
--	I10309 = NAND(WX3587, I10308)
--	I10310 = NAND(WX3251, I10308)
--	I10307 = NAND(I10309, I10310)
--	I10315 = NAND(WX3315, I10307)
--	I10316 = NAND(WX3315, I10315)
--	I10317 = NAND(I10307, I10315)
--	I10306 = NAND(I10316, I10317)
--	I10323 = NAND(WX3379, WX3443)
--	I10324 = NAND(WX3379, I10323)
--	I10325 = NAND(WX3443, I10323)
--	I10322 = NAND(I10324, I10325)
--	I10330 = NAND(I10306, I10322)
--	I10331 = NAND(I10306, I10330)
--	I10332 = NAND(I10322, I10330)
--	WX3496 = NAND(I10331, I10332)
--	I10339 = NAND(WX3587, WX3253)
--	I10340 = NAND(WX3587, I10339)
--	I10341 = NAND(WX3253, I10339)
--	I10338 = NAND(I10340, I10341)
--	I10346 = NAND(WX3317, I10338)
--	I10347 = NAND(WX3317, I10346)
--	I10348 = NAND(I10338, I10346)
--	I10337 = NAND(I10347, I10348)
--	I10354 = NAND(WX3381, WX3445)
--	I10355 = NAND(WX3381, I10354)
--	I10356 = NAND(WX3445, I10354)
--	I10353 = NAND(I10355, I10356)
--	I10361 = NAND(I10337, I10353)
--	I10362 = NAND(I10337, I10361)
--	I10363 = NAND(I10353, I10361)
--	WX3497 = NAND(I10362, I10363)
--	I10370 = NAND(WX3587, WX3255)
--	I10371 = NAND(WX3587, I10370)
--	I10372 = NAND(WX3255, I10370)
--	I10369 = NAND(I10371, I10372)
--	I10377 = NAND(WX3319, I10369)
--	I10378 = NAND(WX3319, I10377)
--	I10379 = NAND(I10369, I10377)
--	I10368 = NAND(I10378, I10379)
--	I10385 = NAND(WX3383, WX3447)
--	I10386 = NAND(WX3383, I10385)
--	I10387 = NAND(WX3447, I10385)
--	I10384 = NAND(I10386, I10387)
--	I10392 = NAND(I10368, I10384)
--	I10393 = NAND(I10368, I10392)
--	I10394 = NAND(I10384, I10392)
--	WX3498 = NAND(I10393, I10394)
--	I10401 = NAND(WX3587, WX3257)
--	I10402 = NAND(WX3587, I10401)
--	I10403 = NAND(WX3257, I10401)
--	I10400 = NAND(I10402, I10403)
--	I10408 = NAND(WX3321, I10400)
--	I10409 = NAND(WX3321, I10408)
--	I10410 = NAND(I10400, I10408)
--	I10399 = NAND(I10409, I10410)
--	I10416 = NAND(WX3385, WX3449)
--	I10417 = NAND(WX3385, I10416)
--	I10418 = NAND(WX3449, I10416)
--	I10415 = NAND(I10417, I10418)
--	I10423 = NAND(I10399, I10415)
--	I10424 = NAND(I10399, I10423)
--	I10425 = NAND(I10415, I10423)
--	WX3499 = NAND(I10424, I10425)
--	I10432 = NAND(WX3587, WX3259)
--	I10433 = NAND(WX3587, I10432)
--	I10434 = NAND(WX3259, I10432)
--	I10431 = NAND(I10433, I10434)
--	I10439 = NAND(WX3323, I10431)
--	I10440 = NAND(WX3323, I10439)
--	I10441 = NAND(I10431, I10439)
--	I10430 = NAND(I10440, I10441)
--	I10447 = NAND(WX3387, WX3451)
--	I10448 = NAND(WX3387, I10447)
--	I10449 = NAND(WX3451, I10447)
--	I10446 = NAND(I10448, I10449)
--	I10454 = NAND(I10430, I10446)
--	I10455 = NAND(I10430, I10454)
--	I10456 = NAND(I10446, I10454)
--	WX3500 = NAND(I10455, I10456)
--	I10463 = NAND(WX3587, WX3261)
--	I10464 = NAND(WX3587, I10463)
--	I10465 = NAND(WX3261, I10463)
--	I10462 = NAND(I10464, I10465)
--	I10470 = NAND(WX3325, I10462)
--	I10471 = NAND(WX3325, I10470)
--	I10472 = NAND(I10462, I10470)
--	I10461 = NAND(I10471, I10472)
--	I10478 = NAND(WX3389, WX3453)
--	I10479 = NAND(WX3389, I10478)
--	I10480 = NAND(WX3453, I10478)
--	I10477 = NAND(I10479, I10480)
--	I10485 = NAND(I10461, I10477)
--	I10486 = NAND(I10461, I10485)
--	I10487 = NAND(I10477, I10485)
--	WX3501 = NAND(I10486, I10487)
--	I10494 = NAND(WX3588, WX3263)
--	I10495 = NAND(WX3588, I10494)
--	I10496 = NAND(WX3263, I10494)
--	I10493 = NAND(I10495, I10496)
--	I10501 = NAND(WX3327, I10493)
--	I10502 = NAND(WX3327, I10501)
--	I10503 = NAND(I10493, I10501)
--	I10492 = NAND(I10502, I10503)
--	I10509 = NAND(WX3391, WX3455)
--	I10510 = NAND(WX3391, I10509)
--	I10511 = NAND(WX3455, I10509)
--	I10508 = NAND(I10510, I10511)
--	I10516 = NAND(I10492, I10508)
--	I10517 = NAND(I10492, I10516)
--	I10518 = NAND(I10508, I10516)
--	WX3502 = NAND(I10517, I10518)
--	I10525 = NAND(WX3588, WX3265)
--	I10526 = NAND(WX3588, I10525)
--	I10527 = NAND(WX3265, I10525)
--	I10524 = NAND(I10526, I10527)
--	I10532 = NAND(WX3329, I10524)
--	I10533 = NAND(WX3329, I10532)
--	I10534 = NAND(I10524, I10532)
--	I10523 = NAND(I10533, I10534)
--	I10540 = NAND(WX3393, WX3457)
--	I10541 = NAND(WX3393, I10540)
--	I10542 = NAND(WX3457, I10540)
--	I10539 = NAND(I10541, I10542)
--	I10547 = NAND(I10523, I10539)
--	I10548 = NAND(I10523, I10547)
--	I10549 = NAND(I10539, I10547)
--	WX3503 = NAND(I10548, I10549)
--	I10556 = NAND(WX3588, WX3267)
--	I10557 = NAND(WX3588, I10556)
--	I10558 = NAND(WX3267, I10556)
--	I10555 = NAND(I10557, I10558)
--	I10563 = NAND(WX3331, I10555)
--	I10564 = NAND(WX3331, I10563)
--	I10565 = NAND(I10555, I10563)
--	I10554 = NAND(I10564, I10565)
--	I10571 = NAND(WX3395, WX3459)
--	I10572 = NAND(WX3395, I10571)
--	I10573 = NAND(WX3459, I10571)
--	I10570 = NAND(I10572, I10573)
--	I10578 = NAND(I10554, I10570)
--	I10579 = NAND(I10554, I10578)
--	I10580 = NAND(I10570, I10578)
--	WX3504 = NAND(I10579, I10580)
--	I10587 = NAND(WX3588, WX3269)
--	I10588 = NAND(WX3588, I10587)
--	I10589 = NAND(WX3269, I10587)
--	I10586 = NAND(I10588, I10589)
--	I10594 = NAND(WX3333, I10586)
--	I10595 = NAND(WX3333, I10594)
--	I10596 = NAND(I10586, I10594)
--	I10585 = NAND(I10595, I10596)
--	I10602 = NAND(WX3397, WX3461)
--	I10603 = NAND(WX3397, I10602)
--	I10604 = NAND(WX3461, I10602)
--	I10601 = NAND(I10603, I10604)
--	I10609 = NAND(I10585, I10601)
--	I10610 = NAND(I10585, I10609)
--	I10611 = NAND(I10601, I10609)
--	WX3505 = NAND(I10610, I10611)
--	I10618 = NAND(WX3588, WX3271)
--	I10619 = NAND(WX3588, I10618)
--	I10620 = NAND(WX3271, I10618)
--	I10617 = NAND(I10619, I10620)
--	I10625 = NAND(WX3335, I10617)
--	I10626 = NAND(WX3335, I10625)
--	I10627 = NAND(I10617, I10625)
--	I10616 = NAND(I10626, I10627)
--	I10633 = NAND(WX3399, WX3463)
--	I10634 = NAND(WX3399, I10633)
--	I10635 = NAND(WX3463, I10633)
--	I10632 = NAND(I10634, I10635)
--	I10640 = NAND(I10616, I10632)
--	I10641 = NAND(I10616, I10640)
--	I10642 = NAND(I10632, I10640)
--	WX3506 = NAND(I10641, I10642)
--	I10649 = NAND(WX3588, WX3273)
--	I10650 = NAND(WX3588, I10649)
--	I10651 = NAND(WX3273, I10649)
--	I10648 = NAND(I10650, I10651)
--	I10656 = NAND(WX3337, I10648)
--	I10657 = NAND(WX3337, I10656)
--	I10658 = NAND(I10648, I10656)
--	I10647 = NAND(I10657, I10658)
--	I10664 = NAND(WX3401, WX3465)
--	I10665 = NAND(WX3401, I10664)
--	I10666 = NAND(WX3465, I10664)
--	I10663 = NAND(I10665, I10666)
--	I10671 = NAND(I10647, I10663)
--	I10672 = NAND(I10647, I10671)
--	I10673 = NAND(I10663, I10671)
--	WX3507 = NAND(I10672, I10673)
--	I10680 = NAND(WX3588, WX3275)
--	I10681 = NAND(WX3588, I10680)
--	I10682 = NAND(WX3275, I10680)
--	I10679 = NAND(I10681, I10682)
--	I10687 = NAND(WX3339, I10679)
--	I10688 = NAND(WX3339, I10687)
--	I10689 = NAND(I10679, I10687)
--	I10678 = NAND(I10688, I10689)
--	I10695 = NAND(WX3403, WX3467)
--	I10696 = NAND(WX3403, I10695)
--	I10697 = NAND(WX3467, I10695)
--	I10694 = NAND(I10696, I10697)
--	I10702 = NAND(I10678, I10694)
--	I10703 = NAND(I10678, I10702)
--	I10704 = NAND(I10694, I10702)
--	WX3508 = NAND(I10703, I10704)
--	I10711 = NAND(WX3588, WX3277)
--	I10712 = NAND(WX3588, I10711)
--	I10713 = NAND(WX3277, I10711)
--	I10710 = NAND(I10712, I10713)
--	I10718 = NAND(WX3341, I10710)
--	I10719 = NAND(WX3341, I10718)
--	I10720 = NAND(I10710, I10718)
--	I10709 = NAND(I10719, I10720)
--	I10726 = NAND(WX3405, WX3469)
--	I10727 = NAND(WX3405, I10726)
--	I10728 = NAND(WX3469, I10726)
--	I10725 = NAND(I10727, I10728)
--	I10733 = NAND(I10709, I10725)
--	I10734 = NAND(I10709, I10733)
--	I10735 = NAND(I10725, I10733)
--	WX3509 = NAND(I10734, I10735)
--	I10742 = NAND(WX3588, WX3279)
--	I10743 = NAND(WX3588, I10742)
--	I10744 = NAND(WX3279, I10742)
--	I10741 = NAND(I10743, I10744)
--	I10749 = NAND(WX3343, I10741)
--	I10750 = NAND(WX3343, I10749)
--	I10751 = NAND(I10741, I10749)
--	I10740 = NAND(I10750, I10751)
--	I10757 = NAND(WX3407, WX3471)
--	I10758 = NAND(WX3407, I10757)
--	I10759 = NAND(WX3471, I10757)
--	I10756 = NAND(I10758, I10759)
--	I10764 = NAND(I10740, I10756)
--	I10765 = NAND(I10740, I10764)
--	I10766 = NAND(I10756, I10764)
--	WX3510 = NAND(I10765, I10766)
--	I10773 = NAND(WX3588, WX3281)
--	I10774 = NAND(WX3588, I10773)
--	I10775 = NAND(WX3281, I10773)
--	I10772 = NAND(I10774, I10775)
--	I10780 = NAND(WX3345, I10772)
--	I10781 = NAND(WX3345, I10780)
--	I10782 = NAND(I10772, I10780)
--	I10771 = NAND(I10781, I10782)
--	I10788 = NAND(WX3409, WX3473)
--	I10789 = NAND(WX3409, I10788)
--	I10790 = NAND(WX3473, I10788)
--	I10787 = NAND(I10789, I10790)
--	I10795 = NAND(I10771, I10787)
--	I10796 = NAND(I10771, I10795)
--	I10797 = NAND(I10787, I10795)
--	WX3511 = NAND(I10796, I10797)
--	I10804 = NAND(WX3588, WX3283)
--	I10805 = NAND(WX3588, I10804)
--	I10806 = NAND(WX3283, I10804)
--	I10803 = NAND(I10805, I10806)
--	I10811 = NAND(WX3347, I10803)
--	I10812 = NAND(WX3347, I10811)
--	I10813 = NAND(I10803, I10811)
--	I10802 = NAND(I10812, I10813)
--	I10819 = NAND(WX3411, WX3475)
--	I10820 = NAND(WX3411, I10819)
--	I10821 = NAND(WX3475, I10819)
--	I10818 = NAND(I10820, I10821)
--	I10826 = NAND(I10802, I10818)
--	I10827 = NAND(I10802, I10826)
--	I10828 = NAND(I10818, I10826)
--	WX3512 = NAND(I10827, I10828)
--	I10835 = NAND(WX3588, WX3285)
--	I10836 = NAND(WX3588, I10835)
--	I10837 = NAND(WX3285, I10835)
--	I10834 = NAND(I10836, I10837)
--	I10842 = NAND(WX3349, I10834)
--	I10843 = NAND(WX3349, I10842)
--	I10844 = NAND(I10834, I10842)
--	I10833 = NAND(I10843, I10844)
--	I10850 = NAND(WX3413, WX3477)
--	I10851 = NAND(WX3413, I10850)
--	I10852 = NAND(WX3477, I10850)
--	I10849 = NAND(I10851, I10852)
--	I10857 = NAND(I10833, I10849)
--	I10858 = NAND(I10833, I10857)
--	I10859 = NAND(I10849, I10857)
--	WX3513 = NAND(I10858, I10859)
--	I10866 = NAND(WX3588, WX3287)
--	I10867 = NAND(WX3588, I10866)
--	I10868 = NAND(WX3287, I10866)
--	I10865 = NAND(I10867, I10868)
--	I10873 = NAND(WX3351, I10865)
--	I10874 = NAND(WX3351, I10873)
--	I10875 = NAND(I10865, I10873)
--	I10864 = NAND(I10874, I10875)
--	I10881 = NAND(WX3415, WX3479)
--	I10882 = NAND(WX3415, I10881)
--	I10883 = NAND(WX3479, I10881)
--	I10880 = NAND(I10882, I10883)
--	I10888 = NAND(I10864, I10880)
--	I10889 = NAND(I10864, I10888)
--	I10890 = NAND(I10880, I10888)
--	WX3514 = NAND(I10889, I10890)
--	I10897 = NAND(WX3588, WX3289)
--	I10898 = NAND(WX3588, I10897)
--	I10899 = NAND(WX3289, I10897)
--	I10896 = NAND(I10898, I10899)
--	I10904 = NAND(WX3353, I10896)
--	I10905 = NAND(WX3353, I10904)
--	I10906 = NAND(I10896, I10904)
--	I10895 = NAND(I10905, I10906)
--	I10912 = NAND(WX3417, WX3481)
--	I10913 = NAND(WX3417, I10912)
--	I10914 = NAND(WX3481, I10912)
--	I10911 = NAND(I10913, I10914)
--	I10919 = NAND(I10895, I10911)
--	I10920 = NAND(I10895, I10919)
--	I10921 = NAND(I10911, I10919)
--	WX3515 = NAND(I10920, I10921)
--	I10928 = NAND(WX3588, WX3291)
--	I10929 = NAND(WX3588, I10928)
--	I10930 = NAND(WX3291, I10928)
--	I10927 = NAND(I10929, I10930)
--	I10935 = NAND(WX3355, I10927)
--	I10936 = NAND(WX3355, I10935)
--	I10937 = NAND(I10927, I10935)
--	I10926 = NAND(I10936, I10937)
--	I10943 = NAND(WX3419, WX3483)
--	I10944 = NAND(WX3419, I10943)
--	I10945 = NAND(WX3483, I10943)
--	I10942 = NAND(I10944, I10945)
--	I10950 = NAND(I10926, I10942)
--	I10951 = NAND(I10926, I10950)
--	I10952 = NAND(I10942, I10950)
--	WX3516 = NAND(I10951, I10952)
--	I10959 = NAND(WX3588, WX3293)
--	I10960 = NAND(WX3588, I10959)
--	I10961 = NAND(WX3293, I10959)
--	I10958 = NAND(I10960, I10961)
--	I10966 = NAND(WX3357, I10958)
--	I10967 = NAND(WX3357, I10966)
--	I10968 = NAND(I10958, I10966)
--	I10957 = NAND(I10967, I10968)
--	I10974 = NAND(WX3421, WX3485)
--	I10975 = NAND(WX3421, I10974)
--	I10976 = NAND(WX3485, I10974)
--	I10973 = NAND(I10975, I10976)
--	I10981 = NAND(I10957, I10973)
--	I10982 = NAND(I10957, I10981)
--	I10983 = NAND(I10973, I10981)
--	WX3517 = NAND(I10982, I10983)
--	I11062 = NAND(WX3166, WX3071)
--	I11063 = NAND(WX3166, I11062)
--	I11064 = NAND(WX3071, I11062)
--	WX3592 = NAND(I11063, I11064)
--	I11075 = NAND(WX3167, WX3073)
--	I11076 = NAND(WX3167, I11075)
--	I11077 = NAND(WX3073, I11075)
--	WX3599 = NAND(I11076, I11077)
--	I11088 = NAND(WX3168, WX3075)
--	I11089 = NAND(WX3168, I11088)
--	I11090 = NAND(WX3075, I11088)
--	WX3606 = NAND(I11089, I11090)
--	I11101 = NAND(WX3169, WX3077)
--	I11102 = NAND(WX3169, I11101)
--	I11103 = NAND(WX3077, I11101)
--	WX3613 = NAND(I11102, I11103)
--	I11114 = NAND(WX3170, WX3079)
--	I11115 = NAND(WX3170, I11114)
--	I11116 = NAND(WX3079, I11114)
--	WX3620 = NAND(I11115, I11116)
--	I11127 = NAND(WX3171, WX3081)
--	I11128 = NAND(WX3171, I11127)
--	I11129 = NAND(WX3081, I11127)
--	WX3627 = NAND(I11128, I11129)
--	I11140 = NAND(WX3172, WX3083)
--	I11141 = NAND(WX3172, I11140)
--	I11142 = NAND(WX3083, I11140)
--	WX3634 = NAND(I11141, I11142)
--	I11153 = NAND(WX3173, WX3085)
--	I11154 = NAND(WX3173, I11153)
--	I11155 = NAND(WX3085, I11153)
--	WX3641 = NAND(I11154, I11155)
--	I11166 = NAND(WX3174, WX3087)
--	I11167 = NAND(WX3174, I11166)
--	I11168 = NAND(WX3087, I11166)
--	WX3648 = NAND(I11167, I11168)
--	I11179 = NAND(WX3175, WX3089)
--	I11180 = NAND(WX3175, I11179)
--	I11181 = NAND(WX3089, I11179)
--	WX3655 = NAND(I11180, I11181)
--	I11192 = NAND(WX3176, WX3091)
--	I11193 = NAND(WX3176, I11192)
--	I11194 = NAND(WX3091, I11192)
--	WX3662 = NAND(I11193, I11194)
--	I11205 = NAND(WX3177, WX3093)
--	I11206 = NAND(WX3177, I11205)
--	I11207 = NAND(WX3093, I11205)
--	WX3669 = NAND(I11206, I11207)
--	I11218 = NAND(WX3178, WX3095)
--	I11219 = NAND(WX3178, I11218)
--	I11220 = NAND(WX3095, I11218)
--	WX3676 = NAND(I11219, I11220)
--	I11231 = NAND(WX3179, WX3097)
--	I11232 = NAND(WX3179, I11231)
--	I11233 = NAND(WX3097, I11231)
--	WX3683 = NAND(I11232, I11233)
--	I11244 = NAND(WX3180, WX3099)
--	I11245 = NAND(WX3180, I11244)
--	I11246 = NAND(WX3099, I11244)
--	WX3690 = NAND(I11245, I11246)
--	I11257 = NAND(WX3181, WX3101)
--	I11258 = NAND(WX3181, I11257)
--	I11259 = NAND(WX3101, I11257)
--	WX3697 = NAND(I11258, I11259)
--	I11270 = NAND(WX3182, WX3103)
--	I11271 = NAND(WX3182, I11270)
--	I11272 = NAND(WX3103, I11270)
--	WX3704 = NAND(I11271, I11272)
--	I11283 = NAND(WX3183, WX3105)
--	I11284 = NAND(WX3183, I11283)
--	I11285 = NAND(WX3105, I11283)
--	WX3711 = NAND(I11284, I11285)
--	I11296 = NAND(WX3184, WX3107)
--	I11297 = NAND(WX3184, I11296)
--	I11298 = NAND(WX3107, I11296)
--	WX3718 = NAND(I11297, I11298)
--	I11309 = NAND(WX3185, WX3109)
--	I11310 = NAND(WX3185, I11309)
--	I11311 = NAND(WX3109, I11309)
--	WX3725 = NAND(I11310, I11311)
--	I11322 = NAND(WX3186, WX3111)
--	I11323 = NAND(WX3186, I11322)
--	I11324 = NAND(WX3111, I11322)
--	WX3732 = NAND(I11323, I11324)
--	I11335 = NAND(WX3187, WX3113)
--	I11336 = NAND(WX3187, I11335)
--	I11337 = NAND(WX3113, I11335)
--	WX3739 = NAND(I11336, I11337)
--	I11348 = NAND(WX3188, WX3115)
--	I11349 = NAND(WX3188, I11348)
--	I11350 = NAND(WX3115, I11348)
--	WX3746 = NAND(I11349, I11350)
--	I11361 = NAND(WX3189, WX3117)
--	I11362 = NAND(WX3189, I11361)
--	I11363 = NAND(WX3117, I11361)
--	WX3753 = NAND(I11362, I11363)
--	I11374 = NAND(WX3190, WX3119)
--	I11375 = NAND(WX3190, I11374)
--	I11376 = NAND(WX3119, I11374)
--	WX3760 = NAND(I11375, I11376)
--	I11387 = NAND(WX3191, WX3121)
--	I11388 = NAND(WX3191, I11387)
--	I11389 = NAND(WX3121, I11387)
--	WX3767 = NAND(I11388, I11389)
--	I11400 = NAND(WX3192, WX3123)
--	I11401 = NAND(WX3192, I11400)
--	I11402 = NAND(WX3123, I11400)
--	WX3774 = NAND(I11401, I11402)
--	I11413 = NAND(WX3193, WX3125)
--	I11414 = NAND(WX3193, I11413)
--	I11415 = NAND(WX3125, I11413)
--	WX3781 = NAND(I11414, I11415)
--	I11426 = NAND(WX3194, WX3127)
--	I11427 = NAND(WX3194, I11426)
--	I11428 = NAND(WX3127, I11426)
--	WX3788 = NAND(I11427, I11428)
--	I11439 = NAND(WX3195, WX3129)
--	I11440 = NAND(WX3195, I11439)
--	I11441 = NAND(WX3129, I11439)
--	WX3795 = NAND(I11440, I11441)
--	I11452 = NAND(WX3196, WX3131)
--	I11453 = NAND(WX3196, I11452)
--	I11454 = NAND(WX3131, I11452)
--	WX3802 = NAND(I11453, I11454)
--	I11465 = NAND(WX3197, WX3133)
--	I11466 = NAND(WX3197, I11465)
--	I11467 = NAND(WX3133, I11465)
--	WX3809 = NAND(I11466, I11467)
--	I11480 = NAND(WX3213, CRC_OUT_7_31)
--	I11481 = NAND(WX3213, I11480)
--	I11482 = NAND(CRC_OUT_7_31, I11480)
--	I11479 = NAND(I11481, I11482)
--	I11487 = NAND(CRC_OUT_7_15, I11479)
--	I11488 = NAND(CRC_OUT_7_15, I11487)
--	I11489 = NAND(I11479, I11487)
--	WX3817 = NAND(I11488, I11489)
--	I11495 = NAND(WX3218, CRC_OUT_7_31)
--	I11496 = NAND(WX3218, I11495)
--	I11497 = NAND(CRC_OUT_7_31, I11495)
--	I11494 = NAND(I11496, I11497)
--	I11502 = NAND(CRC_OUT_7_10, I11494)
--	I11503 = NAND(CRC_OUT_7_10, I11502)
--	I11504 = NAND(I11494, I11502)
--	WX3818 = NAND(I11503, I11504)
--	I11510 = NAND(WX3225, CRC_OUT_7_31)
--	I11511 = NAND(WX3225, I11510)
--	I11512 = NAND(CRC_OUT_7_31, I11510)
--	I11509 = NAND(I11511, I11512)
--	I11517 = NAND(CRC_OUT_7_3, I11509)
--	I11518 = NAND(CRC_OUT_7_3, I11517)
--	I11519 = NAND(I11509, I11517)
--	WX3819 = NAND(I11518, I11519)
--	I11524 = NAND(WX3229, CRC_OUT_7_31)
--	I11525 = NAND(WX3229, I11524)
--	I11526 = NAND(CRC_OUT_7_31, I11524)
--	WX3820 = NAND(I11525, I11526)
--	I11531 = NAND(WX3198, CRC_OUT_7_30)
--	I11532 = NAND(WX3198, I11531)
--	I11533 = NAND(CRC_OUT_7_30, I11531)
--	WX3821 = NAND(I11532, I11533)
--	I11538 = NAND(WX3199, CRC_OUT_7_29)
--	I11539 = NAND(WX3199, I11538)
--	I11540 = NAND(CRC_OUT_7_29, I11538)
--	WX3822 = NAND(I11539, I11540)
--	I11545 = NAND(WX3200, CRC_OUT_7_28)
--	I11546 = NAND(WX3200, I11545)
--	I11547 = NAND(CRC_OUT_7_28, I11545)
--	WX3823 = NAND(I11546, I11547)
--	I11552 = NAND(WX3201, CRC_OUT_7_27)
--	I11553 = NAND(WX3201, I11552)
--	I11554 = NAND(CRC_OUT_7_27, I11552)
--	WX3824 = NAND(I11553, I11554)
--	I11559 = NAND(WX3202, CRC_OUT_7_26)
--	I11560 = NAND(WX3202, I11559)
--	I11561 = NAND(CRC_OUT_7_26, I11559)
--	WX3825 = NAND(I11560, I11561)
--	I11566 = NAND(WX3203, CRC_OUT_7_25)
--	I11567 = NAND(WX3203, I11566)
--	I11568 = NAND(CRC_OUT_7_25, I11566)
--	WX3826 = NAND(I11567, I11568)
--	I11573 = NAND(WX3204, CRC_OUT_7_24)
--	I11574 = NAND(WX3204, I11573)
--	I11575 = NAND(CRC_OUT_7_24, I11573)
--	WX3827 = NAND(I11574, I11575)
--	I11580 = NAND(WX3205, CRC_OUT_7_23)
--	I11581 = NAND(WX3205, I11580)
--	I11582 = NAND(CRC_OUT_7_23, I11580)
--	WX3828 = NAND(I11581, I11582)
--	I11587 = NAND(WX3206, CRC_OUT_7_22)
--	I11588 = NAND(WX3206, I11587)
--	I11589 = NAND(CRC_OUT_7_22, I11587)
--	WX3829 = NAND(I11588, I11589)
--	I11594 = NAND(WX3207, CRC_OUT_7_21)
--	I11595 = NAND(WX3207, I11594)
--	I11596 = NAND(CRC_OUT_7_21, I11594)
--	WX3830 = NAND(I11595, I11596)
--	I11601 = NAND(WX3208, CRC_OUT_7_20)
--	I11602 = NAND(WX3208, I11601)
--	I11603 = NAND(CRC_OUT_7_20, I11601)
--	WX3831 = NAND(I11602, I11603)
--	I11608 = NAND(WX3209, CRC_OUT_7_19)
--	I11609 = NAND(WX3209, I11608)
--	I11610 = NAND(CRC_OUT_7_19, I11608)
--	WX3832 = NAND(I11609, I11610)
--	I11615 = NAND(WX3210, CRC_OUT_7_18)
--	I11616 = NAND(WX3210, I11615)
--	I11617 = NAND(CRC_OUT_7_18, I11615)
--	WX3833 = NAND(I11616, I11617)
--	I11622 = NAND(WX3211, CRC_OUT_7_17)
--	I11623 = NAND(WX3211, I11622)
--	I11624 = NAND(CRC_OUT_7_17, I11622)
--	WX3834 = NAND(I11623, I11624)
--	I11629 = NAND(WX3212, CRC_OUT_7_16)
--	I11630 = NAND(WX3212, I11629)
--	I11631 = NAND(CRC_OUT_7_16, I11629)
--	WX3835 = NAND(I11630, I11631)
--	I11636 = NAND(WX3214, CRC_OUT_7_14)
--	I11637 = NAND(WX3214, I11636)
--	I11638 = NAND(CRC_OUT_7_14, I11636)
--	WX3836 = NAND(I11637, I11638)
--	I11643 = NAND(WX3215, CRC_OUT_7_13)
--	I11644 = NAND(WX3215, I11643)
--	I11645 = NAND(CRC_OUT_7_13, I11643)
--	WX3837 = NAND(I11644, I11645)
--	I11650 = NAND(WX3216, CRC_OUT_7_12)
--	I11651 = NAND(WX3216, I11650)
--	I11652 = NAND(CRC_OUT_7_12, I11650)
--	WX3838 = NAND(I11651, I11652)
--	I11657 = NAND(WX3217, CRC_OUT_7_11)
--	I11658 = NAND(WX3217, I11657)
--	I11659 = NAND(CRC_OUT_7_11, I11657)
--	WX3839 = NAND(I11658, I11659)
--	I11664 = NAND(WX3219, CRC_OUT_7_9)
--	I11665 = NAND(WX3219, I11664)
--	I11666 = NAND(CRC_OUT_7_9, I11664)
--	WX3840 = NAND(I11665, I11666)
--	I11671 = NAND(WX3220, CRC_OUT_7_8)
--	I11672 = NAND(WX3220, I11671)
--	I11673 = NAND(CRC_OUT_7_8, I11671)
--	WX3841 = NAND(I11672, I11673)
--	I11678 = NAND(WX3221, CRC_OUT_7_7)
--	I11679 = NAND(WX3221, I11678)
--	I11680 = NAND(CRC_OUT_7_7, I11678)
--	WX3842 = NAND(I11679, I11680)
--	I11685 = NAND(WX3222, CRC_OUT_7_6)
--	I11686 = NAND(WX3222, I11685)
--	I11687 = NAND(CRC_OUT_7_6, I11685)
--	WX3843 = NAND(I11686, I11687)
--	I11692 = NAND(WX3223, CRC_OUT_7_5)
--	I11693 = NAND(WX3223, I11692)
--	I11694 = NAND(CRC_OUT_7_5, I11692)
--	WX3844 = NAND(I11693, I11694)
--	I11699 = NAND(WX3224, CRC_OUT_7_4)
--	I11700 = NAND(WX3224, I11699)
--	I11701 = NAND(CRC_OUT_7_4, I11699)
--	WX3845 = NAND(I11700, I11701)
--	I11706 = NAND(WX3226, CRC_OUT_7_2)
--	I11707 = NAND(WX3226, I11706)
--	I11708 = NAND(CRC_OUT_7_2, I11706)
--	WX3846 = NAND(I11707, I11708)
--	I11713 = NAND(WX3227, CRC_OUT_7_1)
--	I11714 = NAND(WX3227, I11713)
--	I11715 = NAND(CRC_OUT_7_1, I11713)
--	WX3847 = NAND(I11714, I11715)
--	I11720 = NAND(WX3228, CRC_OUT_7_0)
--	I11721 = NAND(WX3228, I11720)
--	I11722 = NAND(CRC_OUT_7_0, I11720)
--	WX3848 = NAND(I11721, I11722)
--	I14003 = NAND(WX4880, WX4524)
--	I14004 = NAND(WX4880, I14003)
--	I14005 = NAND(WX4524, I14003)
--	I14002 = NAND(I14004, I14005)
--	I14010 = NAND(WX4588, I14002)
--	I14011 = NAND(WX4588, I14010)
--	I14012 = NAND(I14002, I14010)
--	I14001 = NAND(I14011, I14012)
--	I14018 = NAND(WX4652, WX4716)
--	I14019 = NAND(WX4652, I14018)
--	I14020 = NAND(WX4716, I14018)
--	I14017 = NAND(I14019, I14020)
--	I14025 = NAND(I14001, I14017)
--	I14026 = NAND(I14001, I14025)
--	I14027 = NAND(I14017, I14025)
--	WX4779 = NAND(I14026, I14027)
--	I14034 = NAND(WX4880, WX4526)
--	I14035 = NAND(WX4880, I14034)
--	I14036 = NAND(WX4526, I14034)
--	I14033 = NAND(I14035, I14036)
--	I14041 = NAND(WX4590, I14033)
--	I14042 = NAND(WX4590, I14041)
--	I14043 = NAND(I14033, I14041)
--	I14032 = NAND(I14042, I14043)
--	I14049 = NAND(WX4654, WX4718)
--	I14050 = NAND(WX4654, I14049)
--	I14051 = NAND(WX4718, I14049)
--	I14048 = NAND(I14050, I14051)
--	I14056 = NAND(I14032, I14048)
--	I14057 = NAND(I14032, I14056)
--	I14058 = NAND(I14048, I14056)
--	WX4780 = NAND(I14057, I14058)
--	I14065 = NAND(WX4880, WX4528)
--	I14066 = NAND(WX4880, I14065)
--	I14067 = NAND(WX4528, I14065)
--	I14064 = NAND(I14066, I14067)
--	I14072 = NAND(WX4592, I14064)
--	I14073 = NAND(WX4592, I14072)
--	I14074 = NAND(I14064, I14072)
--	I14063 = NAND(I14073, I14074)
--	I14080 = NAND(WX4656, WX4720)
--	I14081 = NAND(WX4656, I14080)
--	I14082 = NAND(WX4720, I14080)
--	I14079 = NAND(I14081, I14082)
--	I14087 = NAND(I14063, I14079)
--	I14088 = NAND(I14063, I14087)
--	I14089 = NAND(I14079, I14087)
--	WX4781 = NAND(I14088, I14089)
--	I14096 = NAND(WX4880, WX4530)
--	I14097 = NAND(WX4880, I14096)
--	I14098 = NAND(WX4530, I14096)
--	I14095 = NAND(I14097, I14098)
--	I14103 = NAND(WX4594, I14095)
--	I14104 = NAND(WX4594, I14103)
--	I14105 = NAND(I14095, I14103)
--	I14094 = NAND(I14104, I14105)
--	I14111 = NAND(WX4658, WX4722)
--	I14112 = NAND(WX4658, I14111)
--	I14113 = NAND(WX4722, I14111)
--	I14110 = NAND(I14112, I14113)
--	I14118 = NAND(I14094, I14110)
--	I14119 = NAND(I14094, I14118)
--	I14120 = NAND(I14110, I14118)
--	WX4782 = NAND(I14119, I14120)
--	I14127 = NAND(WX4880, WX4532)
--	I14128 = NAND(WX4880, I14127)
--	I14129 = NAND(WX4532, I14127)
--	I14126 = NAND(I14128, I14129)
--	I14134 = NAND(WX4596, I14126)
--	I14135 = NAND(WX4596, I14134)
--	I14136 = NAND(I14126, I14134)
--	I14125 = NAND(I14135, I14136)
--	I14142 = NAND(WX4660, WX4724)
--	I14143 = NAND(WX4660, I14142)
--	I14144 = NAND(WX4724, I14142)
--	I14141 = NAND(I14143, I14144)
--	I14149 = NAND(I14125, I14141)
--	I14150 = NAND(I14125, I14149)
--	I14151 = NAND(I14141, I14149)
--	WX4783 = NAND(I14150, I14151)
--	I14158 = NAND(WX4880, WX4534)
--	I14159 = NAND(WX4880, I14158)
--	I14160 = NAND(WX4534, I14158)
--	I14157 = NAND(I14159, I14160)
--	I14165 = NAND(WX4598, I14157)
--	I14166 = NAND(WX4598, I14165)
--	I14167 = NAND(I14157, I14165)
--	I14156 = NAND(I14166, I14167)
--	I14173 = NAND(WX4662, WX4726)
--	I14174 = NAND(WX4662, I14173)
--	I14175 = NAND(WX4726, I14173)
--	I14172 = NAND(I14174, I14175)
--	I14180 = NAND(I14156, I14172)
--	I14181 = NAND(I14156, I14180)
--	I14182 = NAND(I14172, I14180)
--	WX4784 = NAND(I14181, I14182)
--	I14189 = NAND(WX4880, WX4536)
--	I14190 = NAND(WX4880, I14189)
--	I14191 = NAND(WX4536, I14189)
--	I14188 = NAND(I14190, I14191)
--	I14196 = NAND(WX4600, I14188)
--	I14197 = NAND(WX4600, I14196)
--	I14198 = NAND(I14188, I14196)
--	I14187 = NAND(I14197, I14198)
--	I14204 = NAND(WX4664, WX4728)
--	I14205 = NAND(WX4664, I14204)
--	I14206 = NAND(WX4728, I14204)
--	I14203 = NAND(I14205, I14206)
--	I14211 = NAND(I14187, I14203)
--	I14212 = NAND(I14187, I14211)
--	I14213 = NAND(I14203, I14211)
--	WX4785 = NAND(I14212, I14213)
--	I14220 = NAND(WX4880, WX4538)
--	I14221 = NAND(WX4880, I14220)
--	I14222 = NAND(WX4538, I14220)
--	I14219 = NAND(I14221, I14222)
--	I14227 = NAND(WX4602, I14219)
--	I14228 = NAND(WX4602, I14227)
--	I14229 = NAND(I14219, I14227)
--	I14218 = NAND(I14228, I14229)
--	I14235 = NAND(WX4666, WX4730)
--	I14236 = NAND(WX4666, I14235)
--	I14237 = NAND(WX4730, I14235)
--	I14234 = NAND(I14236, I14237)
--	I14242 = NAND(I14218, I14234)
--	I14243 = NAND(I14218, I14242)
--	I14244 = NAND(I14234, I14242)
--	WX4786 = NAND(I14243, I14244)
--	I14251 = NAND(WX4880, WX4540)
--	I14252 = NAND(WX4880, I14251)
--	I14253 = NAND(WX4540, I14251)
--	I14250 = NAND(I14252, I14253)
--	I14258 = NAND(WX4604, I14250)
--	I14259 = NAND(WX4604, I14258)
--	I14260 = NAND(I14250, I14258)
--	I14249 = NAND(I14259, I14260)
--	I14266 = NAND(WX4668, WX4732)
--	I14267 = NAND(WX4668, I14266)
--	I14268 = NAND(WX4732, I14266)
--	I14265 = NAND(I14267, I14268)
--	I14273 = NAND(I14249, I14265)
--	I14274 = NAND(I14249, I14273)
--	I14275 = NAND(I14265, I14273)
--	WX4787 = NAND(I14274, I14275)
--	I14282 = NAND(WX4880, WX4542)
--	I14283 = NAND(WX4880, I14282)
--	I14284 = NAND(WX4542, I14282)
--	I14281 = NAND(I14283, I14284)
--	I14289 = NAND(WX4606, I14281)
--	I14290 = NAND(WX4606, I14289)
--	I14291 = NAND(I14281, I14289)
--	I14280 = NAND(I14290, I14291)
--	I14297 = NAND(WX4670, WX4734)
--	I14298 = NAND(WX4670, I14297)
--	I14299 = NAND(WX4734, I14297)
--	I14296 = NAND(I14298, I14299)
--	I14304 = NAND(I14280, I14296)
--	I14305 = NAND(I14280, I14304)
--	I14306 = NAND(I14296, I14304)
--	WX4788 = NAND(I14305, I14306)
--	I14313 = NAND(WX4880, WX4544)
--	I14314 = NAND(WX4880, I14313)
--	I14315 = NAND(WX4544, I14313)
--	I14312 = NAND(I14314, I14315)
--	I14320 = NAND(WX4608, I14312)
--	I14321 = NAND(WX4608, I14320)
--	I14322 = NAND(I14312, I14320)
--	I14311 = NAND(I14321, I14322)
--	I14328 = NAND(WX4672, WX4736)
--	I14329 = NAND(WX4672, I14328)
--	I14330 = NAND(WX4736, I14328)
--	I14327 = NAND(I14329, I14330)
--	I14335 = NAND(I14311, I14327)
--	I14336 = NAND(I14311, I14335)
--	I14337 = NAND(I14327, I14335)
--	WX4789 = NAND(I14336, I14337)
--	I14344 = NAND(WX4880, WX4546)
--	I14345 = NAND(WX4880, I14344)
--	I14346 = NAND(WX4546, I14344)
--	I14343 = NAND(I14345, I14346)
--	I14351 = NAND(WX4610, I14343)
--	I14352 = NAND(WX4610, I14351)
--	I14353 = NAND(I14343, I14351)
--	I14342 = NAND(I14352, I14353)
--	I14359 = NAND(WX4674, WX4738)
--	I14360 = NAND(WX4674, I14359)
--	I14361 = NAND(WX4738, I14359)
--	I14358 = NAND(I14360, I14361)
--	I14366 = NAND(I14342, I14358)
--	I14367 = NAND(I14342, I14366)
--	I14368 = NAND(I14358, I14366)
--	WX4790 = NAND(I14367, I14368)
--	I14375 = NAND(WX4880, WX4548)
--	I14376 = NAND(WX4880, I14375)
--	I14377 = NAND(WX4548, I14375)
--	I14374 = NAND(I14376, I14377)
--	I14382 = NAND(WX4612, I14374)
--	I14383 = NAND(WX4612, I14382)
--	I14384 = NAND(I14374, I14382)
--	I14373 = NAND(I14383, I14384)
--	I14390 = NAND(WX4676, WX4740)
--	I14391 = NAND(WX4676, I14390)
--	I14392 = NAND(WX4740, I14390)
--	I14389 = NAND(I14391, I14392)
--	I14397 = NAND(I14373, I14389)
--	I14398 = NAND(I14373, I14397)
--	I14399 = NAND(I14389, I14397)
--	WX4791 = NAND(I14398, I14399)
--	I14406 = NAND(WX4880, WX4550)
--	I14407 = NAND(WX4880, I14406)
--	I14408 = NAND(WX4550, I14406)
--	I14405 = NAND(I14407, I14408)
--	I14413 = NAND(WX4614, I14405)
--	I14414 = NAND(WX4614, I14413)
--	I14415 = NAND(I14405, I14413)
--	I14404 = NAND(I14414, I14415)
--	I14421 = NAND(WX4678, WX4742)
--	I14422 = NAND(WX4678, I14421)
--	I14423 = NAND(WX4742, I14421)
--	I14420 = NAND(I14422, I14423)
--	I14428 = NAND(I14404, I14420)
--	I14429 = NAND(I14404, I14428)
--	I14430 = NAND(I14420, I14428)
--	WX4792 = NAND(I14429, I14430)
--	I14437 = NAND(WX4880, WX4552)
--	I14438 = NAND(WX4880, I14437)
--	I14439 = NAND(WX4552, I14437)
--	I14436 = NAND(I14438, I14439)
--	I14444 = NAND(WX4616, I14436)
--	I14445 = NAND(WX4616, I14444)
--	I14446 = NAND(I14436, I14444)
--	I14435 = NAND(I14445, I14446)
--	I14452 = NAND(WX4680, WX4744)
--	I14453 = NAND(WX4680, I14452)
--	I14454 = NAND(WX4744, I14452)
--	I14451 = NAND(I14453, I14454)
--	I14459 = NAND(I14435, I14451)
--	I14460 = NAND(I14435, I14459)
--	I14461 = NAND(I14451, I14459)
--	WX4793 = NAND(I14460, I14461)
--	I14468 = NAND(WX4880, WX4554)
--	I14469 = NAND(WX4880, I14468)
--	I14470 = NAND(WX4554, I14468)
--	I14467 = NAND(I14469, I14470)
--	I14475 = NAND(WX4618, I14467)
--	I14476 = NAND(WX4618, I14475)
--	I14477 = NAND(I14467, I14475)
--	I14466 = NAND(I14476, I14477)
--	I14483 = NAND(WX4682, WX4746)
--	I14484 = NAND(WX4682, I14483)
--	I14485 = NAND(WX4746, I14483)
--	I14482 = NAND(I14484, I14485)
--	I14490 = NAND(I14466, I14482)
--	I14491 = NAND(I14466, I14490)
--	I14492 = NAND(I14482, I14490)
--	WX4794 = NAND(I14491, I14492)
--	I14499 = NAND(WX4881, WX4556)
--	I14500 = NAND(WX4881, I14499)
--	I14501 = NAND(WX4556, I14499)
--	I14498 = NAND(I14500, I14501)
--	I14506 = NAND(WX4620, I14498)
--	I14507 = NAND(WX4620, I14506)
--	I14508 = NAND(I14498, I14506)
--	I14497 = NAND(I14507, I14508)
--	I14514 = NAND(WX4684, WX4748)
--	I14515 = NAND(WX4684, I14514)
--	I14516 = NAND(WX4748, I14514)
--	I14513 = NAND(I14515, I14516)
--	I14521 = NAND(I14497, I14513)
--	I14522 = NAND(I14497, I14521)
--	I14523 = NAND(I14513, I14521)
--	WX4795 = NAND(I14522, I14523)
--	I14530 = NAND(WX4881, WX4558)
--	I14531 = NAND(WX4881, I14530)
--	I14532 = NAND(WX4558, I14530)
--	I14529 = NAND(I14531, I14532)
--	I14537 = NAND(WX4622, I14529)
--	I14538 = NAND(WX4622, I14537)
--	I14539 = NAND(I14529, I14537)
--	I14528 = NAND(I14538, I14539)
--	I14545 = NAND(WX4686, WX4750)
--	I14546 = NAND(WX4686, I14545)
--	I14547 = NAND(WX4750, I14545)
--	I14544 = NAND(I14546, I14547)
--	I14552 = NAND(I14528, I14544)
--	I14553 = NAND(I14528, I14552)
--	I14554 = NAND(I14544, I14552)
--	WX4796 = NAND(I14553, I14554)
--	I14561 = NAND(WX4881, WX4560)
--	I14562 = NAND(WX4881, I14561)
--	I14563 = NAND(WX4560, I14561)
--	I14560 = NAND(I14562, I14563)
--	I14568 = NAND(WX4624, I14560)
--	I14569 = NAND(WX4624, I14568)
--	I14570 = NAND(I14560, I14568)
--	I14559 = NAND(I14569, I14570)
--	I14576 = NAND(WX4688, WX4752)
--	I14577 = NAND(WX4688, I14576)
--	I14578 = NAND(WX4752, I14576)
--	I14575 = NAND(I14577, I14578)
--	I14583 = NAND(I14559, I14575)
--	I14584 = NAND(I14559, I14583)
--	I14585 = NAND(I14575, I14583)
--	WX4797 = NAND(I14584, I14585)
--	I14592 = NAND(WX4881, WX4562)
--	I14593 = NAND(WX4881, I14592)
--	I14594 = NAND(WX4562, I14592)
--	I14591 = NAND(I14593, I14594)
--	I14599 = NAND(WX4626, I14591)
--	I14600 = NAND(WX4626, I14599)
--	I14601 = NAND(I14591, I14599)
--	I14590 = NAND(I14600, I14601)
--	I14607 = NAND(WX4690, WX4754)
--	I14608 = NAND(WX4690, I14607)
--	I14609 = NAND(WX4754, I14607)
--	I14606 = NAND(I14608, I14609)
--	I14614 = NAND(I14590, I14606)
--	I14615 = NAND(I14590, I14614)
--	I14616 = NAND(I14606, I14614)
--	WX4798 = NAND(I14615, I14616)
--	I14623 = NAND(WX4881, WX4564)
--	I14624 = NAND(WX4881, I14623)
--	I14625 = NAND(WX4564, I14623)
--	I14622 = NAND(I14624, I14625)
--	I14630 = NAND(WX4628, I14622)
--	I14631 = NAND(WX4628, I14630)
--	I14632 = NAND(I14622, I14630)
--	I14621 = NAND(I14631, I14632)
--	I14638 = NAND(WX4692, WX4756)
--	I14639 = NAND(WX4692, I14638)
--	I14640 = NAND(WX4756, I14638)
--	I14637 = NAND(I14639, I14640)
--	I14645 = NAND(I14621, I14637)
--	I14646 = NAND(I14621, I14645)
--	I14647 = NAND(I14637, I14645)
--	WX4799 = NAND(I14646, I14647)
--	I14654 = NAND(WX4881, WX4566)
--	I14655 = NAND(WX4881, I14654)
--	I14656 = NAND(WX4566, I14654)
--	I14653 = NAND(I14655, I14656)
--	I14661 = NAND(WX4630, I14653)
--	I14662 = NAND(WX4630, I14661)
--	I14663 = NAND(I14653, I14661)
--	I14652 = NAND(I14662, I14663)
--	I14669 = NAND(WX4694, WX4758)
--	I14670 = NAND(WX4694, I14669)
--	I14671 = NAND(WX4758, I14669)
--	I14668 = NAND(I14670, I14671)
--	I14676 = NAND(I14652, I14668)
--	I14677 = NAND(I14652, I14676)
--	I14678 = NAND(I14668, I14676)
--	WX4800 = NAND(I14677, I14678)
--	I14685 = NAND(WX4881, WX4568)
--	I14686 = NAND(WX4881, I14685)
--	I14687 = NAND(WX4568, I14685)
--	I14684 = NAND(I14686, I14687)
--	I14692 = NAND(WX4632, I14684)
--	I14693 = NAND(WX4632, I14692)
--	I14694 = NAND(I14684, I14692)
--	I14683 = NAND(I14693, I14694)
--	I14700 = NAND(WX4696, WX4760)
--	I14701 = NAND(WX4696, I14700)
--	I14702 = NAND(WX4760, I14700)
--	I14699 = NAND(I14701, I14702)
--	I14707 = NAND(I14683, I14699)
--	I14708 = NAND(I14683, I14707)
--	I14709 = NAND(I14699, I14707)
--	WX4801 = NAND(I14708, I14709)
--	I14716 = NAND(WX4881, WX4570)
--	I14717 = NAND(WX4881, I14716)
--	I14718 = NAND(WX4570, I14716)
--	I14715 = NAND(I14717, I14718)
--	I14723 = NAND(WX4634, I14715)
--	I14724 = NAND(WX4634, I14723)
--	I14725 = NAND(I14715, I14723)
--	I14714 = NAND(I14724, I14725)
--	I14731 = NAND(WX4698, WX4762)
--	I14732 = NAND(WX4698, I14731)
--	I14733 = NAND(WX4762, I14731)
--	I14730 = NAND(I14732, I14733)
--	I14738 = NAND(I14714, I14730)
--	I14739 = NAND(I14714, I14738)
--	I14740 = NAND(I14730, I14738)
--	WX4802 = NAND(I14739, I14740)
--	I14747 = NAND(WX4881, WX4572)
--	I14748 = NAND(WX4881, I14747)
--	I14749 = NAND(WX4572, I14747)
--	I14746 = NAND(I14748, I14749)
--	I14754 = NAND(WX4636, I14746)
--	I14755 = NAND(WX4636, I14754)
--	I14756 = NAND(I14746, I14754)
--	I14745 = NAND(I14755, I14756)
--	I14762 = NAND(WX4700, WX4764)
--	I14763 = NAND(WX4700, I14762)
--	I14764 = NAND(WX4764, I14762)
--	I14761 = NAND(I14763, I14764)
--	I14769 = NAND(I14745, I14761)
--	I14770 = NAND(I14745, I14769)
--	I14771 = NAND(I14761, I14769)
--	WX4803 = NAND(I14770, I14771)
--	I14778 = NAND(WX4881, WX4574)
--	I14779 = NAND(WX4881, I14778)
--	I14780 = NAND(WX4574, I14778)
--	I14777 = NAND(I14779, I14780)
--	I14785 = NAND(WX4638, I14777)
--	I14786 = NAND(WX4638, I14785)
--	I14787 = NAND(I14777, I14785)
--	I14776 = NAND(I14786, I14787)
--	I14793 = NAND(WX4702, WX4766)
--	I14794 = NAND(WX4702, I14793)
--	I14795 = NAND(WX4766, I14793)
--	I14792 = NAND(I14794, I14795)
--	I14800 = NAND(I14776, I14792)
--	I14801 = NAND(I14776, I14800)
--	I14802 = NAND(I14792, I14800)
--	WX4804 = NAND(I14801, I14802)
--	I14809 = NAND(WX4881, WX4576)
--	I14810 = NAND(WX4881, I14809)
--	I14811 = NAND(WX4576, I14809)
--	I14808 = NAND(I14810, I14811)
--	I14816 = NAND(WX4640, I14808)
--	I14817 = NAND(WX4640, I14816)
--	I14818 = NAND(I14808, I14816)
--	I14807 = NAND(I14817, I14818)
--	I14824 = NAND(WX4704, WX4768)
--	I14825 = NAND(WX4704, I14824)
--	I14826 = NAND(WX4768, I14824)
--	I14823 = NAND(I14825, I14826)
--	I14831 = NAND(I14807, I14823)
--	I14832 = NAND(I14807, I14831)
--	I14833 = NAND(I14823, I14831)
--	WX4805 = NAND(I14832, I14833)
--	I14840 = NAND(WX4881, WX4578)
--	I14841 = NAND(WX4881, I14840)
--	I14842 = NAND(WX4578, I14840)
--	I14839 = NAND(I14841, I14842)
--	I14847 = NAND(WX4642, I14839)
--	I14848 = NAND(WX4642, I14847)
--	I14849 = NAND(I14839, I14847)
--	I14838 = NAND(I14848, I14849)
--	I14855 = NAND(WX4706, WX4770)
--	I14856 = NAND(WX4706, I14855)
--	I14857 = NAND(WX4770, I14855)
--	I14854 = NAND(I14856, I14857)
--	I14862 = NAND(I14838, I14854)
--	I14863 = NAND(I14838, I14862)
--	I14864 = NAND(I14854, I14862)
--	WX4806 = NAND(I14863, I14864)
--	I14871 = NAND(WX4881, WX4580)
--	I14872 = NAND(WX4881, I14871)
--	I14873 = NAND(WX4580, I14871)
--	I14870 = NAND(I14872, I14873)
--	I14878 = NAND(WX4644, I14870)
--	I14879 = NAND(WX4644, I14878)
--	I14880 = NAND(I14870, I14878)
--	I14869 = NAND(I14879, I14880)
--	I14886 = NAND(WX4708, WX4772)
--	I14887 = NAND(WX4708, I14886)
--	I14888 = NAND(WX4772, I14886)
--	I14885 = NAND(I14887, I14888)
--	I14893 = NAND(I14869, I14885)
--	I14894 = NAND(I14869, I14893)
--	I14895 = NAND(I14885, I14893)
--	WX4807 = NAND(I14894, I14895)
--	I14902 = NAND(WX4881, WX4582)
--	I14903 = NAND(WX4881, I14902)
--	I14904 = NAND(WX4582, I14902)
--	I14901 = NAND(I14903, I14904)
--	I14909 = NAND(WX4646, I14901)
--	I14910 = NAND(WX4646, I14909)
--	I14911 = NAND(I14901, I14909)
--	I14900 = NAND(I14910, I14911)
--	I14917 = NAND(WX4710, WX4774)
--	I14918 = NAND(WX4710, I14917)
--	I14919 = NAND(WX4774, I14917)
--	I14916 = NAND(I14918, I14919)
--	I14924 = NAND(I14900, I14916)
--	I14925 = NAND(I14900, I14924)
--	I14926 = NAND(I14916, I14924)
--	WX4808 = NAND(I14925, I14926)
--	I14933 = NAND(WX4881, WX4584)
--	I14934 = NAND(WX4881, I14933)
--	I14935 = NAND(WX4584, I14933)
--	I14932 = NAND(I14934, I14935)
--	I14940 = NAND(WX4648, I14932)
--	I14941 = NAND(WX4648, I14940)
--	I14942 = NAND(I14932, I14940)
--	I14931 = NAND(I14941, I14942)
--	I14948 = NAND(WX4712, WX4776)
--	I14949 = NAND(WX4712, I14948)
--	I14950 = NAND(WX4776, I14948)
--	I14947 = NAND(I14949, I14950)
--	I14955 = NAND(I14931, I14947)
--	I14956 = NAND(I14931, I14955)
--	I14957 = NAND(I14947, I14955)
--	WX4809 = NAND(I14956, I14957)
--	I14964 = NAND(WX4881, WX4586)
--	I14965 = NAND(WX4881, I14964)
--	I14966 = NAND(WX4586, I14964)
--	I14963 = NAND(I14965, I14966)
--	I14971 = NAND(WX4650, I14963)
--	I14972 = NAND(WX4650, I14971)
--	I14973 = NAND(I14963, I14971)
--	I14962 = NAND(I14972, I14973)
--	I14979 = NAND(WX4714, WX4778)
--	I14980 = NAND(WX4714, I14979)
--	I14981 = NAND(WX4778, I14979)
--	I14978 = NAND(I14980, I14981)
--	I14986 = NAND(I14962, I14978)
--	I14987 = NAND(I14962, I14986)
--	I14988 = NAND(I14978, I14986)
--	WX4810 = NAND(I14987, I14988)
--	I15067 = NAND(WX4459, WX4364)
--	I15068 = NAND(WX4459, I15067)
--	I15069 = NAND(WX4364, I15067)
--	WX4885 = NAND(I15068, I15069)
--	I15080 = NAND(WX4460, WX4366)
--	I15081 = NAND(WX4460, I15080)
--	I15082 = NAND(WX4366, I15080)
--	WX4892 = NAND(I15081, I15082)
--	I15093 = NAND(WX4461, WX4368)
--	I15094 = NAND(WX4461, I15093)
--	I15095 = NAND(WX4368, I15093)
--	WX4899 = NAND(I15094, I15095)
--	I15106 = NAND(WX4462, WX4370)
--	I15107 = NAND(WX4462, I15106)
--	I15108 = NAND(WX4370, I15106)
--	WX4906 = NAND(I15107, I15108)
--	I15119 = NAND(WX4463, WX4372)
--	I15120 = NAND(WX4463, I15119)
--	I15121 = NAND(WX4372, I15119)
--	WX4913 = NAND(I15120, I15121)
--	I15132 = NAND(WX4464, WX4374)
--	I15133 = NAND(WX4464, I15132)
--	I15134 = NAND(WX4374, I15132)
--	WX4920 = NAND(I15133, I15134)
--	I15145 = NAND(WX4465, WX4376)
--	I15146 = NAND(WX4465, I15145)
--	I15147 = NAND(WX4376, I15145)
--	WX4927 = NAND(I15146, I15147)
--	I15158 = NAND(WX4466, WX4378)
--	I15159 = NAND(WX4466, I15158)
--	I15160 = NAND(WX4378, I15158)
--	WX4934 = NAND(I15159, I15160)
--	I15171 = NAND(WX4467, WX4380)
--	I15172 = NAND(WX4467, I15171)
--	I15173 = NAND(WX4380, I15171)
--	WX4941 = NAND(I15172, I15173)
--	I15184 = NAND(WX4468, WX4382)
--	I15185 = NAND(WX4468, I15184)
--	I15186 = NAND(WX4382, I15184)
--	WX4948 = NAND(I15185, I15186)
--	I15197 = NAND(WX4469, WX4384)
--	I15198 = NAND(WX4469, I15197)
--	I15199 = NAND(WX4384, I15197)
--	WX4955 = NAND(I15198, I15199)
--	I15210 = NAND(WX4470, WX4386)
--	I15211 = NAND(WX4470, I15210)
--	I15212 = NAND(WX4386, I15210)
--	WX4962 = NAND(I15211, I15212)
--	I15223 = NAND(WX4471, WX4388)
--	I15224 = NAND(WX4471, I15223)
--	I15225 = NAND(WX4388, I15223)
--	WX4969 = NAND(I15224, I15225)
--	I15236 = NAND(WX4472, WX4390)
--	I15237 = NAND(WX4472, I15236)
--	I15238 = NAND(WX4390, I15236)
--	WX4976 = NAND(I15237, I15238)
--	I15249 = NAND(WX4473, WX4392)
--	I15250 = NAND(WX4473, I15249)
--	I15251 = NAND(WX4392, I15249)
--	WX4983 = NAND(I15250, I15251)
--	I15262 = NAND(WX4474, WX4394)
--	I15263 = NAND(WX4474, I15262)
--	I15264 = NAND(WX4394, I15262)
--	WX4990 = NAND(I15263, I15264)
--	I15275 = NAND(WX4475, WX4396)
--	I15276 = NAND(WX4475, I15275)
--	I15277 = NAND(WX4396, I15275)
--	WX4997 = NAND(I15276, I15277)
--	I15288 = NAND(WX4476, WX4398)
--	I15289 = NAND(WX4476, I15288)
--	I15290 = NAND(WX4398, I15288)
--	WX5004 = NAND(I15289, I15290)
--	I15301 = NAND(WX4477, WX4400)
--	I15302 = NAND(WX4477, I15301)
--	I15303 = NAND(WX4400, I15301)
--	WX5011 = NAND(I15302, I15303)
--	I15314 = NAND(WX4478, WX4402)
--	I15315 = NAND(WX4478, I15314)
--	I15316 = NAND(WX4402, I15314)
--	WX5018 = NAND(I15315, I15316)
--	I15327 = NAND(WX4479, WX4404)
--	I15328 = NAND(WX4479, I15327)
--	I15329 = NAND(WX4404, I15327)
--	WX5025 = NAND(I15328, I15329)
--	I15340 = NAND(WX4480, WX4406)
--	I15341 = NAND(WX4480, I15340)
--	I15342 = NAND(WX4406, I15340)
--	WX5032 = NAND(I15341, I15342)
--	I15353 = NAND(WX4481, WX4408)
--	I15354 = NAND(WX4481, I15353)
--	I15355 = NAND(WX4408, I15353)
--	WX5039 = NAND(I15354, I15355)
--	I15366 = NAND(WX4482, WX4410)
--	I15367 = NAND(WX4482, I15366)
--	I15368 = NAND(WX4410, I15366)
--	WX5046 = NAND(I15367, I15368)
--	I15379 = NAND(WX4483, WX4412)
--	I15380 = NAND(WX4483, I15379)
--	I15381 = NAND(WX4412, I15379)
--	WX5053 = NAND(I15380, I15381)
--	I15392 = NAND(WX4484, WX4414)
--	I15393 = NAND(WX4484, I15392)
--	I15394 = NAND(WX4414, I15392)
--	WX5060 = NAND(I15393, I15394)
--	I15405 = NAND(WX4485, WX4416)
--	I15406 = NAND(WX4485, I15405)
--	I15407 = NAND(WX4416, I15405)
--	WX5067 = NAND(I15406, I15407)
--	I15418 = NAND(WX4486, WX4418)
--	I15419 = NAND(WX4486, I15418)
--	I15420 = NAND(WX4418, I15418)
--	WX5074 = NAND(I15419, I15420)
--	I15431 = NAND(WX4487, WX4420)
--	I15432 = NAND(WX4487, I15431)
--	I15433 = NAND(WX4420, I15431)
--	WX5081 = NAND(I15432, I15433)
--	I15444 = NAND(WX4488, WX4422)
--	I15445 = NAND(WX4488, I15444)
--	I15446 = NAND(WX4422, I15444)
--	WX5088 = NAND(I15445, I15446)
--	I15457 = NAND(WX4489, WX4424)
--	I15458 = NAND(WX4489, I15457)
--	I15459 = NAND(WX4424, I15457)
--	WX5095 = NAND(I15458, I15459)
--	I15470 = NAND(WX4490, WX4426)
--	I15471 = NAND(WX4490, I15470)
--	I15472 = NAND(WX4426, I15470)
--	WX5102 = NAND(I15471, I15472)
--	I15485 = NAND(WX4506, CRC_OUT_6_31)
--	I15486 = NAND(WX4506, I15485)
--	I15487 = NAND(CRC_OUT_6_31, I15485)
--	I15484 = NAND(I15486, I15487)
--	I15492 = NAND(CRC_OUT_6_15, I15484)
--	I15493 = NAND(CRC_OUT_6_15, I15492)
--	I15494 = NAND(I15484, I15492)
--	WX5110 = NAND(I15493, I15494)
--	I15500 = NAND(WX4511, CRC_OUT_6_31)
--	I15501 = NAND(WX4511, I15500)
--	I15502 = NAND(CRC_OUT_6_31, I15500)
--	I15499 = NAND(I15501, I15502)
--	I15507 = NAND(CRC_OUT_6_10, I15499)
--	I15508 = NAND(CRC_OUT_6_10, I15507)
--	I15509 = NAND(I15499, I15507)
--	WX5111 = NAND(I15508, I15509)
--	I15515 = NAND(WX4518, CRC_OUT_6_31)
--	I15516 = NAND(WX4518, I15515)
--	I15517 = NAND(CRC_OUT_6_31, I15515)
--	I15514 = NAND(I15516, I15517)
--	I15522 = NAND(CRC_OUT_6_3, I15514)
--	I15523 = NAND(CRC_OUT_6_3, I15522)
--	I15524 = NAND(I15514, I15522)
--	WX5112 = NAND(I15523, I15524)
--	I15529 = NAND(WX4522, CRC_OUT_6_31)
--	I15530 = NAND(WX4522, I15529)
--	I15531 = NAND(CRC_OUT_6_31, I15529)
--	WX5113 = NAND(I15530, I15531)
--	I15536 = NAND(WX4491, CRC_OUT_6_30)
--	I15537 = NAND(WX4491, I15536)
--	I15538 = NAND(CRC_OUT_6_30, I15536)
--	WX5114 = NAND(I15537, I15538)
--	I15543 = NAND(WX4492, CRC_OUT_6_29)
--	I15544 = NAND(WX4492, I15543)
--	I15545 = NAND(CRC_OUT_6_29, I15543)
--	WX5115 = NAND(I15544, I15545)
--	I15550 = NAND(WX4493, CRC_OUT_6_28)
--	I15551 = NAND(WX4493, I15550)
--	I15552 = NAND(CRC_OUT_6_28, I15550)
--	WX5116 = NAND(I15551, I15552)
--	I15557 = NAND(WX4494, CRC_OUT_6_27)
--	I15558 = NAND(WX4494, I15557)
--	I15559 = NAND(CRC_OUT_6_27, I15557)
--	WX5117 = NAND(I15558, I15559)
--	I15564 = NAND(WX4495, CRC_OUT_6_26)
--	I15565 = NAND(WX4495, I15564)
--	I15566 = NAND(CRC_OUT_6_26, I15564)
--	WX5118 = NAND(I15565, I15566)
--	I15571 = NAND(WX4496, CRC_OUT_6_25)
--	I15572 = NAND(WX4496, I15571)
--	I15573 = NAND(CRC_OUT_6_25, I15571)
--	WX5119 = NAND(I15572, I15573)
--	I15578 = NAND(WX4497, CRC_OUT_6_24)
--	I15579 = NAND(WX4497, I15578)
--	I15580 = NAND(CRC_OUT_6_24, I15578)
--	WX5120 = NAND(I15579, I15580)
--	I15585 = NAND(WX4498, CRC_OUT_6_23)
--	I15586 = NAND(WX4498, I15585)
--	I15587 = NAND(CRC_OUT_6_23, I15585)
--	WX5121 = NAND(I15586, I15587)
--	I15592 = NAND(WX4499, CRC_OUT_6_22)
--	I15593 = NAND(WX4499, I15592)
--	I15594 = NAND(CRC_OUT_6_22, I15592)
--	WX5122 = NAND(I15593, I15594)
--	I15599 = NAND(WX4500, CRC_OUT_6_21)
--	I15600 = NAND(WX4500, I15599)
--	I15601 = NAND(CRC_OUT_6_21, I15599)
--	WX5123 = NAND(I15600, I15601)
--	I15606 = NAND(WX4501, CRC_OUT_6_20)
--	I15607 = NAND(WX4501, I15606)
--	I15608 = NAND(CRC_OUT_6_20, I15606)
--	WX5124 = NAND(I15607, I15608)
--	I15613 = NAND(WX4502, CRC_OUT_6_19)
--	I15614 = NAND(WX4502, I15613)
--	I15615 = NAND(CRC_OUT_6_19, I15613)
--	WX5125 = NAND(I15614, I15615)
--	I15620 = NAND(WX4503, CRC_OUT_6_18)
--	I15621 = NAND(WX4503, I15620)
--	I15622 = NAND(CRC_OUT_6_18, I15620)
--	WX5126 = NAND(I15621, I15622)
--	I15627 = NAND(WX4504, CRC_OUT_6_17)
--	I15628 = NAND(WX4504, I15627)
--	I15629 = NAND(CRC_OUT_6_17, I15627)
--	WX5127 = NAND(I15628, I15629)
--	I15634 = NAND(WX4505, CRC_OUT_6_16)
--	I15635 = NAND(WX4505, I15634)
--	I15636 = NAND(CRC_OUT_6_16, I15634)
--	WX5128 = NAND(I15635, I15636)
--	I15641 = NAND(WX4507, CRC_OUT_6_14)
--	I15642 = NAND(WX4507, I15641)
--	I15643 = NAND(CRC_OUT_6_14, I15641)
--	WX5129 = NAND(I15642, I15643)
--	I15648 = NAND(WX4508, CRC_OUT_6_13)
--	I15649 = NAND(WX4508, I15648)
--	I15650 = NAND(CRC_OUT_6_13, I15648)
--	WX5130 = NAND(I15649, I15650)
--	I15655 = NAND(WX4509, CRC_OUT_6_12)
--	I15656 = NAND(WX4509, I15655)
--	I15657 = NAND(CRC_OUT_6_12, I15655)
--	WX5131 = NAND(I15656, I15657)
--	I15662 = NAND(WX4510, CRC_OUT_6_11)
--	I15663 = NAND(WX4510, I15662)
--	I15664 = NAND(CRC_OUT_6_11, I15662)
--	WX5132 = NAND(I15663, I15664)
--	I15669 = NAND(WX4512, CRC_OUT_6_9)
--	I15670 = NAND(WX4512, I15669)
--	I15671 = NAND(CRC_OUT_6_9, I15669)
--	WX5133 = NAND(I15670, I15671)
--	I15676 = NAND(WX4513, CRC_OUT_6_8)
--	I15677 = NAND(WX4513, I15676)
--	I15678 = NAND(CRC_OUT_6_8, I15676)
--	WX5134 = NAND(I15677, I15678)
--	I15683 = NAND(WX4514, CRC_OUT_6_7)
--	I15684 = NAND(WX4514, I15683)
--	I15685 = NAND(CRC_OUT_6_7, I15683)
--	WX5135 = NAND(I15684, I15685)
--	I15690 = NAND(WX4515, CRC_OUT_6_6)
--	I15691 = NAND(WX4515, I15690)
--	I15692 = NAND(CRC_OUT_6_6, I15690)
--	WX5136 = NAND(I15691, I15692)
--	I15697 = NAND(WX4516, CRC_OUT_6_5)
--	I15698 = NAND(WX4516, I15697)
--	I15699 = NAND(CRC_OUT_6_5, I15697)
--	WX5137 = NAND(I15698, I15699)
--	I15704 = NAND(WX4517, CRC_OUT_6_4)
--	I15705 = NAND(WX4517, I15704)
--	I15706 = NAND(CRC_OUT_6_4, I15704)
--	WX5138 = NAND(I15705, I15706)
--	I15711 = NAND(WX4519, CRC_OUT_6_2)
--	I15712 = NAND(WX4519, I15711)
--	I15713 = NAND(CRC_OUT_6_2, I15711)
--	WX5139 = NAND(I15712, I15713)
--	I15718 = NAND(WX4520, CRC_OUT_6_1)
--	I15719 = NAND(WX4520, I15718)
--	I15720 = NAND(CRC_OUT_6_1, I15718)
--	WX5140 = NAND(I15719, I15720)
--	I15725 = NAND(WX4521, CRC_OUT_6_0)
--	I15726 = NAND(WX4521, I15725)
--	I15727 = NAND(CRC_OUT_6_0, I15725)
--	WX5141 = NAND(I15726, I15727)
--	I18008 = NAND(WX6173, WX5817)
--	I18009 = NAND(WX6173, I18008)
--	I18010 = NAND(WX5817, I18008)
--	I18007 = NAND(I18009, I18010)
--	I18015 = NAND(WX5881, I18007)
--	I18016 = NAND(WX5881, I18015)
--	I18017 = NAND(I18007, I18015)
--	I18006 = NAND(I18016, I18017)
--	I18023 = NAND(WX5945, WX6009)
--	I18024 = NAND(WX5945, I18023)
--	I18025 = NAND(WX6009, I18023)
--	I18022 = NAND(I18024, I18025)
--	I18030 = NAND(I18006, I18022)
--	I18031 = NAND(I18006, I18030)
--	I18032 = NAND(I18022, I18030)
--	WX6072 = NAND(I18031, I18032)
--	I18039 = NAND(WX6173, WX5819)
--	I18040 = NAND(WX6173, I18039)
--	I18041 = NAND(WX5819, I18039)
--	I18038 = NAND(I18040, I18041)
--	I18046 = NAND(WX5883, I18038)
--	I18047 = NAND(WX5883, I18046)
--	I18048 = NAND(I18038, I18046)
--	I18037 = NAND(I18047, I18048)
--	I18054 = NAND(WX5947, WX6011)
--	I18055 = NAND(WX5947, I18054)
--	I18056 = NAND(WX6011, I18054)
--	I18053 = NAND(I18055, I18056)
--	I18061 = NAND(I18037, I18053)
--	I18062 = NAND(I18037, I18061)
--	I18063 = NAND(I18053, I18061)
--	WX6073 = NAND(I18062, I18063)
--	I18070 = NAND(WX6173, WX5821)
--	I18071 = NAND(WX6173, I18070)
--	I18072 = NAND(WX5821, I18070)
--	I18069 = NAND(I18071, I18072)
--	I18077 = NAND(WX5885, I18069)
--	I18078 = NAND(WX5885, I18077)
--	I18079 = NAND(I18069, I18077)
--	I18068 = NAND(I18078, I18079)
--	I18085 = NAND(WX5949, WX6013)
--	I18086 = NAND(WX5949, I18085)
--	I18087 = NAND(WX6013, I18085)
--	I18084 = NAND(I18086, I18087)
--	I18092 = NAND(I18068, I18084)
--	I18093 = NAND(I18068, I18092)
--	I18094 = NAND(I18084, I18092)
--	WX6074 = NAND(I18093, I18094)
--	I18101 = NAND(WX6173, WX5823)
--	I18102 = NAND(WX6173, I18101)
--	I18103 = NAND(WX5823, I18101)
--	I18100 = NAND(I18102, I18103)
--	I18108 = NAND(WX5887, I18100)
--	I18109 = NAND(WX5887, I18108)
--	I18110 = NAND(I18100, I18108)
--	I18099 = NAND(I18109, I18110)
--	I18116 = NAND(WX5951, WX6015)
--	I18117 = NAND(WX5951, I18116)
--	I18118 = NAND(WX6015, I18116)
--	I18115 = NAND(I18117, I18118)
--	I18123 = NAND(I18099, I18115)
--	I18124 = NAND(I18099, I18123)
--	I18125 = NAND(I18115, I18123)
--	WX6075 = NAND(I18124, I18125)
--	I18132 = NAND(WX6173, WX5825)
--	I18133 = NAND(WX6173, I18132)
--	I18134 = NAND(WX5825, I18132)
--	I18131 = NAND(I18133, I18134)
--	I18139 = NAND(WX5889, I18131)
--	I18140 = NAND(WX5889, I18139)
--	I18141 = NAND(I18131, I18139)
--	I18130 = NAND(I18140, I18141)
--	I18147 = NAND(WX5953, WX6017)
--	I18148 = NAND(WX5953, I18147)
--	I18149 = NAND(WX6017, I18147)
--	I18146 = NAND(I18148, I18149)
--	I18154 = NAND(I18130, I18146)
--	I18155 = NAND(I18130, I18154)
--	I18156 = NAND(I18146, I18154)
--	WX6076 = NAND(I18155, I18156)
--	I18163 = NAND(WX6173, WX5827)
--	I18164 = NAND(WX6173, I18163)
--	I18165 = NAND(WX5827, I18163)
--	I18162 = NAND(I18164, I18165)
--	I18170 = NAND(WX5891, I18162)
--	I18171 = NAND(WX5891, I18170)
--	I18172 = NAND(I18162, I18170)
--	I18161 = NAND(I18171, I18172)
--	I18178 = NAND(WX5955, WX6019)
--	I18179 = NAND(WX5955, I18178)
--	I18180 = NAND(WX6019, I18178)
--	I18177 = NAND(I18179, I18180)
--	I18185 = NAND(I18161, I18177)
--	I18186 = NAND(I18161, I18185)
--	I18187 = NAND(I18177, I18185)
--	WX6077 = NAND(I18186, I18187)
--	I18194 = NAND(WX6173, WX5829)
--	I18195 = NAND(WX6173, I18194)
--	I18196 = NAND(WX5829, I18194)
--	I18193 = NAND(I18195, I18196)
--	I18201 = NAND(WX5893, I18193)
--	I18202 = NAND(WX5893, I18201)
--	I18203 = NAND(I18193, I18201)
--	I18192 = NAND(I18202, I18203)
--	I18209 = NAND(WX5957, WX6021)
--	I18210 = NAND(WX5957, I18209)
--	I18211 = NAND(WX6021, I18209)
--	I18208 = NAND(I18210, I18211)
--	I18216 = NAND(I18192, I18208)
--	I18217 = NAND(I18192, I18216)
--	I18218 = NAND(I18208, I18216)
--	WX6078 = NAND(I18217, I18218)
--	I18225 = NAND(WX6173, WX5831)
--	I18226 = NAND(WX6173, I18225)
--	I18227 = NAND(WX5831, I18225)
--	I18224 = NAND(I18226, I18227)
--	I18232 = NAND(WX5895, I18224)
--	I18233 = NAND(WX5895, I18232)
--	I18234 = NAND(I18224, I18232)
--	I18223 = NAND(I18233, I18234)
--	I18240 = NAND(WX5959, WX6023)
--	I18241 = NAND(WX5959, I18240)
--	I18242 = NAND(WX6023, I18240)
--	I18239 = NAND(I18241, I18242)
--	I18247 = NAND(I18223, I18239)
--	I18248 = NAND(I18223, I18247)
--	I18249 = NAND(I18239, I18247)
--	WX6079 = NAND(I18248, I18249)
--	I18256 = NAND(WX6173, WX5833)
--	I18257 = NAND(WX6173, I18256)
--	I18258 = NAND(WX5833, I18256)
--	I18255 = NAND(I18257, I18258)
--	I18263 = NAND(WX5897, I18255)
--	I18264 = NAND(WX5897, I18263)
--	I18265 = NAND(I18255, I18263)
--	I18254 = NAND(I18264, I18265)
--	I18271 = NAND(WX5961, WX6025)
--	I18272 = NAND(WX5961, I18271)
--	I18273 = NAND(WX6025, I18271)
--	I18270 = NAND(I18272, I18273)
--	I18278 = NAND(I18254, I18270)
--	I18279 = NAND(I18254, I18278)
--	I18280 = NAND(I18270, I18278)
--	WX6080 = NAND(I18279, I18280)
--	I18287 = NAND(WX6173, WX5835)
--	I18288 = NAND(WX6173, I18287)
--	I18289 = NAND(WX5835, I18287)
--	I18286 = NAND(I18288, I18289)
--	I18294 = NAND(WX5899, I18286)
--	I18295 = NAND(WX5899, I18294)
--	I18296 = NAND(I18286, I18294)
--	I18285 = NAND(I18295, I18296)
--	I18302 = NAND(WX5963, WX6027)
--	I18303 = NAND(WX5963, I18302)
--	I18304 = NAND(WX6027, I18302)
--	I18301 = NAND(I18303, I18304)
--	I18309 = NAND(I18285, I18301)
--	I18310 = NAND(I18285, I18309)
--	I18311 = NAND(I18301, I18309)
--	WX6081 = NAND(I18310, I18311)
--	I18318 = NAND(WX6173, WX5837)
--	I18319 = NAND(WX6173, I18318)
--	I18320 = NAND(WX5837, I18318)
--	I18317 = NAND(I18319, I18320)
--	I18325 = NAND(WX5901, I18317)
--	I18326 = NAND(WX5901, I18325)
--	I18327 = NAND(I18317, I18325)
--	I18316 = NAND(I18326, I18327)
--	I18333 = NAND(WX5965, WX6029)
--	I18334 = NAND(WX5965, I18333)
--	I18335 = NAND(WX6029, I18333)
--	I18332 = NAND(I18334, I18335)
--	I18340 = NAND(I18316, I18332)
--	I18341 = NAND(I18316, I18340)
--	I18342 = NAND(I18332, I18340)
--	WX6082 = NAND(I18341, I18342)
--	I18349 = NAND(WX6173, WX5839)
--	I18350 = NAND(WX6173, I18349)
--	I18351 = NAND(WX5839, I18349)
--	I18348 = NAND(I18350, I18351)
--	I18356 = NAND(WX5903, I18348)
--	I18357 = NAND(WX5903, I18356)
--	I18358 = NAND(I18348, I18356)
--	I18347 = NAND(I18357, I18358)
--	I18364 = NAND(WX5967, WX6031)
--	I18365 = NAND(WX5967, I18364)
--	I18366 = NAND(WX6031, I18364)
--	I18363 = NAND(I18365, I18366)
--	I18371 = NAND(I18347, I18363)
--	I18372 = NAND(I18347, I18371)
--	I18373 = NAND(I18363, I18371)
--	WX6083 = NAND(I18372, I18373)
--	I18380 = NAND(WX6173, WX5841)
--	I18381 = NAND(WX6173, I18380)
--	I18382 = NAND(WX5841, I18380)
--	I18379 = NAND(I18381, I18382)
--	I18387 = NAND(WX5905, I18379)
--	I18388 = NAND(WX5905, I18387)
--	I18389 = NAND(I18379, I18387)
--	I18378 = NAND(I18388, I18389)
--	I18395 = NAND(WX5969, WX6033)
--	I18396 = NAND(WX5969, I18395)
--	I18397 = NAND(WX6033, I18395)
--	I18394 = NAND(I18396, I18397)
--	I18402 = NAND(I18378, I18394)
--	I18403 = NAND(I18378, I18402)
--	I18404 = NAND(I18394, I18402)
--	WX6084 = NAND(I18403, I18404)
--	I18411 = NAND(WX6173, WX5843)
--	I18412 = NAND(WX6173, I18411)
--	I18413 = NAND(WX5843, I18411)
--	I18410 = NAND(I18412, I18413)
--	I18418 = NAND(WX5907, I18410)
--	I18419 = NAND(WX5907, I18418)
--	I18420 = NAND(I18410, I18418)
--	I18409 = NAND(I18419, I18420)
--	I18426 = NAND(WX5971, WX6035)
--	I18427 = NAND(WX5971, I18426)
--	I18428 = NAND(WX6035, I18426)
--	I18425 = NAND(I18427, I18428)
--	I18433 = NAND(I18409, I18425)
--	I18434 = NAND(I18409, I18433)
--	I18435 = NAND(I18425, I18433)
--	WX6085 = NAND(I18434, I18435)
--	I18442 = NAND(WX6173, WX5845)
--	I18443 = NAND(WX6173, I18442)
--	I18444 = NAND(WX5845, I18442)
--	I18441 = NAND(I18443, I18444)
--	I18449 = NAND(WX5909, I18441)
--	I18450 = NAND(WX5909, I18449)
--	I18451 = NAND(I18441, I18449)
--	I18440 = NAND(I18450, I18451)
--	I18457 = NAND(WX5973, WX6037)
--	I18458 = NAND(WX5973, I18457)
--	I18459 = NAND(WX6037, I18457)
--	I18456 = NAND(I18458, I18459)
--	I18464 = NAND(I18440, I18456)
--	I18465 = NAND(I18440, I18464)
--	I18466 = NAND(I18456, I18464)
--	WX6086 = NAND(I18465, I18466)
--	I18473 = NAND(WX6173, WX5847)
--	I18474 = NAND(WX6173, I18473)
--	I18475 = NAND(WX5847, I18473)
--	I18472 = NAND(I18474, I18475)
--	I18480 = NAND(WX5911, I18472)
--	I18481 = NAND(WX5911, I18480)
--	I18482 = NAND(I18472, I18480)
--	I18471 = NAND(I18481, I18482)
--	I18488 = NAND(WX5975, WX6039)
--	I18489 = NAND(WX5975, I18488)
--	I18490 = NAND(WX6039, I18488)
--	I18487 = NAND(I18489, I18490)
--	I18495 = NAND(I18471, I18487)
--	I18496 = NAND(I18471, I18495)
--	I18497 = NAND(I18487, I18495)
--	WX6087 = NAND(I18496, I18497)
--	I18504 = NAND(WX6174, WX5849)
--	I18505 = NAND(WX6174, I18504)
--	I18506 = NAND(WX5849, I18504)
--	I18503 = NAND(I18505, I18506)
--	I18511 = NAND(WX5913, I18503)
--	I18512 = NAND(WX5913, I18511)
--	I18513 = NAND(I18503, I18511)
--	I18502 = NAND(I18512, I18513)
--	I18519 = NAND(WX5977, WX6041)
--	I18520 = NAND(WX5977, I18519)
--	I18521 = NAND(WX6041, I18519)
--	I18518 = NAND(I18520, I18521)
--	I18526 = NAND(I18502, I18518)
--	I18527 = NAND(I18502, I18526)
--	I18528 = NAND(I18518, I18526)
--	WX6088 = NAND(I18527, I18528)
--	I18535 = NAND(WX6174, WX5851)
--	I18536 = NAND(WX6174, I18535)
--	I18537 = NAND(WX5851, I18535)
--	I18534 = NAND(I18536, I18537)
--	I18542 = NAND(WX5915, I18534)
--	I18543 = NAND(WX5915, I18542)
--	I18544 = NAND(I18534, I18542)
--	I18533 = NAND(I18543, I18544)
--	I18550 = NAND(WX5979, WX6043)
--	I18551 = NAND(WX5979, I18550)
--	I18552 = NAND(WX6043, I18550)
--	I18549 = NAND(I18551, I18552)
--	I18557 = NAND(I18533, I18549)
--	I18558 = NAND(I18533, I18557)
--	I18559 = NAND(I18549, I18557)
--	WX6089 = NAND(I18558, I18559)
--	I18566 = NAND(WX6174, WX5853)
--	I18567 = NAND(WX6174, I18566)
--	I18568 = NAND(WX5853, I18566)
--	I18565 = NAND(I18567, I18568)
--	I18573 = NAND(WX5917, I18565)
--	I18574 = NAND(WX5917, I18573)
--	I18575 = NAND(I18565, I18573)
--	I18564 = NAND(I18574, I18575)
--	I18581 = NAND(WX5981, WX6045)
--	I18582 = NAND(WX5981, I18581)
--	I18583 = NAND(WX6045, I18581)
--	I18580 = NAND(I18582, I18583)
--	I18588 = NAND(I18564, I18580)
--	I18589 = NAND(I18564, I18588)
--	I18590 = NAND(I18580, I18588)
--	WX6090 = NAND(I18589, I18590)
--	I18597 = NAND(WX6174, WX5855)
--	I18598 = NAND(WX6174, I18597)
--	I18599 = NAND(WX5855, I18597)
--	I18596 = NAND(I18598, I18599)
--	I18604 = NAND(WX5919, I18596)
--	I18605 = NAND(WX5919, I18604)
--	I18606 = NAND(I18596, I18604)
--	I18595 = NAND(I18605, I18606)
--	I18612 = NAND(WX5983, WX6047)
--	I18613 = NAND(WX5983, I18612)
--	I18614 = NAND(WX6047, I18612)
--	I18611 = NAND(I18613, I18614)
--	I18619 = NAND(I18595, I18611)
--	I18620 = NAND(I18595, I18619)
--	I18621 = NAND(I18611, I18619)
--	WX6091 = NAND(I18620, I18621)
--	I18628 = NAND(WX6174, WX5857)
--	I18629 = NAND(WX6174, I18628)
--	I18630 = NAND(WX5857, I18628)
--	I18627 = NAND(I18629, I18630)
--	I18635 = NAND(WX5921, I18627)
--	I18636 = NAND(WX5921, I18635)
--	I18637 = NAND(I18627, I18635)
--	I18626 = NAND(I18636, I18637)
--	I18643 = NAND(WX5985, WX6049)
--	I18644 = NAND(WX5985, I18643)
--	I18645 = NAND(WX6049, I18643)
--	I18642 = NAND(I18644, I18645)
--	I18650 = NAND(I18626, I18642)
--	I18651 = NAND(I18626, I18650)
--	I18652 = NAND(I18642, I18650)
--	WX6092 = NAND(I18651, I18652)
--	I18659 = NAND(WX6174, WX5859)
--	I18660 = NAND(WX6174, I18659)
--	I18661 = NAND(WX5859, I18659)
--	I18658 = NAND(I18660, I18661)
--	I18666 = NAND(WX5923, I18658)
--	I18667 = NAND(WX5923, I18666)
--	I18668 = NAND(I18658, I18666)
--	I18657 = NAND(I18667, I18668)
--	I18674 = NAND(WX5987, WX6051)
--	I18675 = NAND(WX5987, I18674)
--	I18676 = NAND(WX6051, I18674)
--	I18673 = NAND(I18675, I18676)
--	I18681 = NAND(I18657, I18673)
--	I18682 = NAND(I18657, I18681)
--	I18683 = NAND(I18673, I18681)
--	WX6093 = NAND(I18682, I18683)
--	I18690 = NAND(WX6174, WX5861)
--	I18691 = NAND(WX6174, I18690)
--	I18692 = NAND(WX5861, I18690)
--	I18689 = NAND(I18691, I18692)
--	I18697 = NAND(WX5925, I18689)
--	I18698 = NAND(WX5925, I18697)
--	I18699 = NAND(I18689, I18697)
--	I18688 = NAND(I18698, I18699)
--	I18705 = NAND(WX5989, WX6053)
--	I18706 = NAND(WX5989, I18705)
--	I18707 = NAND(WX6053, I18705)
--	I18704 = NAND(I18706, I18707)
--	I18712 = NAND(I18688, I18704)
--	I18713 = NAND(I18688, I18712)
--	I18714 = NAND(I18704, I18712)
--	WX6094 = NAND(I18713, I18714)
--	I18721 = NAND(WX6174, WX5863)
--	I18722 = NAND(WX6174, I18721)
--	I18723 = NAND(WX5863, I18721)
--	I18720 = NAND(I18722, I18723)
--	I18728 = NAND(WX5927, I18720)
--	I18729 = NAND(WX5927, I18728)
--	I18730 = NAND(I18720, I18728)
--	I18719 = NAND(I18729, I18730)
--	I18736 = NAND(WX5991, WX6055)
--	I18737 = NAND(WX5991, I18736)
--	I18738 = NAND(WX6055, I18736)
--	I18735 = NAND(I18737, I18738)
--	I18743 = NAND(I18719, I18735)
--	I18744 = NAND(I18719, I18743)
--	I18745 = NAND(I18735, I18743)
--	WX6095 = NAND(I18744, I18745)
--	I18752 = NAND(WX6174, WX5865)
--	I18753 = NAND(WX6174, I18752)
--	I18754 = NAND(WX5865, I18752)
--	I18751 = NAND(I18753, I18754)
--	I18759 = NAND(WX5929, I18751)
--	I18760 = NAND(WX5929, I18759)
--	I18761 = NAND(I18751, I18759)
--	I18750 = NAND(I18760, I18761)
--	I18767 = NAND(WX5993, WX6057)
--	I18768 = NAND(WX5993, I18767)
--	I18769 = NAND(WX6057, I18767)
--	I18766 = NAND(I18768, I18769)
--	I18774 = NAND(I18750, I18766)
--	I18775 = NAND(I18750, I18774)
--	I18776 = NAND(I18766, I18774)
--	WX6096 = NAND(I18775, I18776)
--	I18783 = NAND(WX6174, WX5867)
--	I18784 = NAND(WX6174, I18783)
--	I18785 = NAND(WX5867, I18783)
--	I18782 = NAND(I18784, I18785)
--	I18790 = NAND(WX5931, I18782)
--	I18791 = NAND(WX5931, I18790)
--	I18792 = NAND(I18782, I18790)
--	I18781 = NAND(I18791, I18792)
--	I18798 = NAND(WX5995, WX6059)
--	I18799 = NAND(WX5995, I18798)
--	I18800 = NAND(WX6059, I18798)
--	I18797 = NAND(I18799, I18800)
--	I18805 = NAND(I18781, I18797)
--	I18806 = NAND(I18781, I18805)
--	I18807 = NAND(I18797, I18805)
--	WX6097 = NAND(I18806, I18807)
--	I18814 = NAND(WX6174, WX5869)
--	I18815 = NAND(WX6174, I18814)
--	I18816 = NAND(WX5869, I18814)
--	I18813 = NAND(I18815, I18816)
--	I18821 = NAND(WX5933, I18813)
--	I18822 = NAND(WX5933, I18821)
--	I18823 = NAND(I18813, I18821)
--	I18812 = NAND(I18822, I18823)
--	I18829 = NAND(WX5997, WX6061)
--	I18830 = NAND(WX5997, I18829)
--	I18831 = NAND(WX6061, I18829)
--	I18828 = NAND(I18830, I18831)
--	I18836 = NAND(I18812, I18828)
--	I18837 = NAND(I18812, I18836)
--	I18838 = NAND(I18828, I18836)
--	WX6098 = NAND(I18837, I18838)
--	I18845 = NAND(WX6174, WX5871)
--	I18846 = NAND(WX6174, I18845)
--	I18847 = NAND(WX5871, I18845)
--	I18844 = NAND(I18846, I18847)
--	I18852 = NAND(WX5935, I18844)
--	I18853 = NAND(WX5935, I18852)
--	I18854 = NAND(I18844, I18852)
--	I18843 = NAND(I18853, I18854)
--	I18860 = NAND(WX5999, WX6063)
--	I18861 = NAND(WX5999, I18860)
--	I18862 = NAND(WX6063, I18860)
--	I18859 = NAND(I18861, I18862)
--	I18867 = NAND(I18843, I18859)
--	I18868 = NAND(I18843, I18867)
--	I18869 = NAND(I18859, I18867)
--	WX6099 = NAND(I18868, I18869)
--	I18876 = NAND(WX6174, WX5873)
--	I18877 = NAND(WX6174, I18876)
--	I18878 = NAND(WX5873, I18876)
--	I18875 = NAND(I18877, I18878)
--	I18883 = NAND(WX5937, I18875)
--	I18884 = NAND(WX5937, I18883)
--	I18885 = NAND(I18875, I18883)
--	I18874 = NAND(I18884, I18885)
--	I18891 = NAND(WX6001, WX6065)
--	I18892 = NAND(WX6001, I18891)
--	I18893 = NAND(WX6065, I18891)
--	I18890 = NAND(I18892, I18893)
--	I18898 = NAND(I18874, I18890)
--	I18899 = NAND(I18874, I18898)
--	I18900 = NAND(I18890, I18898)
--	WX6100 = NAND(I18899, I18900)
--	I18907 = NAND(WX6174, WX5875)
--	I18908 = NAND(WX6174, I18907)
--	I18909 = NAND(WX5875, I18907)
--	I18906 = NAND(I18908, I18909)
--	I18914 = NAND(WX5939, I18906)
--	I18915 = NAND(WX5939, I18914)
--	I18916 = NAND(I18906, I18914)
--	I18905 = NAND(I18915, I18916)
--	I18922 = NAND(WX6003, WX6067)
--	I18923 = NAND(WX6003, I18922)
--	I18924 = NAND(WX6067, I18922)
--	I18921 = NAND(I18923, I18924)
--	I18929 = NAND(I18905, I18921)
--	I18930 = NAND(I18905, I18929)
--	I18931 = NAND(I18921, I18929)
--	WX6101 = NAND(I18930, I18931)
--	I18938 = NAND(WX6174, WX5877)
--	I18939 = NAND(WX6174, I18938)
--	I18940 = NAND(WX5877, I18938)
--	I18937 = NAND(I18939, I18940)
--	I18945 = NAND(WX5941, I18937)
--	I18946 = NAND(WX5941, I18945)
--	I18947 = NAND(I18937, I18945)
--	I18936 = NAND(I18946, I18947)
--	I18953 = NAND(WX6005, WX6069)
--	I18954 = NAND(WX6005, I18953)
--	I18955 = NAND(WX6069, I18953)
--	I18952 = NAND(I18954, I18955)
--	I18960 = NAND(I18936, I18952)
--	I18961 = NAND(I18936, I18960)
--	I18962 = NAND(I18952, I18960)
--	WX6102 = NAND(I18961, I18962)
--	I18969 = NAND(WX6174, WX5879)
--	I18970 = NAND(WX6174, I18969)
--	I18971 = NAND(WX5879, I18969)
--	I18968 = NAND(I18970, I18971)
--	I18976 = NAND(WX5943, I18968)
--	I18977 = NAND(WX5943, I18976)
--	I18978 = NAND(I18968, I18976)
--	I18967 = NAND(I18977, I18978)
--	I18984 = NAND(WX6007, WX6071)
--	I18985 = NAND(WX6007, I18984)
--	I18986 = NAND(WX6071, I18984)
--	I18983 = NAND(I18985, I18986)
--	I18991 = NAND(I18967, I18983)
--	I18992 = NAND(I18967, I18991)
--	I18993 = NAND(I18983, I18991)
--	WX6103 = NAND(I18992, I18993)
--	I19072 = NAND(WX5752, WX5657)
--	I19073 = NAND(WX5752, I19072)
--	I19074 = NAND(WX5657, I19072)
--	WX6178 = NAND(I19073, I19074)
--	I19085 = NAND(WX5753, WX5659)
--	I19086 = NAND(WX5753, I19085)
--	I19087 = NAND(WX5659, I19085)
--	WX6185 = NAND(I19086, I19087)
--	I19098 = NAND(WX5754, WX5661)
--	I19099 = NAND(WX5754, I19098)
--	I19100 = NAND(WX5661, I19098)
--	WX6192 = NAND(I19099, I19100)
--	I19111 = NAND(WX5755, WX5663)
--	I19112 = NAND(WX5755, I19111)
--	I19113 = NAND(WX5663, I19111)
--	WX6199 = NAND(I19112, I19113)
--	I19124 = NAND(WX5756, WX5665)
--	I19125 = NAND(WX5756, I19124)
--	I19126 = NAND(WX5665, I19124)
--	WX6206 = NAND(I19125, I19126)
--	I19137 = NAND(WX5757, WX5667)
--	I19138 = NAND(WX5757, I19137)
--	I19139 = NAND(WX5667, I19137)
--	WX6213 = NAND(I19138, I19139)
--	I19150 = NAND(WX5758, WX5669)
--	I19151 = NAND(WX5758, I19150)
--	I19152 = NAND(WX5669, I19150)
--	WX6220 = NAND(I19151, I19152)
--	I19163 = NAND(WX5759, WX5671)
--	I19164 = NAND(WX5759, I19163)
--	I19165 = NAND(WX5671, I19163)
--	WX6227 = NAND(I19164, I19165)
--	I19176 = NAND(WX5760, WX5673)
--	I19177 = NAND(WX5760, I19176)
--	I19178 = NAND(WX5673, I19176)
--	WX6234 = NAND(I19177, I19178)
--	I19189 = NAND(WX5761, WX5675)
--	I19190 = NAND(WX5761, I19189)
--	I19191 = NAND(WX5675, I19189)
--	WX6241 = NAND(I19190, I19191)
--	I19202 = NAND(WX5762, WX5677)
--	I19203 = NAND(WX5762, I19202)
--	I19204 = NAND(WX5677, I19202)
--	WX6248 = NAND(I19203, I19204)
--	I19215 = NAND(WX5763, WX5679)
--	I19216 = NAND(WX5763, I19215)
--	I19217 = NAND(WX5679, I19215)
--	WX6255 = NAND(I19216, I19217)
--	I19228 = NAND(WX5764, WX5681)
--	I19229 = NAND(WX5764, I19228)
--	I19230 = NAND(WX5681, I19228)
--	WX6262 = NAND(I19229, I19230)
--	I19241 = NAND(WX5765, WX5683)
--	I19242 = NAND(WX5765, I19241)
--	I19243 = NAND(WX5683, I19241)
--	WX6269 = NAND(I19242, I19243)
--	I19254 = NAND(WX5766, WX5685)
--	I19255 = NAND(WX5766, I19254)
--	I19256 = NAND(WX5685, I19254)
--	WX6276 = NAND(I19255, I19256)
--	I19267 = NAND(WX5767, WX5687)
--	I19268 = NAND(WX5767, I19267)
--	I19269 = NAND(WX5687, I19267)
--	WX6283 = NAND(I19268, I19269)
--	I19280 = NAND(WX5768, WX5689)
--	I19281 = NAND(WX5768, I19280)
--	I19282 = NAND(WX5689, I19280)
--	WX6290 = NAND(I19281, I19282)
--	I19293 = NAND(WX5769, WX5691)
--	I19294 = NAND(WX5769, I19293)
--	I19295 = NAND(WX5691, I19293)
--	WX6297 = NAND(I19294, I19295)
--	I19306 = NAND(WX5770, WX5693)
--	I19307 = NAND(WX5770, I19306)
--	I19308 = NAND(WX5693, I19306)
--	WX6304 = NAND(I19307, I19308)
--	I19319 = NAND(WX5771, WX5695)
--	I19320 = NAND(WX5771, I19319)
--	I19321 = NAND(WX5695, I19319)
--	WX6311 = NAND(I19320, I19321)
--	I19332 = NAND(WX5772, WX5697)
--	I19333 = NAND(WX5772, I19332)
--	I19334 = NAND(WX5697, I19332)
--	WX6318 = NAND(I19333, I19334)
--	I19345 = NAND(WX5773, WX5699)
--	I19346 = NAND(WX5773, I19345)
--	I19347 = NAND(WX5699, I19345)
--	WX6325 = NAND(I19346, I19347)
--	I19358 = NAND(WX5774, WX5701)
--	I19359 = NAND(WX5774, I19358)
--	I19360 = NAND(WX5701, I19358)
--	WX6332 = NAND(I19359, I19360)
--	I19371 = NAND(WX5775, WX5703)
--	I19372 = NAND(WX5775, I19371)
--	I19373 = NAND(WX5703, I19371)
--	WX6339 = NAND(I19372, I19373)
--	I19384 = NAND(WX5776, WX5705)
--	I19385 = NAND(WX5776, I19384)
--	I19386 = NAND(WX5705, I19384)
--	WX6346 = NAND(I19385, I19386)
--	I19397 = NAND(WX5777, WX5707)
--	I19398 = NAND(WX5777, I19397)
--	I19399 = NAND(WX5707, I19397)
--	WX6353 = NAND(I19398, I19399)
--	I19410 = NAND(WX5778, WX5709)
--	I19411 = NAND(WX5778, I19410)
--	I19412 = NAND(WX5709, I19410)
--	WX6360 = NAND(I19411, I19412)
--	I19423 = NAND(WX5779, WX5711)
--	I19424 = NAND(WX5779, I19423)
--	I19425 = NAND(WX5711, I19423)
--	WX6367 = NAND(I19424, I19425)
--	I19436 = NAND(WX5780, WX5713)
--	I19437 = NAND(WX5780, I19436)
--	I19438 = NAND(WX5713, I19436)
--	WX6374 = NAND(I19437, I19438)
--	I19449 = NAND(WX5781, WX5715)
--	I19450 = NAND(WX5781, I19449)
--	I19451 = NAND(WX5715, I19449)
--	WX6381 = NAND(I19450, I19451)
--	I19462 = NAND(WX5782, WX5717)
--	I19463 = NAND(WX5782, I19462)
--	I19464 = NAND(WX5717, I19462)
--	WX6388 = NAND(I19463, I19464)
--	I19475 = NAND(WX5783, WX5719)
--	I19476 = NAND(WX5783, I19475)
--	I19477 = NAND(WX5719, I19475)
--	WX6395 = NAND(I19476, I19477)
--	I19490 = NAND(WX5799, CRC_OUT_5_31)
--	I19491 = NAND(WX5799, I19490)
--	I19492 = NAND(CRC_OUT_5_31, I19490)
--	I19489 = NAND(I19491, I19492)
--	I19497 = NAND(CRC_OUT_5_15, I19489)
--	I19498 = NAND(CRC_OUT_5_15, I19497)
--	I19499 = NAND(I19489, I19497)
--	WX6403 = NAND(I19498, I19499)
--	I19505 = NAND(WX5804, CRC_OUT_5_31)
--	I19506 = NAND(WX5804, I19505)
--	I19507 = NAND(CRC_OUT_5_31, I19505)
--	I19504 = NAND(I19506, I19507)
--	I19512 = NAND(CRC_OUT_5_10, I19504)
--	I19513 = NAND(CRC_OUT_5_10, I19512)
--	I19514 = NAND(I19504, I19512)
--	WX6404 = NAND(I19513, I19514)
--	I19520 = NAND(WX5811, CRC_OUT_5_31)
--	I19521 = NAND(WX5811, I19520)
--	I19522 = NAND(CRC_OUT_5_31, I19520)
--	I19519 = NAND(I19521, I19522)
--	I19527 = NAND(CRC_OUT_5_3, I19519)
--	I19528 = NAND(CRC_OUT_5_3, I19527)
--	I19529 = NAND(I19519, I19527)
--	WX6405 = NAND(I19528, I19529)
--	I19534 = NAND(WX5815, CRC_OUT_5_31)
--	I19535 = NAND(WX5815, I19534)
--	I19536 = NAND(CRC_OUT_5_31, I19534)
--	WX6406 = NAND(I19535, I19536)
--	I19541 = NAND(WX5784, CRC_OUT_5_30)
--	I19542 = NAND(WX5784, I19541)
--	I19543 = NAND(CRC_OUT_5_30, I19541)
--	WX6407 = NAND(I19542, I19543)
--	I19548 = NAND(WX5785, CRC_OUT_5_29)
--	I19549 = NAND(WX5785, I19548)
--	I19550 = NAND(CRC_OUT_5_29, I19548)
--	WX6408 = NAND(I19549, I19550)
--	I19555 = NAND(WX5786, CRC_OUT_5_28)
--	I19556 = NAND(WX5786, I19555)
--	I19557 = NAND(CRC_OUT_5_28, I19555)
--	WX6409 = NAND(I19556, I19557)
--	I19562 = NAND(WX5787, CRC_OUT_5_27)
--	I19563 = NAND(WX5787, I19562)
--	I19564 = NAND(CRC_OUT_5_27, I19562)
--	WX6410 = NAND(I19563, I19564)
--	I19569 = NAND(WX5788, CRC_OUT_5_26)
--	I19570 = NAND(WX5788, I19569)
--	I19571 = NAND(CRC_OUT_5_26, I19569)
--	WX6411 = NAND(I19570, I19571)
--	I19576 = NAND(WX5789, CRC_OUT_5_25)
--	I19577 = NAND(WX5789, I19576)
--	I19578 = NAND(CRC_OUT_5_25, I19576)
--	WX6412 = NAND(I19577, I19578)
--	I19583 = NAND(WX5790, CRC_OUT_5_24)
--	I19584 = NAND(WX5790, I19583)
--	I19585 = NAND(CRC_OUT_5_24, I19583)
--	WX6413 = NAND(I19584, I19585)
--	I19590 = NAND(WX5791, CRC_OUT_5_23)
--	I19591 = NAND(WX5791, I19590)
--	I19592 = NAND(CRC_OUT_5_23, I19590)
--	WX6414 = NAND(I19591, I19592)
--	I19597 = NAND(WX5792, CRC_OUT_5_22)
--	I19598 = NAND(WX5792, I19597)
--	I19599 = NAND(CRC_OUT_5_22, I19597)
--	WX6415 = NAND(I19598, I19599)
--	I19604 = NAND(WX5793, CRC_OUT_5_21)
--	I19605 = NAND(WX5793, I19604)
--	I19606 = NAND(CRC_OUT_5_21, I19604)
--	WX6416 = NAND(I19605, I19606)
--	I19611 = NAND(WX5794, CRC_OUT_5_20)
--	I19612 = NAND(WX5794, I19611)
--	I19613 = NAND(CRC_OUT_5_20, I19611)
--	WX6417 = NAND(I19612, I19613)
--	I19618 = NAND(WX5795, CRC_OUT_5_19)
--	I19619 = NAND(WX5795, I19618)
--	I19620 = NAND(CRC_OUT_5_19, I19618)
--	WX6418 = NAND(I19619, I19620)
--	I19625 = NAND(WX5796, CRC_OUT_5_18)
--	I19626 = NAND(WX5796, I19625)
--	I19627 = NAND(CRC_OUT_5_18, I19625)
--	WX6419 = NAND(I19626, I19627)
--	I19632 = NAND(WX5797, CRC_OUT_5_17)
--	I19633 = NAND(WX5797, I19632)
--	I19634 = NAND(CRC_OUT_5_17, I19632)
--	WX6420 = NAND(I19633, I19634)
--	I19639 = NAND(WX5798, CRC_OUT_5_16)
--	I19640 = NAND(WX5798, I19639)
--	I19641 = NAND(CRC_OUT_5_16, I19639)
--	WX6421 = NAND(I19640, I19641)
--	I19646 = NAND(WX5800, CRC_OUT_5_14)
--	I19647 = NAND(WX5800, I19646)
--	I19648 = NAND(CRC_OUT_5_14, I19646)
--	WX6422 = NAND(I19647, I19648)
--	I19653 = NAND(WX5801, CRC_OUT_5_13)
--	I19654 = NAND(WX5801, I19653)
--	I19655 = NAND(CRC_OUT_5_13, I19653)
--	WX6423 = NAND(I19654, I19655)
--	I19660 = NAND(WX5802, CRC_OUT_5_12)
--	I19661 = NAND(WX5802, I19660)
--	I19662 = NAND(CRC_OUT_5_12, I19660)
--	WX6424 = NAND(I19661, I19662)
--	I19667 = NAND(WX5803, CRC_OUT_5_11)
--	I19668 = NAND(WX5803, I19667)
--	I19669 = NAND(CRC_OUT_5_11, I19667)
--	WX6425 = NAND(I19668, I19669)
--	I19674 = NAND(WX5805, CRC_OUT_5_9)
--	I19675 = NAND(WX5805, I19674)
--	I19676 = NAND(CRC_OUT_5_9, I19674)
--	WX6426 = NAND(I19675, I19676)
--	I19681 = NAND(WX5806, CRC_OUT_5_8)
--	I19682 = NAND(WX5806, I19681)
--	I19683 = NAND(CRC_OUT_5_8, I19681)
--	WX6427 = NAND(I19682, I19683)
--	I19688 = NAND(WX5807, CRC_OUT_5_7)
--	I19689 = NAND(WX5807, I19688)
--	I19690 = NAND(CRC_OUT_5_7, I19688)
--	WX6428 = NAND(I19689, I19690)
--	I19695 = NAND(WX5808, CRC_OUT_5_6)
--	I19696 = NAND(WX5808, I19695)
--	I19697 = NAND(CRC_OUT_5_6, I19695)
--	WX6429 = NAND(I19696, I19697)
--	I19702 = NAND(WX5809, CRC_OUT_5_5)
--	I19703 = NAND(WX5809, I19702)
--	I19704 = NAND(CRC_OUT_5_5, I19702)
--	WX6430 = NAND(I19703, I19704)
--	I19709 = NAND(WX5810, CRC_OUT_5_4)
--	I19710 = NAND(WX5810, I19709)
--	I19711 = NAND(CRC_OUT_5_4, I19709)
--	WX6431 = NAND(I19710, I19711)
--	I19716 = NAND(WX5812, CRC_OUT_5_2)
--	I19717 = NAND(WX5812, I19716)
--	I19718 = NAND(CRC_OUT_5_2, I19716)
--	WX6432 = NAND(I19717, I19718)
--	I19723 = NAND(WX5813, CRC_OUT_5_1)
--	I19724 = NAND(WX5813, I19723)
--	I19725 = NAND(CRC_OUT_5_1, I19723)
--	WX6433 = NAND(I19724, I19725)
--	I19730 = NAND(WX5814, CRC_OUT_5_0)
--	I19731 = NAND(WX5814, I19730)
--	I19732 = NAND(CRC_OUT_5_0, I19730)
--	WX6434 = NAND(I19731, I19732)
--	I22013 = NAND(WX7466, WX7110)
--	I22014 = NAND(WX7466, I22013)
--	I22015 = NAND(WX7110, I22013)
--	I22012 = NAND(I22014, I22015)
--	I22020 = NAND(WX7174, I22012)
--	I22021 = NAND(WX7174, I22020)
--	I22022 = NAND(I22012, I22020)
--	I22011 = NAND(I22021, I22022)
--	I22028 = NAND(WX7238, WX7302)
--	I22029 = NAND(WX7238, I22028)
--	I22030 = NAND(WX7302, I22028)
--	I22027 = NAND(I22029, I22030)
--	I22035 = NAND(I22011, I22027)
--	I22036 = NAND(I22011, I22035)
--	I22037 = NAND(I22027, I22035)
--	WX7365 = NAND(I22036, I22037)
--	I22044 = NAND(WX7466, WX7112)
--	I22045 = NAND(WX7466, I22044)
--	I22046 = NAND(WX7112, I22044)
--	I22043 = NAND(I22045, I22046)
--	I22051 = NAND(WX7176, I22043)
--	I22052 = NAND(WX7176, I22051)
--	I22053 = NAND(I22043, I22051)
--	I22042 = NAND(I22052, I22053)
--	I22059 = NAND(WX7240, WX7304)
--	I22060 = NAND(WX7240, I22059)
--	I22061 = NAND(WX7304, I22059)
--	I22058 = NAND(I22060, I22061)
--	I22066 = NAND(I22042, I22058)
--	I22067 = NAND(I22042, I22066)
--	I22068 = NAND(I22058, I22066)
--	WX7366 = NAND(I22067, I22068)
--	I22075 = NAND(WX7466, WX7114)
--	I22076 = NAND(WX7466, I22075)
--	I22077 = NAND(WX7114, I22075)
--	I22074 = NAND(I22076, I22077)
--	I22082 = NAND(WX7178, I22074)
--	I22083 = NAND(WX7178, I22082)
--	I22084 = NAND(I22074, I22082)
--	I22073 = NAND(I22083, I22084)
--	I22090 = NAND(WX7242, WX7306)
--	I22091 = NAND(WX7242, I22090)
--	I22092 = NAND(WX7306, I22090)
--	I22089 = NAND(I22091, I22092)
--	I22097 = NAND(I22073, I22089)
--	I22098 = NAND(I22073, I22097)
--	I22099 = NAND(I22089, I22097)
--	WX7367 = NAND(I22098, I22099)
--	I22106 = NAND(WX7466, WX7116)
--	I22107 = NAND(WX7466, I22106)
--	I22108 = NAND(WX7116, I22106)
--	I22105 = NAND(I22107, I22108)
--	I22113 = NAND(WX7180, I22105)
--	I22114 = NAND(WX7180, I22113)
--	I22115 = NAND(I22105, I22113)
--	I22104 = NAND(I22114, I22115)
--	I22121 = NAND(WX7244, WX7308)
--	I22122 = NAND(WX7244, I22121)
--	I22123 = NAND(WX7308, I22121)
--	I22120 = NAND(I22122, I22123)
--	I22128 = NAND(I22104, I22120)
--	I22129 = NAND(I22104, I22128)
--	I22130 = NAND(I22120, I22128)
--	WX7368 = NAND(I22129, I22130)
--	I22137 = NAND(WX7466, WX7118)
--	I22138 = NAND(WX7466, I22137)
--	I22139 = NAND(WX7118, I22137)
--	I22136 = NAND(I22138, I22139)
--	I22144 = NAND(WX7182, I22136)
--	I22145 = NAND(WX7182, I22144)
--	I22146 = NAND(I22136, I22144)
--	I22135 = NAND(I22145, I22146)
--	I22152 = NAND(WX7246, WX7310)
--	I22153 = NAND(WX7246, I22152)
--	I22154 = NAND(WX7310, I22152)
--	I22151 = NAND(I22153, I22154)
--	I22159 = NAND(I22135, I22151)
--	I22160 = NAND(I22135, I22159)
--	I22161 = NAND(I22151, I22159)
--	WX7369 = NAND(I22160, I22161)
--	I22168 = NAND(WX7466, WX7120)
--	I22169 = NAND(WX7466, I22168)
--	I22170 = NAND(WX7120, I22168)
--	I22167 = NAND(I22169, I22170)
--	I22175 = NAND(WX7184, I22167)
--	I22176 = NAND(WX7184, I22175)
--	I22177 = NAND(I22167, I22175)
--	I22166 = NAND(I22176, I22177)
--	I22183 = NAND(WX7248, WX7312)
--	I22184 = NAND(WX7248, I22183)
--	I22185 = NAND(WX7312, I22183)
--	I22182 = NAND(I22184, I22185)
--	I22190 = NAND(I22166, I22182)
--	I22191 = NAND(I22166, I22190)
--	I22192 = NAND(I22182, I22190)
--	WX7370 = NAND(I22191, I22192)
--	I22199 = NAND(WX7466, WX7122)
--	I22200 = NAND(WX7466, I22199)
--	I22201 = NAND(WX7122, I22199)
--	I22198 = NAND(I22200, I22201)
--	I22206 = NAND(WX7186, I22198)
--	I22207 = NAND(WX7186, I22206)
--	I22208 = NAND(I22198, I22206)
--	I22197 = NAND(I22207, I22208)
--	I22214 = NAND(WX7250, WX7314)
--	I22215 = NAND(WX7250, I22214)
--	I22216 = NAND(WX7314, I22214)
--	I22213 = NAND(I22215, I22216)
--	I22221 = NAND(I22197, I22213)
--	I22222 = NAND(I22197, I22221)
--	I22223 = NAND(I22213, I22221)
--	WX7371 = NAND(I22222, I22223)
--	I22230 = NAND(WX7466, WX7124)
--	I22231 = NAND(WX7466, I22230)
--	I22232 = NAND(WX7124, I22230)
--	I22229 = NAND(I22231, I22232)
--	I22237 = NAND(WX7188, I22229)
--	I22238 = NAND(WX7188, I22237)
--	I22239 = NAND(I22229, I22237)
--	I22228 = NAND(I22238, I22239)
--	I22245 = NAND(WX7252, WX7316)
--	I22246 = NAND(WX7252, I22245)
--	I22247 = NAND(WX7316, I22245)
--	I22244 = NAND(I22246, I22247)
--	I22252 = NAND(I22228, I22244)
--	I22253 = NAND(I22228, I22252)
--	I22254 = NAND(I22244, I22252)
--	WX7372 = NAND(I22253, I22254)
--	I22261 = NAND(WX7466, WX7126)
--	I22262 = NAND(WX7466, I22261)
--	I22263 = NAND(WX7126, I22261)
--	I22260 = NAND(I22262, I22263)
--	I22268 = NAND(WX7190, I22260)
--	I22269 = NAND(WX7190, I22268)
--	I22270 = NAND(I22260, I22268)
--	I22259 = NAND(I22269, I22270)
--	I22276 = NAND(WX7254, WX7318)
--	I22277 = NAND(WX7254, I22276)
--	I22278 = NAND(WX7318, I22276)
--	I22275 = NAND(I22277, I22278)
--	I22283 = NAND(I22259, I22275)
--	I22284 = NAND(I22259, I22283)
--	I22285 = NAND(I22275, I22283)
--	WX7373 = NAND(I22284, I22285)
--	I22292 = NAND(WX7466, WX7128)
--	I22293 = NAND(WX7466, I22292)
--	I22294 = NAND(WX7128, I22292)
--	I22291 = NAND(I22293, I22294)
--	I22299 = NAND(WX7192, I22291)
--	I22300 = NAND(WX7192, I22299)
--	I22301 = NAND(I22291, I22299)
--	I22290 = NAND(I22300, I22301)
--	I22307 = NAND(WX7256, WX7320)
--	I22308 = NAND(WX7256, I22307)
--	I22309 = NAND(WX7320, I22307)
--	I22306 = NAND(I22308, I22309)
--	I22314 = NAND(I22290, I22306)
--	I22315 = NAND(I22290, I22314)
--	I22316 = NAND(I22306, I22314)
--	WX7374 = NAND(I22315, I22316)
--	I22323 = NAND(WX7466, WX7130)
--	I22324 = NAND(WX7466, I22323)
--	I22325 = NAND(WX7130, I22323)
--	I22322 = NAND(I22324, I22325)
--	I22330 = NAND(WX7194, I22322)
--	I22331 = NAND(WX7194, I22330)
--	I22332 = NAND(I22322, I22330)
--	I22321 = NAND(I22331, I22332)
--	I22338 = NAND(WX7258, WX7322)
--	I22339 = NAND(WX7258, I22338)
--	I22340 = NAND(WX7322, I22338)
--	I22337 = NAND(I22339, I22340)
--	I22345 = NAND(I22321, I22337)
--	I22346 = NAND(I22321, I22345)
--	I22347 = NAND(I22337, I22345)
--	WX7375 = NAND(I22346, I22347)
--	I22354 = NAND(WX7466, WX7132)
--	I22355 = NAND(WX7466, I22354)
--	I22356 = NAND(WX7132, I22354)
--	I22353 = NAND(I22355, I22356)
--	I22361 = NAND(WX7196, I22353)
--	I22362 = NAND(WX7196, I22361)
--	I22363 = NAND(I22353, I22361)
--	I22352 = NAND(I22362, I22363)
--	I22369 = NAND(WX7260, WX7324)
--	I22370 = NAND(WX7260, I22369)
--	I22371 = NAND(WX7324, I22369)
--	I22368 = NAND(I22370, I22371)
--	I22376 = NAND(I22352, I22368)
--	I22377 = NAND(I22352, I22376)
--	I22378 = NAND(I22368, I22376)
--	WX7376 = NAND(I22377, I22378)
--	I22385 = NAND(WX7466, WX7134)
--	I22386 = NAND(WX7466, I22385)
--	I22387 = NAND(WX7134, I22385)
--	I22384 = NAND(I22386, I22387)
--	I22392 = NAND(WX7198, I22384)
--	I22393 = NAND(WX7198, I22392)
--	I22394 = NAND(I22384, I22392)
--	I22383 = NAND(I22393, I22394)
--	I22400 = NAND(WX7262, WX7326)
--	I22401 = NAND(WX7262, I22400)
--	I22402 = NAND(WX7326, I22400)
--	I22399 = NAND(I22401, I22402)
--	I22407 = NAND(I22383, I22399)
--	I22408 = NAND(I22383, I22407)
--	I22409 = NAND(I22399, I22407)
--	WX7377 = NAND(I22408, I22409)
--	I22416 = NAND(WX7466, WX7136)
--	I22417 = NAND(WX7466, I22416)
--	I22418 = NAND(WX7136, I22416)
--	I22415 = NAND(I22417, I22418)
--	I22423 = NAND(WX7200, I22415)
--	I22424 = NAND(WX7200, I22423)
--	I22425 = NAND(I22415, I22423)
--	I22414 = NAND(I22424, I22425)
--	I22431 = NAND(WX7264, WX7328)
--	I22432 = NAND(WX7264, I22431)
--	I22433 = NAND(WX7328, I22431)
--	I22430 = NAND(I22432, I22433)
--	I22438 = NAND(I22414, I22430)
--	I22439 = NAND(I22414, I22438)
--	I22440 = NAND(I22430, I22438)
--	WX7378 = NAND(I22439, I22440)
--	I22447 = NAND(WX7466, WX7138)
--	I22448 = NAND(WX7466, I22447)
--	I22449 = NAND(WX7138, I22447)
--	I22446 = NAND(I22448, I22449)
--	I22454 = NAND(WX7202, I22446)
--	I22455 = NAND(WX7202, I22454)
--	I22456 = NAND(I22446, I22454)
--	I22445 = NAND(I22455, I22456)
--	I22462 = NAND(WX7266, WX7330)
--	I22463 = NAND(WX7266, I22462)
--	I22464 = NAND(WX7330, I22462)
--	I22461 = NAND(I22463, I22464)
--	I22469 = NAND(I22445, I22461)
--	I22470 = NAND(I22445, I22469)
--	I22471 = NAND(I22461, I22469)
--	WX7379 = NAND(I22470, I22471)
--	I22478 = NAND(WX7466, WX7140)
--	I22479 = NAND(WX7466, I22478)
--	I22480 = NAND(WX7140, I22478)
--	I22477 = NAND(I22479, I22480)
--	I22485 = NAND(WX7204, I22477)
--	I22486 = NAND(WX7204, I22485)
--	I22487 = NAND(I22477, I22485)
--	I22476 = NAND(I22486, I22487)
--	I22493 = NAND(WX7268, WX7332)
--	I22494 = NAND(WX7268, I22493)
--	I22495 = NAND(WX7332, I22493)
--	I22492 = NAND(I22494, I22495)
--	I22500 = NAND(I22476, I22492)
--	I22501 = NAND(I22476, I22500)
--	I22502 = NAND(I22492, I22500)
--	WX7380 = NAND(I22501, I22502)
--	I22509 = NAND(WX7467, WX7142)
--	I22510 = NAND(WX7467, I22509)
--	I22511 = NAND(WX7142, I22509)
--	I22508 = NAND(I22510, I22511)
--	I22516 = NAND(WX7206, I22508)
--	I22517 = NAND(WX7206, I22516)
--	I22518 = NAND(I22508, I22516)
--	I22507 = NAND(I22517, I22518)
--	I22524 = NAND(WX7270, WX7334)
--	I22525 = NAND(WX7270, I22524)
--	I22526 = NAND(WX7334, I22524)
--	I22523 = NAND(I22525, I22526)
--	I22531 = NAND(I22507, I22523)
--	I22532 = NAND(I22507, I22531)
--	I22533 = NAND(I22523, I22531)
--	WX7381 = NAND(I22532, I22533)
--	I22540 = NAND(WX7467, WX7144)
--	I22541 = NAND(WX7467, I22540)
--	I22542 = NAND(WX7144, I22540)
--	I22539 = NAND(I22541, I22542)
--	I22547 = NAND(WX7208, I22539)
--	I22548 = NAND(WX7208, I22547)
--	I22549 = NAND(I22539, I22547)
--	I22538 = NAND(I22548, I22549)
--	I22555 = NAND(WX7272, WX7336)
--	I22556 = NAND(WX7272, I22555)
--	I22557 = NAND(WX7336, I22555)
--	I22554 = NAND(I22556, I22557)
--	I22562 = NAND(I22538, I22554)
--	I22563 = NAND(I22538, I22562)
--	I22564 = NAND(I22554, I22562)
--	WX7382 = NAND(I22563, I22564)
--	I22571 = NAND(WX7467, WX7146)
--	I22572 = NAND(WX7467, I22571)
--	I22573 = NAND(WX7146, I22571)
--	I22570 = NAND(I22572, I22573)
--	I22578 = NAND(WX7210, I22570)
--	I22579 = NAND(WX7210, I22578)
--	I22580 = NAND(I22570, I22578)
--	I22569 = NAND(I22579, I22580)
--	I22586 = NAND(WX7274, WX7338)
--	I22587 = NAND(WX7274, I22586)
--	I22588 = NAND(WX7338, I22586)
--	I22585 = NAND(I22587, I22588)
--	I22593 = NAND(I22569, I22585)
--	I22594 = NAND(I22569, I22593)
--	I22595 = NAND(I22585, I22593)
--	WX7383 = NAND(I22594, I22595)
--	I22602 = NAND(WX7467, WX7148)
--	I22603 = NAND(WX7467, I22602)
--	I22604 = NAND(WX7148, I22602)
--	I22601 = NAND(I22603, I22604)
--	I22609 = NAND(WX7212, I22601)
--	I22610 = NAND(WX7212, I22609)
--	I22611 = NAND(I22601, I22609)
--	I22600 = NAND(I22610, I22611)
--	I22617 = NAND(WX7276, WX7340)
--	I22618 = NAND(WX7276, I22617)
--	I22619 = NAND(WX7340, I22617)
--	I22616 = NAND(I22618, I22619)
--	I22624 = NAND(I22600, I22616)
--	I22625 = NAND(I22600, I22624)
--	I22626 = NAND(I22616, I22624)
--	WX7384 = NAND(I22625, I22626)
--	I22633 = NAND(WX7467, WX7150)
--	I22634 = NAND(WX7467, I22633)
--	I22635 = NAND(WX7150, I22633)
--	I22632 = NAND(I22634, I22635)
--	I22640 = NAND(WX7214, I22632)
--	I22641 = NAND(WX7214, I22640)
--	I22642 = NAND(I22632, I22640)
--	I22631 = NAND(I22641, I22642)
--	I22648 = NAND(WX7278, WX7342)
--	I22649 = NAND(WX7278, I22648)
--	I22650 = NAND(WX7342, I22648)
--	I22647 = NAND(I22649, I22650)
--	I22655 = NAND(I22631, I22647)
--	I22656 = NAND(I22631, I22655)
--	I22657 = NAND(I22647, I22655)
--	WX7385 = NAND(I22656, I22657)
--	I22664 = NAND(WX7467, WX7152)
--	I22665 = NAND(WX7467, I22664)
--	I22666 = NAND(WX7152, I22664)
--	I22663 = NAND(I22665, I22666)
--	I22671 = NAND(WX7216, I22663)
--	I22672 = NAND(WX7216, I22671)
--	I22673 = NAND(I22663, I22671)
--	I22662 = NAND(I22672, I22673)
--	I22679 = NAND(WX7280, WX7344)
--	I22680 = NAND(WX7280, I22679)
--	I22681 = NAND(WX7344, I22679)
--	I22678 = NAND(I22680, I22681)
--	I22686 = NAND(I22662, I22678)
--	I22687 = NAND(I22662, I22686)
--	I22688 = NAND(I22678, I22686)
--	WX7386 = NAND(I22687, I22688)
--	I22695 = NAND(WX7467, WX7154)
--	I22696 = NAND(WX7467, I22695)
--	I22697 = NAND(WX7154, I22695)
--	I22694 = NAND(I22696, I22697)
--	I22702 = NAND(WX7218, I22694)
--	I22703 = NAND(WX7218, I22702)
--	I22704 = NAND(I22694, I22702)
--	I22693 = NAND(I22703, I22704)
--	I22710 = NAND(WX7282, WX7346)
--	I22711 = NAND(WX7282, I22710)
--	I22712 = NAND(WX7346, I22710)
--	I22709 = NAND(I22711, I22712)
--	I22717 = NAND(I22693, I22709)
--	I22718 = NAND(I22693, I22717)
--	I22719 = NAND(I22709, I22717)
--	WX7387 = NAND(I22718, I22719)
--	I22726 = NAND(WX7467, WX7156)
--	I22727 = NAND(WX7467, I22726)
--	I22728 = NAND(WX7156, I22726)
--	I22725 = NAND(I22727, I22728)
--	I22733 = NAND(WX7220, I22725)
--	I22734 = NAND(WX7220, I22733)
--	I22735 = NAND(I22725, I22733)
--	I22724 = NAND(I22734, I22735)
--	I22741 = NAND(WX7284, WX7348)
--	I22742 = NAND(WX7284, I22741)
--	I22743 = NAND(WX7348, I22741)
--	I22740 = NAND(I22742, I22743)
--	I22748 = NAND(I22724, I22740)
--	I22749 = NAND(I22724, I22748)
--	I22750 = NAND(I22740, I22748)
--	WX7388 = NAND(I22749, I22750)
--	I22757 = NAND(WX7467, WX7158)
--	I22758 = NAND(WX7467, I22757)
--	I22759 = NAND(WX7158, I22757)
--	I22756 = NAND(I22758, I22759)
--	I22764 = NAND(WX7222, I22756)
--	I22765 = NAND(WX7222, I22764)
--	I22766 = NAND(I22756, I22764)
--	I22755 = NAND(I22765, I22766)
--	I22772 = NAND(WX7286, WX7350)
--	I22773 = NAND(WX7286, I22772)
--	I22774 = NAND(WX7350, I22772)
--	I22771 = NAND(I22773, I22774)
--	I22779 = NAND(I22755, I22771)
--	I22780 = NAND(I22755, I22779)
--	I22781 = NAND(I22771, I22779)
--	WX7389 = NAND(I22780, I22781)
--	I22788 = NAND(WX7467, WX7160)
--	I22789 = NAND(WX7467, I22788)
--	I22790 = NAND(WX7160, I22788)
--	I22787 = NAND(I22789, I22790)
--	I22795 = NAND(WX7224, I22787)
--	I22796 = NAND(WX7224, I22795)
--	I22797 = NAND(I22787, I22795)
--	I22786 = NAND(I22796, I22797)
--	I22803 = NAND(WX7288, WX7352)
--	I22804 = NAND(WX7288, I22803)
--	I22805 = NAND(WX7352, I22803)
--	I22802 = NAND(I22804, I22805)
--	I22810 = NAND(I22786, I22802)
--	I22811 = NAND(I22786, I22810)
--	I22812 = NAND(I22802, I22810)
--	WX7390 = NAND(I22811, I22812)
--	I22819 = NAND(WX7467, WX7162)
--	I22820 = NAND(WX7467, I22819)
--	I22821 = NAND(WX7162, I22819)
--	I22818 = NAND(I22820, I22821)
--	I22826 = NAND(WX7226, I22818)
--	I22827 = NAND(WX7226, I22826)
--	I22828 = NAND(I22818, I22826)
--	I22817 = NAND(I22827, I22828)
--	I22834 = NAND(WX7290, WX7354)
--	I22835 = NAND(WX7290, I22834)
--	I22836 = NAND(WX7354, I22834)
--	I22833 = NAND(I22835, I22836)
--	I22841 = NAND(I22817, I22833)
--	I22842 = NAND(I22817, I22841)
--	I22843 = NAND(I22833, I22841)
--	WX7391 = NAND(I22842, I22843)
--	I22850 = NAND(WX7467, WX7164)
--	I22851 = NAND(WX7467, I22850)
--	I22852 = NAND(WX7164, I22850)
--	I22849 = NAND(I22851, I22852)
--	I22857 = NAND(WX7228, I22849)
--	I22858 = NAND(WX7228, I22857)
--	I22859 = NAND(I22849, I22857)
--	I22848 = NAND(I22858, I22859)
--	I22865 = NAND(WX7292, WX7356)
--	I22866 = NAND(WX7292, I22865)
--	I22867 = NAND(WX7356, I22865)
--	I22864 = NAND(I22866, I22867)
--	I22872 = NAND(I22848, I22864)
--	I22873 = NAND(I22848, I22872)
--	I22874 = NAND(I22864, I22872)
--	WX7392 = NAND(I22873, I22874)
--	I22881 = NAND(WX7467, WX7166)
--	I22882 = NAND(WX7467, I22881)
--	I22883 = NAND(WX7166, I22881)
--	I22880 = NAND(I22882, I22883)
--	I22888 = NAND(WX7230, I22880)
--	I22889 = NAND(WX7230, I22888)
--	I22890 = NAND(I22880, I22888)
--	I22879 = NAND(I22889, I22890)
--	I22896 = NAND(WX7294, WX7358)
--	I22897 = NAND(WX7294, I22896)
--	I22898 = NAND(WX7358, I22896)
--	I22895 = NAND(I22897, I22898)
--	I22903 = NAND(I22879, I22895)
--	I22904 = NAND(I22879, I22903)
--	I22905 = NAND(I22895, I22903)
--	WX7393 = NAND(I22904, I22905)
--	I22912 = NAND(WX7467, WX7168)
--	I22913 = NAND(WX7467, I22912)
--	I22914 = NAND(WX7168, I22912)
--	I22911 = NAND(I22913, I22914)
--	I22919 = NAND(WX7232, I22911)
--	I22920 = NAND(WX7232, I22919)
--	I22921 = NAND(I22911, I22919)
--	I22910 = NAND(I22920, I22921)
--	I22927 = NAND(WX7296, WX7360)
--	I22928 = NAND(WX7296, I22927)
--	I22929 = NAND(WX7360, I22927)
--	I22926 = NAND(I22928, I22929)
--	I22934 = NAND(I22910, I22926)
--	I22935 = NAND(I22910, I22934)
--	I22936 = NAND(I22926, I22934)
--	WX7394 = NAND(I22935, I22936)
--	I22943 = NAND(WX7467, WX7170)
--	I22944 = NAND(WX7467, I22943)
--	I22945 = NAND(WX7170, I22943)
--	I22942 = NAND(I22944, I22945)
--	I22950 = NAND(WX7234, I22942)
--	I22951 = NAND(WX7234, I22950)
--	I22952 = NAND(I22942, I22950)
--	I22941 = NAND(I22951, I22952)
--	I22958 = NAND(WX7298, WX7362)
--	I22959 = NAND(WX7298, I22958)
--	I22960 = NAND(WX7362, I22958)
--	I22957 = NAND(I22959, I22960)
--	I22965 = NAND(I22941, I22957)
--	I22966 = NAND(I22941, I22965)
--	I22967 = NAND(I22957, I22965)
--	WX7395 = NAND(I22966, I22967)
--	I22974 = NAND(WX7467, WX7172)
--	I22975 = NAND(WX7467, I22974)
--	I22976 = NAND(WX7172, I22974)
--	I22973 = NAND(I22975, I22976)
--	I22981 = NAND(WX7236, I22973)
--	I22982 = NAND(WX7236, I22981)
--	I22983 = NAND(I22973, I22981)
--	I22972 = NAND(I22982, I22983)
--	I22989 = NAND(WX7300, WX7364)
--	I22990 = NAND(WX7300, I22989)
--	I22991 = NAND(WX7364, I22989)
--	I22988 = NAND(I22990, I22991)
--	I22996 = NAND(I22972, I22988)
--	I22997 = NAND(I22972, I22996)
--	I22998 = NAND(I22988, I22996)
--	WX7396 = NAND(I22997, I22998)
--	I23077 = NAND(WX7045, WX6950)
--	I23078 = NAND(WX7045, I23077)
--	I23079 = NAND(WX6950, I23077)
--	WX7471 = NAND(I23078, I23079)
--	I23090 = NAND(WX7046, WX6952)
--	I23091 = NAND(WX7046, I23090)
--	I23092 = NAND(WX6952, I23090)
--	WX7478 = NAND(I23091, I23092)
--	I23103 = NAND(WX7047, WX6954)
--	I23104 = NAND(WX7047, I23103)
--	I23105 = NAND(WX6954, I23103)
--	WX7485 = NAND(I23104, I23105)
--	I23116 = NAND(WX7048, WX6956)
--	I23117 = NAND(WX7048, I23116)
--	I23118 = NAND(WX6956, I23116)
--	WX7492 = NAND(I23117, I23118)
--	I23129 = NAND(WX7049, WX6958)
--	I23130 = NAND(WX7049, I23129)
--	I23131 = NAND(WX6958, I23129)
--	WX7499 = NAND(I23130, I23131)
--	I23142 = NAND(WX7050, WX6960)
--	I23143 = NAND(WX7050, I23142)
--	I23144 = NAND(WX6960, I23142)
--	WX7506 = NAND(I23143, I23144)
--	I23155 = NAND(WX7051, WX6962)
--	I23156 = NAND(WX7051, I23155)
--	I23157 = NAND(WX6962, I23155)
--	WX7513 = NAND(I23156, I23157)
--	I23168 = NAND(WX7052, WX6964)
--	I23169 = NAND(WX7052, I23168)
--	I23170 = NAND(WX6964, I23168)
--	WX7520 = NAND(I23169, I23170)
--	I23181 = NAND(WX7053, WX6966)
--	I23182 = NAND(WX7053, I23181)
--	I23183 = NAND(WX6966, I23181)
--	WX7527 = NAND(I23182, I23183)
--	I23194 = NAND(WX7054, WX6968)
--	I23195 = NAND(WX7054, I23194)
--	I23196 = NAND(WX6968, I23194)
--	WX7534 = NAND(I23195, I23196)
--	I23207 = NAND(WX7055, WX6970)
--	I23208 = NAND(WX7055, I23207)
--	I23209 = NAND(WX6970, I23207)
--	WX7541 = NAND(I23208, I23209)
--	I23220 = NAND(WX7056, WX6972)
--	I23221 = NAND(WX7056, I23220)
--	I23222 = NAND(WX6972, I23220)
--	WX7548 = NAND(I23221, I23222)
--	I23233 = NAND(WX7057, WX6974)
--	I23234 = NAND(WX7057, I23233)
--	I23235 = NAND(WX6974, I23233)
--	WX7555 = NAND(I23234, I23235)
--	I23246 = NAND(WX7058, WX6976)
--	I23247 = NAND(WX7058, I23246)
--	I23248 = NAND(WX6976, I23246)
--	WX7562 = NAND(I23247, I23248)
--	I23259 = NAND(WX7059, WX6978)
--	I23260 = NAND(WX7059, I23259)
--	I23261 = NAND(WX6978, I23259)
--	WX7569 = NAND(I23260, I23261)
--	I23272 = NAND(WX7060, WX6980)
--	I23273 = NAND(WX7060, I23272)
--	I23274 = NAND(WX6980, I23272)
--	WX7576 = NAND(I23273, I23274)
--	I23285 = NAND(WX7061, WX6982)
--	I23286 = NAND(WX7061, I23285)
--	I23287 = NAND(WX6982, I23285)
--	WX7583 = NAND(I23286, I23287)
--	I23298 = NAND(WX7062, WX6984)
--	I23299 = NAND(WX7062, I23298)
--	I23300 = NAND(WX6984, I23298)
--	WX7590 = NAND(I23299, I23300)
--	I23311 = NAND(WX7063, WX6986)
--	I23312 = NAND(WX7063, I23311)
--	I23313 = NAND(WX6986, I23311)
--	WX7597 = NAND(I23312, I23313)
--	I23324 = NAND(WX7064, WX6988)
--	I23325 = NAND(WX7064, I23324)
--	I23326 = NAND(WX6988, I23324)
--	WX7604 = NAND(I23325, I23326)
--	I23337 = NAND(WX7065, WX6990)
--	I23338 = NAND(WX7065, I23337)
--	I23339 = NAND(WX6990, I23337)
--	WX7611 = NAND(I23338, I23339)
--	I23350 = NAND(WX7066, WX6992)
--	I23351 = NAND(WX7066, I23350)
--	I23352 = NAND(WX6992, I23350)
--	WX7618 = NAND(I23351, I23352)
--	I23363 = NAND(WX7067, WX6994)
--	I23364 = NAND(WX7067, I23363)
--	I23365 = NAND(WX6994, I23363)
--	WX7625 = NAND(I23364, I23365)
--	I23376 = NAND(WX7068, WX6996)
--	I23377 = NAND(WX7068, I23376)
--	I23378 = NAND(WX6996, I23376)
--	WX7632 = NAND(I23377, I23378)
--	I23389 = NAND(WX7069, WX6998)
--	I23390 = NAND(WX7069, I23389)
--	I23391 = NAND(WX6998, I23389)
--	WX7639 = NAND(I23390, I23391)
--	I23402 = NAND(WX7070, WX7000)
--	I23403 = NAND(WX7070, I23402)
--	I23404 = NAND(WX7000, I23402)
--	WX7646 = NAND(I23403, I23404)
--	I23415 = NAND(WX7071, WX7002)
--	I23416 = NAND(WX7071, I23415)
--	I23417 = NAND(WX7002, I23415)
--	WX7653 = NAND(I23416, I23417)
--	I23428 = NAND(WX7072, WX7004)
--	I23429 = NAND(WX7072, I23428)
--	I23430 = NAND(WX7004, I23428)
--	WX7660 = NAND(I23429, I23430)
--	I23441 = NAND(WX7073, WX7006)
--	I23442 = NAND(WX7073, I23441)
--	I23443 = NAND(WX7006, I23441)
--	WX7667 = NAND(I23442, I23443)
--	I23454 = NAND(WX7074, WX7008)
--	I23455 = NAND(WX7074, I23454)
--	I23456 = NAND(WX7008, I23454)
--	WX7674 = NAND(I23455, I23456)
--	I23467 = NAND(WX7075, WX7010)
--	I23468 = NAND(WX7075, I23467)
--	I23469 = NAND(WX7010, I23467)
--	WX7681 = NAND(I23468, I23469)
--	I23480 = NAND(WX7076, WX7012)
--	I23481 = NAND(WX7076, I23480)
--	I23482 = NAND(WX7012, I23480)
--	WX7688 = NAND(I23481, I23482)
--	I23495 = NAND(WX7092, CRC_OUT_4_31)
--	I23496 = NAND(WX7092, I23495)
--	I23497 = NAND(CRC_OUT_4_31, I23495)
--	I23494 = NAND(I23496, I23497)
--	I23502 = NAND(CRC_OUT_4_15, I23494)
--	I23503 = NAND(CRC_OUT_4_15, I23502)
--	I23504 = NAND(I23494, I23502)
--	WX7696 = NAND(I23503, I23504)
--	I23510 = NAND(WX7097, CRC_OUT_4_31)
--	I23511 = NAND(WX7097, I23510)
--	I23512 = NAND(CRC_OUT_4_31, I23510)
--	I23509 = NAND(I23511, I23512)
--	I23517 = NAND(CRC_OUT_4_10, I23509)
--	I23518 = NAND(CRC_OUT_4_10, I23517)
--	I23519 = NAND(I23509, I23517)
--	WX7697 = NAND(I23518, I23519)
--	I23525 = NAND(WX7104, CRC_OUT_4_31)
--	I23526 = NAND(WX7104, I23525)
--	I23527 = NAND(CRC_OUT_4_31, I23525)
--	I23524 = NAND(I23526, I23527)
--	I23532 = NAND(CRC_OUT_4_3, I23524)
--	I23533 = NAND(CRC_OUT_4_3, I23532)
--	I23534 = NAND(I23524, I23532)
--	WX7698 = NAND(I23533, I23534)
--	I23539 = NAND(WX7108, CRC_OUT_4_31)
--	I23540 = NAND(WX7108, I23539)
--	I23541 = NAND(CRC_OUT_4_31, I23539)
--	WX7699 = NAND(I23540, I23541)
--	I23546 = NAND(WX7077, CRC_OUT_4_30)
--	I23547 = NAND(WX7077, I23546)
--	I23548 = NAND(CRC_OUT_4_30, I23546)
--	WX7700 = NAND(I23547, I23548)
--	I23553 = NAND(WX7078, CRC_OUT_4_29)
--	I23554 = NAND(WX7078, I23553)
--	I23555 = NAND(CRC_OUT_4_29, I23553)
--	WX7701 = NAND(I23554, I23555)
--	I23560 = NAND(WX7079, CRC_OUT_4_28)
--	I23561 = NAND(WX7079, I23560)
--	I23562 = NAND(CRC_OUT_4_28, I23560)
--	WX7702 = NAND(I23561, I23562)
--	I23567 = NAND(WX7080, CRC_OUT_4_27)
--	I23568 = NAND(WX7080, I23567)
--	I23569 = NAND(CRC_OUT_4_27, I23567)
--	WX7703 = NAND(I23568, I23569)
--	I23574 = NAND(WX7081, CRC_OUT_4_26)
--	I23575 = NAND(WX7081, I23574)
--	I23576 = NAND(CRC_OUT_4_26, I23574)
--	WX7704 = NAND(I23575, I23576)
--	I23581 = NAND(WX7082, CRC_OUT_4_25)
--	I23582 = NAND(WX7082, I23581)
--	I23583 = NAND(CRC_OUT_4_25, I23581)
--	WX7705 = NAND(I23582, I23583)
--	I23588 = NAND(WX7083, CRC_OUT_4_24)
--	I23589 = NAND(WX7083, I23588)
--	I23590 = NAND(CRC_OUT_4_24, I23588)
--	WX7706 = NAND(I23589, I23590)
--	I23595 = NAND(WX7084, CRC_OUT_4_23)
--	I23596 = NAND(WX7084, I23595)
--	I23597 = NAND(CRC_OUT_4_23, I23595)
--	WX7707 = NAND(I23596, I23597)
--	I23602 = NAND(WX7085, CRC_OUT_4_22)
--	I23603 = NAND(WX7085, I23602)
--	I23604 = NAND(CRC_OUT_4_22, I23602)
--	WX7708 = NAND(I23603, I23604)
--	I23609 = NAND(WX7086, CRC_OUT_4_21)
--	I23610 = NAND(WX7086, I23609)
--	I23611 = NAND(CRC_OUT_4_21, I23609)
--	WX7709 = NAND(I23610, I23611)
--	I23616 = NAND(WX7087, CRC_OUT_4_20)
--	I23617 = NAND(WX7087, I23616)
--	I23618 = NAND(CRC_OUT_4_20, I23616)
--	WX7710 = NAND(I23617, I23618)
--	I23623 = NAND(WX7088, CRC_OUT_4_19)
--	I23624 = NAND(WX7088, I23623)
--	I23625 = NAND(CRC_OUT_4_19, I23623)
--	WX7711 = NAND(I23624, I23625)
--	I23630 = NAND(WX7089, CRC_OUT_4_18)
--	I23631 = NAND(WX7089, I23630)
--	I23632 = NAND(CRC_OUT_4_18, I23630)
--	WX7712 = NAND(I23631, I23632)
--	I23637 = NAND(WX7090, CRC_OUT_4_17)
--	I23638 = NAND(WX7090, I23637)
--	I23639 = NAND(CRC_OUT_4_17, I23637)
--	WX7713 = NAND(I23638, I23639)
--	I23644 = NAND(WX7091, CRC_OUT_4_16)
--	I23645 = NAND(WX7091, I23644)
--	I23646 = NAND(CRC_OUT_4_16, I23644)
--	WX7714 = NAND(I23645, I23646)
--	I23651 = NAND(WX7093, CRC_OUT_4_14)
--	I23652 = NAND(WX7093, I23651)
--	I23653 = NAND(CRC_OUT_4_14, I23651)
--	WX7715 = NAND(I23652, I23653)
--	I23658 = NAND(WX7094, CRC_OUT_4_13)
--	I23659 = NAND(WX7094, I23658)
--	I23660 = NAND(CRC_OUT_4_13, I23658)
--	WX7716 = NAND(I23659, I23660)
--	I23665 = NAND(WX7095, CRC_OUT_4_12)
--	I23666 = NAND(WX7095, I23665)
--	I23667 = NAND(CRC_OUT_4_12, I23665)
--	WX7717 = NAND(I23666, I23667)
--	I23672 = NAND(WX7096, CRC_OUT_4_11)
--	I23673 = NAND(WX7096, I23672)
--	I23674 = NAND(CRC_OUT_4_11, I23672)
--	WX7718 = NAND(I23673, I23674)
--	I23679 = NAND(WX7098, CRC_OUT_4_9)
--	I23680 = NAND(WX7098, I23679)
--	I23681 = NAND(CRC_OUT_4_9, I23679)
--	WX7719 = NAND(I23680, I23681)
--	I23686 = NAND(WX7099, CRC_OUT_4_8)
--	I23687 = NAND(WX7099, I23686)
--	I23688 = NAND(CRC_OUT_4_8, I23686)
--	WX7720 = NAND(I23687, I23688)
--	I23693 = NAND(WX7100, CRC_OUT_4_7)
--	I23694 = NAND(WX7100, I23693)
--	I23695 = NAND(CRC_OUT_4_7, I23693)
--	WX7721 = NAND(I23694, I23695)
--	I23700 = NAND(WX7101, CRC_OUT_4_6)
--	I23701 = NAND(WX7101, I23700)
--	I23702 = NAND(CRC_OUT_4_6, I23700)
--	WX7722 = NAND(I23701, I23702)
--	I23707 = NAND(WX7102, CRC_OUT_4_5)
--	I23708 = NAND(WX7102, I23707)
--	I23709 = NAND(CRC_OUT_4_5, I23707)
--	WX7723 = NAND(I23708, I23709)
--	I23714 = NAND(WX7103, CRC_OUT_4_4)
--	I23715 = NAND(WX7103, I23714)
--	I23716 = NAND(CRC_OUT_4_4, I23714)
--	WX7724 = NAND(I23715, I23716)
--	I23721 = NAND(WX7105, CRC_OUT_4_2)
--	I23722 = NAND(WX7105, I23721)
--	I23723 = NAND(CRC_OUT_4_2, I23721)
--	WX7725 = NAND(I23722, I23723)
--	I23728 = NAND(WX7106, CRC_OUT_4_1)
--	I23729 = NAND(WX7106, I23728)
--	I23730 = NAND(CRC_OUT_4_1, I23728)
--	WX7726 = NAND(I23729, I23730)
--	I23735 = NAND(WX7107, CRC_OUT_4_0)
--	I23736 = NAND(WX7107, I23735)
--	I23737 = NAND(CRC_OUT_4_0, I23735)
--	WX7727 = NAND(I23736, I23737)
--	I26018 = NAND(WX8759, WX8403)
--	I26019 = NAND(WX8759, I26018)
--	I26020 = NAND(WX8403, I26018)
--	I26017 = NAND(I26019, I26020)
--	I26025 = NAND(WX8467, I26017)
--	I26026 = NAND(WX8467, I26025)
--	I26027 = NAND(I26017, I26025)
--	I26016 = NAND(I26026, I26027)
--	I26033 = NAND(WX8531, WX8595)
--	I26034 = NAND(WX8531, I26033)
--	I26035 = NAND(WX8595, I26033)
--	I26032 = NAND(I26034, I26035)
--	I26040 = NAND(I26016, I26032)
--	I26041 = NAND(I26016, I26040)
--	I26042 = NAND(I26032, I26040)
--	WX8658 = NAND(I26041, I26042)
--	I26049 = NAND(WX8759, WX8405)
--	I26050 = NAND(WX8759, I26049)
--	I26051 = NAND(WX8405, I26049)
--	I26048 = NAND(I26050, I26051)
--	I26056 = NAND(WX8469, I26048)
--	I26057 = NAND(WX8469, I26056)
--	I26058 = NAND(I26048, I26056)
--	I26047 = NAND(I26057, I26058)
--	I26064 = NAND(WX8533, WX8597)
--	I26065 = NAND(WX8533, I26064)
--	I26066 = NAND(WX8597, I26064)
--	I26063 = NAND(I26065, I26066)
--	I26071 = NAND(I26047, I26063)
--	I26072 = NAND(I26047, I26071)
--	I26073 = NAND(I26063, I26071)
--	WX8659 = NAND(I26072, I26073)
--	I26080 = NAND(WX8759, WX8407)
--	I26081 = NAND(WX8759, I26080)
--	I26082 = NAND(WX8407, I26080)
--	I26079 = NAND(I26081, I26082)
--	I26087 = NAND(WX8471, I26079)
--	I26088 = NAND(WX8471, I26087)
--	I26089 = NAND(I26079, I26087)
--	I26078 = NAND(I26088, I26089)
--	I26095 = NAND(WX8535, WX8599)
--	I26096 = NAND(WX8535, I26095)
--	I26097 = NAND(WX8599, I26095)
--	I26094 = NAND(I26096, I26097)
--	I26102 = NAND(I26078, I26094)
--	I26103 = NAND(I26078, I26102)
--	I26104 = NAND(I26094, I26102)
--	WX8660 = NAND(I26103, I26104)
--	I26111 = NAND(WX8759, WX8409)
--	I26112 = NAND(WX8759, I26111)
--	I26113 = NAND(WX8409, I26111)
--	I26110 = NAND(I26112, I26113)
--	I26118 = NAND(WX8473, I26110)
--	I26119 = NAND(WX8473, I26118)
--	I26120 = NAND(I26110, I26118)
--	I26109 = NAND(I26119, I26120)
--	I26126 = NAND(WX8537, WX8601)
--	I26127 = NAND(WX8537, I26126)
--	I26128 = NAND(WX8601, I26126)
--	I26125 = NAND(I26127, I26128)
--	I26133 = NAND(I26109, I26125)
--	I26134 = NAND(I26109, I26133)
--	I26135 = NAND(I26125, I26133)
--	WX8661 = NAND(I26134, I26135)
--	I26142 = NAND(WX8759, WX8411)
--	I26143 = NAND(WX8759, I26142)
--	I26144 = NAND(WX8411, I26142)
--	I26141 = NAND(I26143, I26144)
--	I26149 = NAND(WX8475, I26141)
--	I26150 = NAND(WX8475, I26149)
--	I26151 = NAND(I26141, I26149)
--	I26140 = NAND(I26150, I26151)
--	I26157 = NAND(WX8539, WX8603)
--	I26158 = NAND(WX8539, I26157)
--	I26159 = NAND(WX8603, I26157)
--	I26156 = NAND(I26158, I26159)
--	I26164 = NAND(I26140, I26156)
--	I26165 = NAND(I26140, I26164)
--	I26166 = NAND(I26156, I26164)
--	WX8662 = NAND(I26165, I26166)
--	I26173 = NAND(WX8759, WX8413)
--	I26174 = NAND(WX8759, I26173)
--	I26175 = NAND(WX8413, I26173)
--	I26172 = NAND(I26174, I26175)
--	I26180 = NAND(WX8477, I26172)
--	I26181 = NAND(WX8477, I26180)
--	I26182 = NAND(I26172, I26180)
--	I26171 = NAND(I26181, I26182)
--	I26188 = NAND(WX8541, WX8605)
--	I26189 = NAND(WX8541, I26188)
--	I26190 = NAND(WX8605, I26188)
--	I26187 = NAND(I26189, I26190)
--	I26195 = NAND(I26171, I26187)
--	I26196 = NAND(I26171, I26195)
--	I26197 = NAND(I26187, I26195)
--	WX8663 = NAND(I26196, I26197)
--	I26204 = NAND(WX8759, WX8415)
--	I26205 = NAND(WX8759, I26204)
--	I26206 = NAND(WX8415, I26204)
--	I26203 = NAND(I26205, I26206)
--	I26211 = NAND(WX8479, I26203)
--	I26212 = NAND(WX8479, I26211)
--	I26213 = NAND(I26203, I26211)
--	I26202 = NAND(I26212, I26213)
--	I26219 = NAND(WX8543, WX8607)
--	I26220 = NAND(WX8543, I26219)
--	I26221 = NAND(WX8607, I26219)
--	I26218 = NAND(I26220, I26221)
--	I26226 = NAND(I26202, I26218)
--	I26227 = NAND(I26202, I26226)
--	I26228 = NAND(I26218, I26226)
--	WX8664 = NAND(I26227, I26228)
--	I26235 = NAND(WX8759, WX8417)
--	I26236 = NAND(WX8759, I26235)
--	I26237 = NAND(WX8417, I26235)
--	I26234 = NAND(I26236, I26237)
--	I26242 = NAND(WX8481, I26234)
--	I26243 = NAND(WX8481, I26242)
--	I26244 = NAND(I26234, I26242)
--	I26233 = NAND(I26243, I26244)
--	I26250 = NAND(WX8545, WX8609)
--	I26251 = NAND(WX8545, I26250)
--	I26252 = NAND(WX8609, I26250)
--	I26249 = NAND(I26251, I26252)
--	I26257 = NAND(I26233, I26249)
--	I26258 = NAND(I26233, I26257)
--	I26259 = NAND(I26249, I26257)
--	WX8665 = NAND(I26258, I26259)
--	I26266 = NAND(WX8759, WX8419)
--	I26267 = NAND(WX8759, I26266)
--	I26268 = NAND(WX8419, I26266)
--	I26265 = NAND(I26267, I26268)
--	I26273 = NAND(WX8483, I26265)
--	I26274 = NAND(WX8483, I26273)
--	I26275 = NAND(I26265, I26273)
--	I26264 = NAND(I26274, I26275)
--	I26281 = NAND(WX8547, WX8611)
--	I26282 = NAND(WX8547, I26281)
--	I26283 = NAND(WX8611, I26281)
--	I26280 = NAND(I26282, I26283)
--	I26288 = NAND(I26264, I26280)
--	I26289 = NAND(I26264, I26288)
--	I26290 = NAND(I26280, I26288)
--	WX8666 = NAND(I26289, I26290)
--	I26297 = NAND(WX8759, WX8421)
--	I26298 = NAND(WX8759, I26297)
--	I26299 = NAND(WX8421, I26297)
--	I26296 = NAND(I26298, I26299)
--	I26304 = NAND(WX8485, I26296)
--	I26305 = NAND(WX8485, I26304)
--	I26306 = NAND(I26296, I26304)
--	I26295 = NAND(I26305, I26306)
--	I26312 = NAND(WX8549, WX8613)
--	I26313 = NAND(WX8549, I26312)
--	I26314 = NAND(WX8613, I26312)
--	I26311 = NAND(I26313, I26314)
--	I26319 = NAND(I26295, I26311)
--	I26320 = NAND(I26295, I26319)
--	I26321 = NAND(I26311, I26319)
--	WX8667 = NAND(I26320, I26321)
--	I26328 = NAND(WX8759, WX8423)
--	I26329 = NAND(WX8759, I26328)
--	I26330 = NAND(WX8423, I26328)
--	I26327 = NAND(I26329, I26330)
--	I26335 = NAND(WX8487, I26327)
--	I26336 = NAND(WX8487, I26335)
--	I26337 = NAND(I26327, I26335)
--	I26326 = NAND(I26336, I26337)
--	I26343 = NAND(WX8551, WX8615)
--	I26344 = NAND(WX8551, I26343)
--	I26345 = NAND(WX8615, I26343)
--	I26342 = NAND(I26344, I26345)
--	I26350 = NAND(I26326, I26342)
--	I26351 = NAND(I26326, I26350)
--	I26352 = NAND(I26342, I26350)
--	WX8668 = NAND(I26351, I26352)
--	I26359 = NAND(WX8759, WX8425)
--	I26360 = NAND(WX8759, I26359)
--	I26361 = NAND(WX8425, I26359)
--	I26358 = NAND(I26360, I26361)
--	I26366 = NAND(WX8489, I26358)
--	I26367 = NAND(WX8489, I26366)
--	I26368 = NAND(I26358, I26366)
--	I26357 = NAND(I26367, I26368)
--	I26374 = NAND(WX8553, WX8617)
--	I26375 = NAND(WX8553, I26374)
--	I26376 = NAND(WX8617, I26374)
--	I26373 = NAND(I26375, I26376)
--	I26381 = NAND(I26357, I26373)
--	I26382 = NAND(I26357, I26381)
--	I26383 = NAND(I26373, I26381)
--	WX8669 = NAND(I26382, I26383)
--	I26390 = NAND(WX8759, WX8427)
--	I26391 = NAND(WX8759, I26390)
--	I26392 = NAND(WX8427, I26390)
--	I26389 = NAND(I26391, I26392)
--	I26397 = NAND(WX8491, I26389)
--	I26398 = NAND(WX8491, I26397)
--	I26399 = NAND(I26389, I26397)
--	I26388 = NAND(I26398, I26399)
--	I26405 = NAND(WX8555, WX8619)
--	I26406 = NAND(WX8555, I26405)
--	I26407 = NAND(WX8619, I26405)
--	I26404 = NAND(I26406, I26407)
--	I26412 = NAND(I26388, I26404)
--	I26413 = NAND(I26388, I26412)
--	I26414 = NAND(I26404, I26412)
--	WX8670 = NAND(I26413, I26414)
--	I26421 = NAND(WX8759, WX8429)
--	I26422 = NAND(WX8759, I26421)
--	I26423 = NAND(WX8429, I26421)
--	I26420 = NAND(I26422, I26423)
--	I26428 = NAND(WX8493, I26420)
--	I26429 = NAND(WX8493, I26428)
--	I26430 = NAND(I26420, I26428)
--	I26419 = NAND(I26429, I26430)
--	I26436 = NAND(WX8557, WX8621)
--	I26437 = NAND(WX8557, I26436)
--	I26438 = NAND(WX8621, I26436)
--	I26435 = NAND(I26437, I26438)
--	I26443 = NAND(I26419, I26435)
--	I26444 = NAND(I26419, I26443)
--	I26445 = NAND(I26435, I26443)
--	WX8671 = NAND(I26444, I26445)
--	I26452 = NAND(WX8759, WX8431)
--	I26453 = NAND(WX8759, I26452)
--	I26454 = NAND(WX8431, I26452)
--	I26451 = NAND(I26453, I26454)
--	I26459 = NAND(WX8495, I26451)
--	I26460 = NAND(WX8495, I26459)
--	I26461 = NAND(I26451, I26459)
--	I26450 = NAND(I26460, I26461)
--	I26467 = NAND(WX8559, WX8623)
--	I26468 = NAND(WX8559, I26467)
--	I26469 = NAND(WX8623, I26467)
--	I26466 = NAND(I26468, I26469)
--	I26474 = NAND(I26450, I26466)
--	I26475 = NAND(I26450, I26474)
--	I26476 = NAND(I26466, I26474)
--	WX8672 = NAND(I26475, I26476)
--	I26483 = NAND(WX8759, WX8433)
--	I26484 = NAND(WX8759, I26483)
--	I26485 = NAND(WX8433, I26483)
--	I26482 = NAND(I26484, I26485)
--	I26490 = NAND(WX8497, I26482)
--	I26491 = NAND(WX8497, I26490)
--	I26492 = NAND(I26482, I26490)
--	I26481 = NAND(I26491, I26492)
--	I26498 = NAND(WX8561, WX8625)
--	I26499 = NAND(WX8561, I26498)
--	I26500 = NAND(WX8625, I26498)
--	I26497 = NAND(I26499, I26500)
--	I26505 = NAND(I26481, I26497)
--	I26506 = NAND(I26481, I26505)
--	I26507 = NAND(I26497, I26505)
--	WX8673 = NAND(I26506, I26507)
--	I26514 = NAND(WX8760, WX8435)
--	I26515 = NAND(WX8760, I26514)
--	I26516 = NAND(WX8435, I26514)
--	I26513 = NAND(I26515, I26516)
--	I26521 = NAND(WX8499, I26513)
--	I26522 = NAND(WX8499, I26521)
--	I26523 = NAND(I26513, I26521)
--	I26512 = NAND(I26522, I26523)
--	I26529 = NAND(WX8563, WX8627)
--	I26530 = NAND(WX8563, I26529)
--	I26531 = NAND(WX8627, I26529)
--	I26528 = NAND(I26530, I26531)
--	I26536 = NAND(I26512, I26528)
--	I26537 = NAND(I26512, I26536)
--	I26538 = NAND(I26528, I26536)
--	WX8674 = NAND(I26537, I26538)
--	I26545 = NAND(WX8760, WX8437)
--	I26546 = NAND(WX8760, I26545)
--	I26547 = NAND(WX8437, I26545)
--	I26544 = NAND(I26546, I26547)
--	I26552 = NAND(WX8501, I26544)
--	I26553 = NAND(WX8501, I26552)
--	I26554 = NAND(I26544, I26552)
--	I26543 = NAND(I26553, I26554)
--	I26560 = NAND(WX8565, WX8629)
--	I26561 = NAND(WX8565, I26560)
--	I26562 = NAND(WX8629, I26560)
--	I26559 = NAND(I26561, I26562)
--	I26567 = NAND(I26543, I26559)
--	I26568 = NAND(I26543, I26567)
--	I26569 = NAND(I26559, I26567)
--	WX8675 = NAND(I26568, I26569)
--	I26576 = NAND(WX8760, WX8439)
--	I26577 = NAND(WX8760, I26576)
--	I26578 = NAND(WX8439, I26576)
--	I26575 = NAND(I26577, I26578)
--	I26583 = NAND(WX8503, I26575)
--	I26584 = NAND(WX8503, I26583)
--	I26585 = NAND(I26575, I26583)
--	I26574 = NAND(I26584, I26585)
--	I26591 = NAND(WX8567, WX8631)
--	I26592 = NAND(WX8567, I26591)
--	I26593 = NAND(WX8631, I26591)
--	I26590 = NAND(I26592, I26593)
--	I26598 = NAND(I26574, I26590)
--	I26599 = NAND(I26574, I26598)
--	I26600 = NAND(I26590, I26598)
--	WX8676 = NAND(I26599, I26600)
--	I26607 = NAND(WX8760, WX8441)
--	I26608 = NAND(WX8760, I26607)
--	I26609 = NAND(WX8441, I26607)
--	I26606 = NAND(I26608, I26609)
--	I26614 = NAND(WX8505, I26606)
--	I26615 = NAND(WX8505, I26614)
--	I26616 = NAND(I26606, I26614)
--	I26605 = NAND(I26615, I26616)
--	I26622 = NAND(WX8569, WX8633)
--	I26623 = NAND(WX8569, I26622)
--	I26624 = NAND(WX8633, I26622)
--	I26621 = NAND(I26623, I26624)
--	I26629 = NAND(I26605, I26621)
--	I26630 = NAND(I26605, I26629)
--	I26631 = NAND(I26621, I26629)
--	WX8677 = NAND(I26630, I26631)
--	I26638 = NAND(WX8760, WX8443)
--	I26639 = NAND(WX8760, I26638)
--	I26640 = NAND(WX8443, I26638)
--	I26637 = NAND(I26639, I26640)
--	I26645 = NAND(WX8507, I26637)
--	I26646 = NAND(WX8507, I26645)
--	I26647 = NAND(I26637, I26645)
--	I26636 = NAND(I26646, I26647)
--	I26653 = NAND(WX8571, WX8635)
--	I26654 = NAND(WX8571, I26653)
--	I26655 = NAND(WX8635, I26653)
--	I26652 = NAND(I26654, I26655)
--	I26660 = NAND(I26636, I26652)
--	I26661 = NAND(I26636, I26660)
--	I26662 = NAND(I26652, I26660)
--	WX8678 = NAND(I26661, I26662)
--	I26669 = NAND(WX8760, WX8445)
--	I26670 = NAND(WX8760, I26669)
--	I26671 = NAND(WX8445, I26669)
--	I26668 = NAND(I26670, I26671)
--	I26676 = NAND(WX8509, I26668)
--	I26677 = NAND(WX8509, I26676)
--	I26678 = NAND(I26668, I26676)
--	I26667 = NAND(I26677, I26678)
--	I26684 = NAND(WX8573, WX8637)
--	I26685 = NAND(WX8573, I26684)
--	I26686 = NAND(WX8637, I26684)
--	I26683 = NAND(I26685, I26686)
--	I26691 = NAND(I26667, I26683)
--	I26692 = NAND(I26667, I26691)
--	I26693 = NAND(I26683, I26691)
--	WX8679 = NAND(I26692, I26693)
--	I26700 = NAND(WX8760, WX8447)
--	I26701 = NAND(WX8760, I26700)
--	I26702 = NAND(WX8447, I26700)
--	I26699 = NAND(I26701, I26702)
--	I26707 = NAND(WX8511, I26699)
--	I26708 = NAND(WX8511, I26707)
--	I26709 = NAND(I26699, I26707)
--	I26698 = NAND(I26708, I26709)
--	I26715 = NAND(WX8575, WX8639)
--	I26716 = NAND(WX8575, I26715)
--	I26717 = NAND(WX8639, I26715)
--	I26714 = NAND(I26716, I26717)
--	I26722 = NAND(I26698, I26714)
--	I26723 = NAND(I26698, I26722)
--	I26724 = NAND(I26714, I26722)
--	WX8680 = NAND(I26723, I26724)
--	I26731 = NAND(WX8760, WX8449)
--	I26732 = NAND(WX8760, I26731)
--	I26733 = NAND(WX8449, I26731)
--	I26730 = NAND(I26732, I26733)
--	I26738 = NAND(WX8513, I26730)
--	I26739 = NAND(WX8513, I26738)
--	I26740 = NAND(I26730, I26738)
--	I26729 = NAND(I26739, I26740)
--	I26746 = NAND(WX8577, WX8641)
--	I26747 = NAND(WX8577, I26746)
--	I26748 = NAND(WX8641, I26746)
--	I26745 = NAND(I26747, I26748)
--	I26753 = NAND(I26729, I26745)
--	I26754 = NAND(I26729, I26753)
--	I26755 = NAND(I26745, I26753)
--	WX8681 = NAND(I26754, I26755)
--	I26762 = NAND(WX8760, WX8451)
--	I26763 = NAND(WX8760, I26762)
--	I26764 = NAND(WX8451, I26762)
--	I26761 = NAND(I26763, I26764)
--	I26769 = NAND(WX8515, I26761)
--	I26770 = NAND(WX8515, I26769)
--	I26771 = NAND(I26761, I26769)
--	I26760 = NAND(I26770, I26771)
--	I26777 = NAND(WX8579, WX8643)
--	I26778 = NAND(WX8579, I26777)
--	I26779 = NAND(WX8643, I26777)
--	I26776 = NAND(I26778, I26779)
--	I26784 = NAND(I26760, I26776)
--	I26785 = NAND(I26760, I26784)
--	I26786 = NAND(I26776, I26784)
--	WX8682 = NAND(I26785, I26786)
--	I26793 = NAND(WX8760, WX8453)
--	I26794 = NAND(WX8760, I26793)
--	I26795 = NAND(WX8453, I26793)
--	I26792 = NAND(I26794, I26795)
--	I26800 = NAND(WX8517, I26792)
--	I26801 = NAND(WX8517, I26800)
--	I26802 = NAND(I26792, I26800)
--	I26791 = NAND(I26801, I26802)
--	I26808 = NAND(WX8581, WX8645)
--	I26809 = NAND(WX8581, I26808)
--	I26810 = NAND(WX8645, I26808)
--	I26807 = NAND(I26809, I26810)
--	I26815 = NAND(I26791, I26807)
--	I26816 = NAND(I26791, I26815)
--	I26817 = NAND(I26807, I26815)
--	WX8683 = NAND(I26816, I26817)
--	I26824 = NAND(WX8760, WX8455)
--	I26825 = NAND(WX8760, I26824)
--	I26826 = NAND(WX8455, I26824)
--	I26823 = NAND(I26825, I26826)
--	I26831 = NAND(WX8519, I26823)
--	I26832 = NAND(WX8519, I26831)
--	I26833 = NAND(I26823, I26831)
--	I26822 = NAND(I26832, I26833)
--	I26839 = NAND(WX8583, WX8647)
--	I26840 = NAND(WX8583, I26839)
--	I26841 = NAND(WX8647, I26839)
--	I26838 = NAND(I26840, I26841)
--	I26846 = NAND(I26822, I26838)
--	I26847 = NAND(I26822, I26846)
--	I26848 = NAND(I26838, I26846)
--	WX8684 = NAND(I26847, I26848)
--	I26855 = NAND(WX8760, WX8457)
--	I26856 = NAND(WX8760, I26855)
--	I26857 = NAND(WX8457, I26855)
--	I26854 = NAND(I26856, I26857)
--	I26862 = NAND(WX8521, I26854)
--	I26863 = NAND(WX8521, I26862)
--	I26864 = NAND(I26854, I26862)
--	I26853 = NAND(I26863, I26864)
--	I26870 = NAND(WX8585, WX8649)
--	I26871 = NAND(WX8585, I26870)
--	I26872 = NAND(WX8649, I26870)
--	I26869 = NAND(I26871, I26872)
--	I26877 = NAND(I26853, I26869)
--	I26878 = NAND(I26853, I26877)
--	I26879 = NAND(I26869, I26877)
--	WX8685 = NAND(I26878, I26879)
--	I26886 = NAND(WX8760, WX8459)
--	I26887 = NAND(WX8760, I26886)
--	I26888 = NAND(WX8459, I26886)
--	I26885 = NAND(I26887, I26888)
--	I26893 = NAND(WX8523, I26885)
--	I26894 = NAND(WX8523, I26893)
--	I26895 = NAND(I26885, I26893)
--	I26884 = NAND(I26894, I26895)
--	I26901 = NAND(WX8587, WX8651)
--	I26902 = NAND(WX8587, I26901)
--	I26903 = NAND(WX8651, I26901)
--	I26900 = NAND(I26902, I26903)
--	I26908 = NAND(I26884, I26900)
--	I26909 = NAND(I26884, I26908)
--	I26910 = NAND(I26900, I26908)
--	WX8686 = NAND(I26909, I26910)
--	I26917 = NAND(WX8760, WX8461)
--	I26918 = NAND(WX8760, I26917)
--	I26919 = NAND(WX8461, I26917)
--	I26916 = NAND(I26918, I26919)
--	I26924 = NAND(WX8525, I26916)
--	I26925 = NAND(WX8525, I26924)
--	I26926 = NAND(I26916, I26924)
--	I26915 = NAND(I26925, I26926)
--	I26932 = NAND(WX8589, WX8653)
--	I26933 = NAND(WX8589, I26932)
--	I26934 = NAND(WX8653, I26932)
--	I26931 = NAND(I26933, I26934)
--	I26939 = NAND(I26915, I26931)
--	I26940 = NAND(I26915, I26939)
--	I26941 = NAND(I26931, I26939)
--	WX8687 = NAND(I26940, I26941)
--	I26948 = NAND(WX8760, WX8463)
--	I26949 = NAND(WX8760, I26948)
--	I26950 = NAND(WX8463, I26948)
--	I26947 = NAND(I26949, I26950)
--	I26955 = NAND(WX8527, I26947)
--	I26956 = NAND(WX8527, I26955)
--	I26957 = NAND(I26947, I26955)
--	I26946 = NAND(I26956, I26957)
--	I26963 = NAND(WX8591, WX8655)
--	I26964 = NAND(WX8591, I26963)
--	I26965 = NAND(WX8655, I26963)
--	I26962 = NAND(I26964, I26965)
--	I26970 = NAND(I26946, I26962)
--	I26971 = NAND(I26946, I26970)
--	I26972 = NAND(I26962, I26970)
--	WX8688 = NAND(I26971, I26972)
--	I26979 = NAND(WX8760, WX8465)
--	I26980 = NAND(WX8760, I26979)
--	I26981 = NAND(WX8465, I26979)
--	I26978 = NAND(I26980, I26981)
--	I26986 = NAND(WX8529, I26978)
--	I26987 = NAND(WX8529, I26986)
--	I26988 = NAND(I26978, I26986)
--	I26977 = NAND(I26987, I26988)
--	I26994 = NAND(WX8593, WX8657)
--	I26995 = NAND(WX8593, I26994)
--	I26996 = NAND(WX8657, I26994)
--	I26993 = NAND(I26995, I26996)
--	I27001 = NAND(I26977, I26993)
--	I27002 = NAND(I26977, I27001)
--	I27003 = NAND(I26993, I27001)
--	WX8689 = NAND(I27002, I27003)
--	I27082 = NAND(WX8338, WX8243)
--	I27083 = NAND(WX8338, I27082)
--	I27084 = NAND(WX8243, I27082)
--	WX8764 = NAND(I27083, I27084)
--	I27095 = NAND(WX8339, WX8245)
--	I27096 = NAND(WX8339, I27095)
--	I27097 = NAND(WX8245, I27095)
--	WX8771 = NAND(I27096, I27097)
--	I27108 = NAND(WX8340, WX8247)
--	I27109 = NAND(WX8340, I27108)
--	I27110 = NAND(WX8247, I27108)
--	WX8778 = NAND(I27109, I27110)
--	I27121 = NAND(WX8341, WX8249)
--	I27122 = NAND(WX8341, I27121)
--	I27123 = NAND(WX8249, I27121)
--	WX8785 = NAND(I27122, I27123)
--	I27134 = NAND(WX8342, WX8251)
--	I27135 = NAND(WX8342, I27134)
--	I27136 = NAND(WX8251, I27134)
--	WX8792 = NAND(I27135, I27136)
--	I27147 = NAND(WX8343, WX8253)
--	I27148 = NAND(WX8343, I27147)
--	I27149 = NAND(WX8253, I27147)
--	WX8799 = NAND(I27148, I27149)
--	I27160 = NAND(WX8344, WX8255)
--	I27161 = NAND(WX8344, I27160)
--	I27162 = NAND(WX8255, I27160)
--	WX8806 = NAND(I27161, I27162)
--	I27173 = NAND(WX8345, WX8257)
--	I27174 = NAND(WX8345, I27173)
--	I27175 = NAND(WX8257, I27173)
--	WX8813 = NAND(I27174, I27175)
--	I27186 = NAND(WX8346, WX8259)
--	I27187 = NAND(WX8346, I27186)
--	I27188 = NAND(WX8259, I27186)
--	WX8820 = NAND(I27187, I27188)
--	I27199 = NAND(WX8347, WX8261)
--	I27200 = NAND(WX8347, I27199)
--	I27201 = NAND(WX8261, I27199)
--	WX8827 = NAND(I27200, I27201)
--	I27212 = NAND(WX8348, WX8263)
--	I27213 = NAND(WX8348, I27212)
--	I27214 = NAND(WX8263, I27212)
--	WX8834 = NAND(I27213, I27214)
--	I27225 = NAND(WX8349, WX8265)
--	I27226 = NAND(WX8349, I27225)
--	I27227 = NAND(WX8265, I27225)
--	WX8841 = NAND(I27226, I27227)
--	I27238 = NAND(WX8350, WX8267)
--	I27239 = NAND(WX8350, I27238)
--	I27240 = NAND(WX8267, I27238)
--	WX8848 = NAND(I27239, I27240)
--	I27251 = NAND(WX8351, WX8269)
--	I27252 = NAND(WX8351, I27251)
--	I27253 = NAND(WX8269, I27251)
--	WX8855 = NAND(I27252, I27253)
--	I27264 = NAND(WX8352, WX8271)
--	I27265 = NAND(WX8352, I27264)
--	I27266 = NAND(WX8271, I27264)
--	WX8862 = NAND(I27265, I27266)
--	I27277 = NAND(WX8353, WX8273)
--	I27278 = NAND(WX8353, I27277)
--	I27279 = NAND(WX8273, I27277)
--	WX8869 = NAND(I27278, I27279)
--	I27290 = NAND(WX8354, WX8275)
--	I27291 = NAND(WX8354, I27290)
--	I27292 = NAND(WX8275, I27290)
--	WX8876 = NAND(I27291, I27292)
--	I27303 = NAND(WX8355, WX8277)
--	I27304 = NAND(WX8355, I27303)
--	I27305 = NAND(WX8277, I27303)
--	WX8883 = NAND(I27304, I27305)
--	I27316 = NAND(WX8356, WX8279)
--	I27317 = NAND(WX8356, I27316)
--	I27318 = NAND(WX8279, I27316)
--	WX8890 = NAND(I27317, I27318)
--	I27329 = NAND(WX8357, WX8281)
--	I27330 = NAND(WX8357, I27329)
--	I27331 = NAND(WX8281, I27329)
--	WX8897 = NAND(I27330, I27331)
--	I27342 = NAND(WX8358, WX8283)
--	I27343 = NAND(WX8358, I27342)
--	I27344 = NAND(WX8283, I27342)
--	WX8904 = NAND(I27343, I27344)
--	I27355 = NAND(WX8359, WX8285)
--	I27356 = NAND(WX8359, I27355)
--	I27357 = NAND(WX8285, I27355)
--	WX8911 = NAND(I27356, I27357)
--	I27368 = NAND(WX8360, WX8287)
--	I27369 = NAND(WX8360, I27368)
--	I27370 = NAND(WX8287, I27368)
--	WX8918 = NAND(I27369, I27370)
--	I27381 = NAND(WX8361, WX8289)
--	I27382 = NAND(WX8361, I27381)
--	I27383 = NAND(WX8289, I27381)
--	WX8925 = NAND(I27382, I27383)
--	I27394 = NAND(WX8362, WX8291)
--	I27395 = NAND(WX8362, I27394)
--	I27396 = NAND(WX8291, I27394)
--	WX8932 = NAND(I27395, I27396)
--	I27407 = NAND(WX8363, WX8293)
--	I27408 = NAND(WX8363, I27407)
--	I27409 = NAND(WX8293, I27407)
--	WX8939 = NAND(I27408, I27409)
--	I27420 = NAND(WX8364, WX8295)
--	I27421 = NAND(WX8364, I27420)
--	I27422 = NAND(WX8295, I27420)
--	WX8946 = NAND(I27421, I27422)
--	I27433 = NAND(WX8365, WX8297)
--	I27434 = NAND(WX8365, I27433)
--	I27435 = NAND(WX8297, I27433)
--	WX8953 = NAND(I27434, I27435)
--	I27446 = NAND(WX8366, WX8299)
--	I27447 = NAND(WX8366, I27446)
--	I27448 = NAND(WX8299, I27446)
--	WX8960 = NAND(I27447, I27448)
--	I27459 = NAND(WX8367, WX8301)
--	I27460 = NAND(WX8367, I27459)
--	I27461 = NAND(WX8301, I27459)
--	WX8967 = NAND(I27460, I27461)
--	I27472 = NAND(WX8368, WX8303)
--	I27473 = NAND(WX8368, I27472)
--	I27474 = NAND(WX8303, I27472)
--	WX8974 = NAND(I27473, I27474)
--	I27485 = NAND(WX8369, WX8305)
--	I27486 = NAND(WX8369, I27485)
--	I27487 = NAND(WX8305, I27485)
--	WX8981 = NAND(I27486, I27487)
--	I27500 = NAND(WX8385, CRC_OUT_3_31)
--	I27501 = NAND(WX8385, I27500)
--	I27502 = NAND(CRC_OUT_3_31, I27500)
--	I27499 = NAND(I27501, I27502)
--	I27507 = NAND(CRC_OUT_3_15, I27499)
--	I27508 = NAND(CRC_OUT_3_15, I27507)
--	I27509 = NAND(I27499, I27507)
--	WX8989 = NAND(I27508, I27509)
--	I27515 = NAND(WX8390, CRC_OUT_3_31)
--	I27516 = NAND(WX8390, I27515)
--	I27517 = NAND(CRC_OUT_3_31, I27515)
--	I27514 = NAND(I27516, I27517)
--	I27522 = NAND(CRC_OUT_3_10, I27514)
--	I27523 = NAND(CRC_OUT_3_10, I27522)
--	I27524 = NAND(I27514, I27522)
--	WX8990 = NAND(I27523, I27524)
--	I27530 = NAND(WX8397, CRC_OUT_3_31)
--	I27531 = NAND(WX8397, I27530)
--	I27532 = NAND(CRC_OUT_3_31, I27530)
--	I27529 = NAND(I27531, I27532)
--	I27537 = NAND(CRC_OUT_3_3, I27529)
--	I27538 = NAND(CRC_OUT_3_3, I27537)
--	I27539 = NAND(I27529, I27537)
--	WX8991 = NAND(I27538, I27539)
--	I27544 = NAND(WX8401, CRC_OUT_3_31)
--	I27545 = NAND(WX8401, I27544)
--	I27546 = NAND(CRC_OUT_3_31, I27544)
--	WX8992 = NAND(I27545, I27546)
--	I27551 = NAND(WX8370, CRC_OUT_3_30)
--	I27552 = NAND(WX8370, I27551)
--	I27553 = NAND(CRC_OUT_3_30, I27551)
--	WX8993 = NAND(I27552, I27553)
--	I27558 = NAND(WX8371, CRC_OUT_3_29)
--	I27559 = NAND(WX8371, I27558)
--	I27560 = NAND(CRC_OUT_3_29, I27558)
--	WX8994 = NAND(I27559, I27560)
--	I27565 = NAND(WX8372, CRC_OUT_3_28)
--	I27566 = NAND(WX8372, I27565)
--	I27567 = NAND(CRC_OUT_3_28, I27565)
--	WX8995 = NAND(I27566, I27567)
--	I27572 = NAND(WX8373, CRC_OUT_3_27)
--	I27573 = NAND(WX8373, I27572)
--	I27574 = NAND(CRC_OUT_3_27, I27572)
--	WX8996 = NAND(I27573, I27574)
--	I27579 = NAND(WX8374, CRC_OUT_3_26)
--	I27580 = NAND(WX8374, I27579)
--	I27581 = NAND(CRC_OUT_3_26, I27579)
--	WX8997 = NAND(I27580, I27581)
--	I27586 = NAND(WX8375, CRC_OUT_3_25)
--	I27587 = NAND(WX8375, I27586)
--	I27588 = NAND(CRC_OUT_3_25, I27586)
--	WX8998 = NAND(I27587, I27588)
--	I27593 = NAND(WX8376, CRC_OUT_3_24)
--	I27594 = NAND(WX8376, I27593)
--	I27595 = NAND(CRC_OUT_3_24, I27593)
--	WX8999 = NAND(I27594, I27595)
--	I27600 = NAND(WX8377, CRC_OUT_3_23)
--	I27601 = NAND(WX8377, I27600)
--	I27602 = NAND(CRC_OUT_3_23, I27600)
--	WX9000 = NAND(I27601, I27602)
--	I27607 = NAND(WX8378, CRC_OUT_3_22)
--	I27608 = NAND(WX8378, I27607)
--	I27609 = NAND(CRC_OUT_3_22, I27607)
--	WX9001 = NAND(I27608, I27609)
--	I27614 = NAND(WX8379, CRC_OUT_3_21)
--	I27615 = NAND(WX8379, I27614)
--	I27616 = NAND(CRC_OUT_3_21, I27614)
--	WX9002 = NAND(I27615, I27616)
--	I27621 = NAND(WX8380, CRC_OUT_3_20)
--	I27622 = NAND(WX8380, I27621)
--	I27623 = NAND(CRC_OUT_3_20, I27621)
--	WX9003 = NAND(I27622, I27623)
--	I27628 = NAND(WX8381, CRC_OUT_3_19)
--	I27629 = NAND(WX8381, I27628)
--	I27630 = NAND(CRC_OUT_3_19, I27628)
--	WX9004 = NAND(I27629, I27630)
--	I27635 = NAND(WX8382, CRC_OUT_3_18)
--	I27636 = NAND(WX8382, I27635)
--	I27637 = NAND(CRC_OUT_3_18, I27635)
--	WX9005 = NAND(I27636, I27637)
--	I27642 = NAND(WX8383, CRC_OUT_3_17)
--	I27643 = NAND(WX8383, I27642)
--	I27644 = NAND(CRC_OUT_3_17, I27642)
--	WX9006 = NAND(I27643, I27644)
--	I27649 = NAND(WX8384, CRC_OUT_3_16)
--	I27650 = NAND(WX8384, I27649)
--	I27651 = NAND(CRC_OUT_3_16, I27649)
--	WX9007 = NAND(I27650, I27651)
--	I27656 = NAND(WX8386, CRC_OUT_3_14)
--	I27657 = NAND(WX8386, I27656)
--	I27658 = NAND(CRC_OUT_3_14, I27656)
--	WX9008 = NAND(I27657, I27658)
--	I27663 = NAND(WX8387, CRC_OUT_3_13)
--	I27664 = NAND(WX8387, I27663)
--	I27665 = NAND(CRC_OUT_3_13, I27663)
--	WX9009 = NAND(I27664, I27665)
--	I27670 = NAND(WX8388, CRC_OUT_3_12)
--	I27671 = NAND(WX8388, I27670)
--	I27672 = NAND(CRC_OUT_3_12, I27670)
--	WX9010 = NAND(I27671, I27672)
--	I27677 = NAND(WX8389, CRC_OUT_3_11)
--	I27678 = NAND(WX8389, I27677)
--	I27679 = NAND(CRC_OUT_3_11, I27677)
--	WX9011 = NAND(I27678, I27679)
--	I27684 = NAND(WX8391, CRC_OUT_3_9)
--	I27685 = NAND(WX8391, I27684)
--	I27686 = NAND(CRC_OUT_3_9, I27684)
--	WX9012 = NAND(I27685, I27686)
--	I27691 = NAND(WX8392, CRC_OUT_3_8)
--	I27692 = NAND(WX8392, I27691)
--	I27693 = NAND(CRC_OUT_3_8, I27691)
--	WX9013 = NAND(I27692, I27693)
--	I27698 = NAND(WX8393, CRC_OUT_3_7)
--	I27699 = NAND(WX8393, I27698)
--	I27700 = NAND(CRC_OUT_3_7, I27698)
--	WX9014 = NAND(I27699, I27700)
--	I27705 = NAND(WX8394, CRC_OUT_3_6)
--	I27706 = NAND(WX8394, I27705)
--	I27707 = NAND(CRC_OUT_3_6, I27705)
--	WX9015 = NAND(I27706, I27707)
--	I27712 = NAND(WX8395, CRC_OUT_3_5)
--	I27713 = NAND(WX8395, I27712)
--	I27714 = NAND(CRC_OUT_3_5, I27712)
--	WX9016 = NAND(I27713, I27714)
--	I27719 = NAND(WX8396, CRC_OUT_3_4)
--	I27720 = NAND(WX8396, I27719)
--	I27721 = NAND(CRC_OUT_3_4, I27719)
--	WX9017 = NAND(I27720, I27721)
--	I27726 = NAND(WX8398, CRC_OUT_3_2)
--	I27727 = NAND(WX8398, I27726)
--	I27728 = NAND(CRC_OUT_3_2, I27726)
--	WX9018 = NAND(I27727, I27728)
--	I27733 = NAND(WX8399, CRC_OUT_3_1)
--	I27734 = NAND(WX8399, I27733)
--	I27735 = NAND(CRC_OUT_3_1, I27733)
--	WX9019 = NAND(I27734, I27735)
--	I27740 = NAND(WX8400, CRC_OUT_3_0)
--	I27741 = NAND(WX8400, I27740)
--	I27742 = NAND(CRC_OUT_3_0, I27740)
--	WX9020 = NAND(I27741, I27742)
--	I30023 = NAND(WX10052, WX9696)
--	I30024 = NAND(WX10052, I30023)
--	I30025 = NAND(WX9696, I30023)
--	I30022 = NAND(I30024, I30025)
--	I30030 = NAND(WX9760, I30022)
--	I30031 = NAND(WX9760, I30030)
--	I30032 = NAND(I30022, I30030)
--	I30021 = NAND(I30031, I30032)
--	I30038 = NAND(WX9824, WX9888)
--	I30039 = NAND(WX9824, I30038)
--	I30040 = NAND(WX9888, I30038)
--	I30037 = NAND(I30039, I30040)
--	I30045 = NAND(I30021, I30037)
--	I30046 = NAND(I30021, I30045)
--	I30047 = NAND(I30037, I30045)
--	WX9951 = NAND(I30046, I30047)
--	I30054 = NAND(WX10052, WX9698)
--	I30055 = NAND(WX10052, I30054)
--	I30056 = NAND(WX9698, I30054)
--	I30053 = NAND(I30055, I30056)
--	I30061 = NAND(WX9762, I30053)
--	I30062 = NAND(WX9762, I30061)
--	I30063 = NAND(I30053, I30061)
--	I30052 = NAND(I30062, I30063)
--	I30069 = NAND(WX9826, WX9890)
--	I30070 = NAND(WX9826, I30069)
--	I30071 = NAND(WX9890, I30069)
--	I30068 = NAND(I30070, I30071)
--	I30076 = NAND(I30052, I30068)
--	I30077 = NAND(I30052, I30076)
--	I30078 = NAND(I30068, I30076)
--	WX9952 = NAND(I30077, I30078)
--	I30085 = NAND(WX10052, WX9700)
--	I30086 = NAND(WX10052, I30085)
--	I30087 = NAND(WX9700, I30085)
--	I30084 = NAND(I30086, I30087)
--	I30092 = NAND(WX9764, I30084)
--	I30093 = NAND(WX9764, I30092)
--	I30094 = NAND(I30084, I30092)
--	I30083 = NAND(I30093, I30094)
--	I30100 = NAND(WX9828, WX9892)
--	I30101 = NAND(WX9828, I30100)
--	I30102 = NAND(WX9892, I30100)
--	I30099 = NAND(I30101, I30102)
--	I30107 = NAND(I30083, I30099)
--	I30108 = NAND(I30083, I30107)
--	I30109 = NAND(I30099, I30107)
--	WX9953 = NAND(I30108, I30109)
--	I30116 = NAND(WX10052, WX9702)
--	I30117 = NAND(WX10052, I30116)
--	I30118 = NAND(WX9702, I30116)
--	I30115 = NAND(I30117, I30118)
--	I30123 = NAND(WX9766, I30115)
--	I30124 = NAND(WX9766, I30123)
--	I30125 = NAND(I30115, I30123)
--	I30114 = NAND(I30124, I30125)
--	I30131 = NAND(WX9830, WX9894)
--	I30132 = NAND(WX9830, I30131)
--	I30133 = NAND(WX9894, I30131)
--	I30130 = NAND(I30132, I30133)
--	I30138 = NAND(I30114, I30130)
--	I30139 = NAND(I30114, I30138)
--	I30140 = NAND(I30130, I30138)
--	WX9954 = NAND(I30139, I30140)
--	I30147 = NAND(WX10052, WX9704)
--	I30148 = NAND(WX10052, I30147)
--	I30149 = NAND(WX9704, I30147)
--	I30146 = NAND(I30148, I30149)
--	I30154 = NAND(WX9768, I30146)
--	I30155 = NAND(WX9768, I30154)
--	I30156 = NAND(I30146, I30154)
--	I30145 = NAND(I30155, I30156)
--	I30162 = NAND(WX9832, WX9896)
--	I30163 = NAND(WX9832, I30162)
--	I30164 = NAND(WX9896, I30162)
--	I30161 = NAND(I30163, I30164)
--	I30169 = NAND(I30145, I30161)
--	I30170 = NAND(I30145, I30169)
--	I30171 = NAND(I30161, I30169)
--	WX9955 = NAND(I30170, I30171)
--	I30178 = NAND(WX10052, WX9706)
--	I30179 = NAND(WX10052, I30178)
--	I30180 = NAND(WX9706, I30178)
--	I30177 = NAND(I30179, I30180)
--	I30185 = NAND(WX9770, I30177)
--	I30186 = NAND(WX9770, I30185)
--	I30187 = NAND(I30177, I30185)
--	I30176 = NAND(I30186, I30187)
--	I30193 = NAND(WX9834, WX9898)
--	I30194 = NAND(WX9834, I30193)
--	I30195 = NAND(WX9898, I30193)
--	I30192 = NAND(I30194, I30195)
--	I30200 = NAND(I30176, I30192)
--	I30201 = NAND(I30176, I30200)
--	I30202 = NAND(I30192, I30200)
--	WX9956 = NAND(I30201, I30202)
--	I30209 = NAND(WX10052, WX9708)
--	I30210 = NAND(WX10052, I30209)
--	I30211 = NAND(WX9708, I30209)
--	I30208 = NAND(I30210, I30211)
--	I30216 = NAND(WX9772, I30208)
--	I30217 = NAND(WX9772, I30216)
--	I30218 = NAND(I30208, I30216)
--	I30207 = NAND(I30217, I30218)
--	I30224 = NAND(WX9836, WX9900)
--	I30225 = NAND(WX9836, I30224)
--	I30226 = NAND(WX9900, I30224)
--	I30223 = NAND(I30225, I30226)
--	I30231 = NAND(I30207, I30223)
--	I30232 = NAND(I30207, I30231)
--	I30233 = NAND(I30223, I30231)
--	WX9957 = NAND(I30232, I30233)
--	I30240 = NAND(WX10052, WX9710)
--	I30241 = NAND(WX10052, I30240)
--	I30242 = NAND(WX9710, I30240)
--	I30239 = NAND(I30241, I30242)
--	I30247 = NAND(WX9774, I30239)
--	I30248 = NAND(WX9774, I30247)
--	I30249 = NAND(I30239, I30247)
--	I30238 = NAND(I30248, I30249)
--	I30255 = NAND(WX9838, WX9902)
--	I30256 = NAND(WX9838, I30255)
--	I30257 = NAND(WX9902, I30255)
--	I30254 = NAND(I30256, I30257)
--	I30262 = NAND(I30238, I30254)
--	I30263 = NAND(I30238, I30262)
--	I30264 = NAND(I30254, I30262)
--	WX9958 = NAND(I30263, I30264)
--	I30271 = NAND(WX10052, WX9712)
--	I30272 = NAND(WX10052, I30271)
--	I30273 = NAND(WX9712, I30271)
--	I30270 = NAND(I30272, I30273)
--	I30278 = NAND(WX9776, I30270)
--	I30279 = NAND(WX9776, I30278)
--	I30280 = NAND(I30270, I30278)
--	I30269 = NAND(I30279, I30280)
--	I30286 = NAND(WX9840, WX9904)
--	I30287 = NAND(WX9840, I30286)
--	I30288 = NAND(WX9904, I30286)
--	I30285 = NAND(I30287, I30288)
--	I30293 = NAND(I30269, I30285)
--	I30294 = NAND(I30269, I30293)
--	I30295 = NAND(I30285, I30293)
--	WX9959 = NAND(I30294, I30295)
--	I30302 = NAND(WX10052, WX9714)
--	I30303 = NAND(WX10052, I30302)
--	I30304 = NAND(WX9714, I30302)
--	I30301 = NAND(I30303, I30304)
--	I30309 = NAND(WX9778, I30301)
--	I30310 = NAND(WX9778, I30309)
--	I30311 = NAND(I30301, I30309)
--	I30300 = NAND(I30310, I30311)
--	I30317 = NAND(WX9842, WX9906)
--	I30318 = NAND(WX9842, I30317)
--	I30319 = NAND(WX9906, I30317)
--	I30316 = NAND(I30318, I30319)
--	I30324 = NAND(I30300, I30316)
--	I30325 = NAND(I30300, I30324)
--	I30326 = NAND(I30316, I30324)
--	WX9960 = NAND(I30325, I30326)
--	I30333 = NAND(WX10052, WX9716)
--	I30334 = NAND(WX10052, I30333)
--	I30335 = NAND(WX9716, I30333)
--	I30332 = NAND(I30334, I30335)
--	I30340 = NAND(WX9780, I30332)
--	I30341 = NAND(WX9780, I30340)
--	I30342 = NAND(I30332, I30340)
--	I30331 = NAND(I30341, I30342)
--	I30348 = NAND(WX9844, WX9908)
--	I30349 = NAND(WX9844, I30348)
--	I30350 = NAND(WX9908, I30348)
--	I30347 = NAND(I30349, I30350)
--	I30355 = NAND(I30331, I30347)
--	I30356 = NAND(I30331, I30355)
--	I30357 = NAND(I30347, I30355)
--	WX9961 = NAND(I30356, I30357)
--	I30364 = NAND(WX10052, WX9718)
--	I30365 = NAND(WX10052, I30364)
--	I30366 = NAND(WX9718, I30364)
--	I30363 = NAND(I30365, I30366)
--	I30371 = NAND(WX9782, I30363)
--	I30372 = NAND(WX9782, I30371)
--	I30373 = NAND(I30363, I30371)
--	I30362 = NAND(I30372, I30373)
--	I30379 = NAND(WX9846, WX9910)
--	I30380 = NAND(WX9846, I30379)
--	I30381 = NAND(WX9910, I30379)
--	I30378 = NAND(I30380, I30381)
--	I30386 = NAND(I30362, I30378)
--	I30387 = NAND(I30362, I30386)
--	I30388 = NAND(I30378, I30386)
--	WX9962 = NAND(I30387, I30388)
--	I30395 = NAND(WX10052, WX9720)
--	I30396 = NAND(WX10052, I30395)
--	I30397 = NAND(WX9720, I30395)
--	I30394 = NAND(I30396, I30397)
--	I30402 = NAND(WX9784, I30394)
--	I30403 = NAND(WX9784, I30402)
--	I30404 = NAND(I30394, I30402)
--	I30393 = NAND(I30403, I30404)
--	I30410 = NAND(WX9848, WX9912)
--	I30411 = NAND(WX9848, I30410)
--	I30412 = NAND(WX9912, I30410)
--	I30409 = NAND(I30411, I30412)
--	I30417 = NAND(I30393, I30409)
--	I30418 = NAND(I30393, I30417)
--	I30419 = NAND(I30409, I30417)
--	WX9963 = NAND(I30418, I30419)
--	I30426 = NAND(WX10052, WX9722)
--	I30427 = NAND(WX10052, I30426)
--	I30428 = NAND(WX9722, I30426)
--	I30425 = NAND(I30427, I30428)
--	I30433 = NAND(WX9786, I30425)
--	I30434 = NAND(WX9786, I30433)
--	I30435 = NAND(I30425, I30433)
--	I30424 = NAND(I30434, I30435)
--	I30441 = NAND(WX9850, WX9914)
--	I30442 = NAND(WX9850, I30441)
--	I30443 = NAND(WX9914, I30441)
--	I30440 = NAND(I30442, I30443)
--	I30448 = NAND(I30424, I30440)
--	I30449 = NAND(I30424, I30448)
--	I30450 = NAND(I30440, I30448)
--	WX9964 = NAND(I30449, I30450)
--	I30457 = NAND(WX10052, WX9724)
--	I30458 = NAND(WX10052, I30457)
--	I30459 = NAND(WX9724, I30457)
--	I30456 = NAND(I30458, I30459)
--	I30464 = NAND(WX9788, I30456)
--	I30465 = NAND(WX9788, I30464)
--	I30466 = NAND(I30456, I30464)
--	I30455 = NAND(I30465, I30466)
--	I30472 = NAND(WX9852, WX9916)
--	I30473 = NAND(WX9852, I30472)
--	I30474 = NAND(WX9916, I30472)
--	I30471 = NAND(I30473, I30474)
--	I30479 = NAND(I30455, I30471)
--	I30480 = NAND(I30455, I30479)
--	I30481 = NAND(I30471, I30479)
--	WX9965 = NAND(I30480, I30481)
--	I30488 = NAND(WX10052, WX9726)
--	I30489 = NAND(WX10052, I30488)
--	I30490 = NAND(WX9726, I30488)
--	I30487 = NAND(I30489, I30490)
--	I30495 = NAND(WX9790, I30487)
--	I30496 = NAND(WX9790, I30495)
--	I30497 = NAND(I30487, I30495)
--	I30486 = NAND(I30496, I30497)
--	I30503 = NAND(WX9854, WX9918)
--	I30504 = NAND(WX9854, I30503)
--	I30505 = NAND(WX9918, I30503)
--	I30502 = NAND(I30504, I30505)
--	I30510 = NAND(I30486, I30502)
--	I30511 = NAND(I30486, I30510)
--	I30512 = NAND(I30502, I30510)
--	WX9966 = NAND(I30511, I30512)
--	I30519 = NAND(WX10053, WX9728)
--	I30520 = NAND(WX10053, I30519)
--	I30521 = NAND(WX9728, I30519)
--	I30518 = NAND(I30520, I30521)
--	I30526 = NAND(WX9792, I30518)
--	I30527 = NAND(WX9792, I30526)
--	I30528 = NAND(I30518, I30526)
--	I30517 = NAND(I30527, I30528)
--	I30534 = NAND(WX9856, WX9920)
--	I30535 = NAND(WX9856, I30534)
--	I30536 = NAND(WX9920, I30534)
--	I30533 = NAND(I30535, I30536)
--	I30541 = NAND(I30517, I30533)
--	I30542 = NAND(I30517, I30541)
--	I30543 = NAND(I30533, I30541)
--	WX9967 = NAND(I30542, I30543)
--	I30550 = NAND(WX10053, WX9730)
--	I30551 = NAND(WX10053, I30550)
--	I30552 = NAND(WX9730, I30550)
--	I30549 = NAND(I30551, I30552)
--	I30557 = NAND(WX9794, I30549)
--	I30558 = NAND(WX9794, I30557)
--	I30559 = NAND(I30549, I30557)
--	I30548 = NAND(I30558, I30559)
--	I30565 = NAND(WX9858, WX9922)
--	I30566 = NAND(WX9858, I30565)
--	I30567 = NAND(WX9922, I30565)
--	I30564 = NAND(I30566, I30567)
--	I30572 = NAND(I30548, I30564)
--	I30573 = NAND(I30548, I30572)
--	I30574 = NAND(I30564, I30572)
--	WX9968 = NAND(I30573, I30574)
--	I30581 = NAND(WX10053, WX9732)
--	I30582 = NAND(WX10053, I30581)
--	I30583 = NAND(WX9732, I30581)
--	I30580 = NAND(I30582, I30583)
--	I30588 = NAND(WX9796, I30580)
--	I30589 = NAND(WX9796, I30588)
--	I30590 = NAND(I30580, I30588)
--	I30579 = NAND(I30589, I30590)
--	I30596 = NAND(WX9860, WX9924)
--	I30597 = NAND(WX9860, I30596)
--	I30598 = NAND(WX9924, I30596)
--	I30595 = NAND(I30597, I30598)
--	I30603 = NAND(I30579, I30595)
--	I30604 = NAND(I30579, I30603)
--	I30605 = NAND(I30595, I30603)
--	WX9969 = NAND(I30604, I30605)
--	I30612 = NAND(WX10053, WX9734)
--	I30613 = NAND(WX10053, I30612)
--	I30614 = NAND(WX9734, I30612)
--	I30611 = NAND(I30613, I30614)
--	I30619 = NAND(WX9798, I30611)
--	I30620 = NAND(WX9798, I30619)
--	I30621 = NAND(I30611, I30619)
--	I30610 = NAND(I30620, I30621)
--	I30627 = NAND(WX9862, WX9926)
--	I30628 = NAND(WX9862, I30627)
--	I30629 = NAND(WX9926, I30627)
--	I30626 = NAND(I30628, I30629)
--	I30634 = NAND(I30610, I30626)
--	I30635 = NAND(I30610, I30634)
--	I30636 = NAND(I30626, I30634)
--	WX9970 = NAND(I30635, I30636)
--	I30643 = NAND(WX10053, WX9736)
--	I30644 = NAND(WX10053, I30643)
--	I30645 = NAND(WX9736, I30643)
--	I30642 = NAND(I30644, I30645)
--	I30650 = NAND(WX9800, I30642)
--	I30651 = NAND(WX9800, I30650)
--	I30652 = NAND(I30642, I30650)
--	I30641 = NAND(I30651, I30652)
--	I30658 = NAND(WX9864, WX9928)
--	I30659 = NAND(WX9864, I30658)
--	I30660 = NAND(WX9928, I30658)
--	I30657 = NAND(I30659, I30660)
--	I30665 = NAND(I30641, I30657)
--	I30666 = NAND(I30641, I30665)
--	I30667 = NAND(I30657, I30665)
--	WX9971 = NAND(I30666, I30667)
--	I30674 = NAND(WX10053, WX9738)
--	I30675 = NAND(WX10053, I30674)
--	I30676 = NAND(WX9738, I30674)
--	I30673 = NAND(I30675, I30676)
--	I30681 = NAND(WX9802, I30673)
--	I30682 = NAND(WX9802, I30681)
--	I30683 = NAND(I30673, I30681)
--	I30672 = NAND(I30682, I30683)
--	I30689 = NAND(WX9866, WX9930)
--	I30690 = NAND(WX9866, I30689)
--	I30691 = NAND(WX9930, I30689)
--	I30688 = NAND(I30690, I30691)
--	I30696 = NAND(I30672, I30688)
--	I30697 = NAND(I30672, I30696)
--	I30698 = NAND(I30688, I30696)
--	WX9972 = NAND(I30697, I30698)
--	I30705 = NAND(WX10053, WX9740)
--	I30706 = NAND(WX10053, I30705)
--	I30707 = NAND(WX9740, I30705)
--	I30704 = NAND(I30706, I30707)
--	I30712 = NAND(WX9804, I30704)
--	I30713 = NAND(WX9804, I30712)
--	I30714 = NAND(I30704, I30712)
--	I30703 = NAND(I30713, I30714)
--	I30720 = NAND(WX9868, WX9932)
--	I30721 = NAND(WX9868, I30720)
--	I30722 = NAND(WX9932, I30720)
--	I30719 = NAND(I30721, I30722)
--	I30727 = NAND(I30703, I30719)
--	I30728 = NAND(I30703, I30727)
--	I30729 = NAND(I30719, I30727)
--	WX9973 = NAND(I30728, I30729)
--	I30736 = NAND(WX10053, WX9742)
--	I30737 = NAND(WX10053, I30736)
--	I30738 = NAND(WX9742, I30736)
--	I30735 = NAND(I30737, I30738)
--	I30743 = NAND(WX9806, I30735)
--	I30744 = NAND(WX9806, I30743)
--	I30745 = NAND(I30735, I30743)
--	I30734 = NAND(I30744, I30745)
--	I30751 = NAND(WX9870, WX9934)
--	I30752 = NAND(WX9870, I30751)
--	I30753 = NAND(WX9934, I30751)
--	I30750 = NAND(I30752, I30753)
--	I30758 = NAND(I30734, I30750)
--	I30759 = NAND(I30734, I30758)
--	I30760 = NAND(I30750, I30758)
--	WX9974 = NAND(I30759, I30760)
--	I30767 = NAND(WX10053, WX9744)
--	I30768 = NAND(WX10053, I30767)
--	I30769 = NAND(WX9744, I30767)
--	I30766 = NAND(I30768, I30769)
--	I30774 = NAND(WX9808, I30766)
--	I30775 = NAND(WX9808, I30774)
--	I30776 = NAND(I30766, I30774)
--	I30765 = NAND(I30775, I30776)
--	I30782 = NAND(WX9872, WX9936)
--	I30783 = NAND(WX9872, I30782)
--	I30784 = NAND(WX9936, I30782)
--	I30781 = NAND(I30783, I30784)
--	I30789 = NAND(I30765, I30781)
--	I30790 = NAND(I30765, I30789)
--	I30791 = NAND(I30781, I30789)
--	WX9975 = NAND(I30790, I30791)
--	I30798 = NAND(WX10053, WX9746)
--	I30799 = NAND(WX10053, I30798)
--	I30800 = NAND(WX9746, I30798)
--	I30797 = NAND(I30799, I30800)
--	I30805 = NAND(WX9810, I30797)
--	I30806 = NAND(WX9810, I30805)
--	I30807 = NAND(I30797, I30805)
--	I30796 = NAND(I30806, I30807)
--	I30813 = NAND(WX9874, WX9938)
--	I30814 = NAND(WX9874, I30813)
--	I30815 = NAND(WX9938, I30813)
--	I30812 = NAND(I30814, I30815)
--	I30820 = NAND(I30796, I30812)
--	I30821 = NAND(I30796, I30820)
--	I30822 = NAND(I30812, I30820)
--	WX9976 = NAND(I30821, I30822)
--	I30829 = NAND(WX10053, WX9748)
--	I30830 = NAND(WX10053, I30829)
--	I30831 = NAND(WX9748, I30829)
--	I30828 = NAND(I30830, I30831)
--	I30836 = NAND(WX9812, I30828)
--	I30837 = NAND(WX9812, I30836)
--	I30838 = NAND(I30828, I30836)
--	I30827 = NAND(I30837, I30838)
--	I30844 = NAND(WX9876, WX9940)
--	I30845 = NAND(WX9876, I30844)
--	I30846 = NAND(WX9940, I30844)
--	I30843 = NAND(I30845, I30846)
--	I30851 = NAND(I30827, I30843)
--	I30852 = NAND(I30827, I30851)
--	I30853 = NAND(I30843, I30851)
--	WX9977 = NAND(I30852, I30853)
--	I30860 = NAND(WX10053, WX9750)
--	I30861 = NAND(WX10053, I30860)
--	I30862 = NAND(WX9750, I30860)
--	I30859 = NAND(I30861, I30862)
--	I30867 = NAND(WX9814, I30859)
--	I30868 = NAND(WX9814, I30867)
--	I30869 = NAND(I30859, I30867)
--	I30858 = NAND(I30868, I30869)
--	I30875 = NAND(WX9878, WX9942)
--	I30876 = NAND(WX9878, I30875)
--	I30877 = NAND(WX9942, I30875)
--	I30874 = NAND(I30876, I30877)
--	I30882 = NAND(I30858, I30874)
--	I30883 = NAND(I30858, I30882)
--	I30884 = NAND(I30874, I30882)
--	WX9978 = NAND(I30883, I30884)
--	I30891 = NAND(WX10053, WX9752)
--	I30892 = NAND(WX10053, I30891)
--	I30893 = NAND(WX9752, I30891)
--	I30890 = NAND(I30892, I30893)
--	I30898 = NAND(WX9816, I30890)
--	I30899 = NAND(WX9816, I30898)
--	I30900 = NAND(I30890, I30898)
--	I30889 = NAND(I30899, I30900)
--	I30906 = NAND(WX9880, WX9944)
--	I30907 = NAND(WX9880, I30906)
--	I30908 = NAND(WX9944, I30906)
--	I30905 = NAND(I30907, I30908)
--	I30913 = NAND(I30889, I30905)
--	I30914 = NAND(I30889, I30913)
--	I30915 = NAND(I30905, I30913)
--	WX9979 = NAND(I30914, I30915)
--	I30922 = NAND(WX10053, WX9754)
--	I30923 = NAND(WX10053, I30922)
--	I30924 = NAND(WX9754, I30922)
--	I30921 = NAND(I30923, I30924)
--	I30929 = NAND(WX9818, I30921)
--	I30930 = NAND(WX9818, I30929)
--	I30931 = NAND(I30921, I30929)
--	I30920 = NAND(I30930, I30931)
--	I30937 = NAND(WX9882, WX9946)
--	I30938 = NAND(WX9882, I30937)
--	I30939 = NAND(WX9946, I30937)
--	I30936 = NAND(I30938, I30939)
--	I30944 = NAND(I30920, I30936)
--	I30945 = NAND(I30920, I30944)
--	I30946 = NAND(I30936, I30944)
--	WX9980 = NAND(I30945, I30946)
--	I30953 = NAND(WX10053, WX9756)
--	I30954 = NAND(WX10053, I30953)
--	I30955 = NAND(WX9756, I30953)
--	I30952 = NAND(I30954, I30955)
--	I30960 = NAND(WX9820, I30952)
--	I30961 = NAND(WX9820, I30960)
--	I30962 = NAND(I30952, I30960)
--	I30951 = NAND(I30961, I30962)
--	I30968 = NAND(WX9884, WX9948)
--	I30969 = NAND(WX9884, I30968)
--	I30970 = NAND(WX9948, I30968)
--	I30967 = NAND(I30969, I30970)
--	I30975 = NAND(I30951, I30967)
--	I30976 = NAND(I30951, I30975)
--	I30977 = NAND(I30967, I30975)
--	WX9981 = NAND(I30976, I30977)
--	I30984 = NAND(WX10053, WX9758)
--	I30985 = NAND(WX10053, I30984)
--	I30986 = NAND(WX9758, I30984)
--	I30983 = NAND(I30985, I30986)
--	I30991 = NAND(WX9822, I30983)
--	I30992 = NAND(WX9822, I30991)
--	I30993 = NAND(I30983, I30991)
--	I30982 = NAND(I30992, I30993)
--	I30999 = NAND(WX9886, WX9950)
--	I31000 = NAND(WX9886, I30999)
--	I31001 = NAND(WX9950, I30999)
--	I30998 = NAND(I31000, I31001)
--	I31006 = NAND(I30982, I30998)
--	I31007 = NAND(I30982, I31006)
--	I31008 = NAND(I30998, I31006)
--	WX9982 = NAND(I31007, I31008)
--	I31087 = NAND(WX9631, WX9536)
--	I31088 = NAND(WX9631, I31087)
--	I31089 = NAND(WX9536, I31087)
--	WX10057 = NAND(I31088, I31089)
--	I31100 = NAND(WX9632, WX9538)
--	I31101 = NAND(WX9632, I31100)
--	I31102 = NAND(WX9538, I31100)
--	WX10064 = NAND(I31101, I31102)
--	I31113 = NAND(WX9633, WX9540)
--	I31114 = NAND(WX9633, I31113)
--	I31115 = NAND(WX9540, I31113)
--	WX10071 = NAND(I31114, I31115)
--	I31126 = NAND(WX9634, WX9542)
--	I31127 = NAND(WX9634, I31126)
--	I31128 = NAND(WX9542, I31126)
--	WX10078 = NAND(I31127, I31128)
--	I31139 = NAND(WX9635, WX9544)
--	I31140 = NAND(WX9635, I31139)
--	I31141 = NAND(WX9544, I31139)
--	WX10085 = NAND(I31140, I31141)
--	I31152 = NAND(WX9636, WX9546)
--	I31153 = NAND(WX9636, I31152)
--	I31154 = NAND(WX9546, I31152)
--	WX10092 = NAND(I31153, I31154)
--	I31165 = NAND(WX9637, WX9548)
--	I31166 = NAND(WX9637, I31165)
--	I31167 = NAND(WX9548, I31165)
--	WX10099 = NAND(I31166, I31167)
--	I31178 = NAND(WX9638, WX9550)
--	I31179 = NAND(WX9638, I31178)
--	I31180 = NAND(WX9550, I31178)
--	WX10106 = NAND(I31179, I31180)
--	I31191 = NAND(WX9639, WX9552)
--	I31192 = NAND(WX9639, I31191)
--	I31193 = NAND(WX9552, I31191)
--	WX10113 = NAND(I31192, I31193)
--	I31204 = NAND(WX9640, WX9554)
--	I31205 = NAND(WX9640, I31204)
--	I31206 = NAND(WX9554, I31204)
--	WX10120 = NAND(I31205, I31206)
--	I31217 = NAND(WX9641, WX9556)
--	I31218 = NAND(WX9641, I31217)
--	I31219 = NAND(WX9556, I31217)
--	WX10127 = NAND(I31218, I31219)
--	I31230 = NAND(WX9642, WX9558)
--	I31231 = NAND(WX9642, I31230)
--	I31232 = NAND(WX9558, I31230)
--	WX10134 = NAND(I31231, I31232)
--	I31243 = NAND(WX9643, WX9560)
--	I31244 = NAND(WX9643, I31243)
--	I31245 = NAND(WX9560, I31243)
--	WX10141 = NAND(I31244, I31245)
--	I31256 = NAND(WX9644, WX9562)
--	I31257 = NAND(WX9644, I31256)
--	I31258 = NAND(WX9562, I31256)
--	WX10148 = NAND(I31257, I31258)
--	I31269 = NAND(WX9645, WX9564)
--	I31270 = NAND(WX9645, I31269)
--	I31271 = NAND(WX9564, I31269)
--	WX10155 = NAND(I31270, I31271)
--	I31282 = NAND(WX9646, WX9566)
--	I31283 = NAND(WX9646, I31282)
--	I31284 = NAND(WX9566, I31282)
--	WX10162 = NAND(I31283, I31284)
--	I31295 = NAND(WX9647, WX9568)
--	I31296 = NAND(WX9647, I31295)
--	I31297 = NAND(WX9568, I31295)
--	WX10169 = NAND(I31296, I31297)
--	I31308 = NAND(WX9648, WX9570)
--	I31309 = NAND(WX9648, I31308)
--	I31310 = NAND(WX9570, I31308)
--	WX10176 = NAND(I31309, I31310)
--	I31321 = NAND(WX9649, WX9572)
--	I31322 = NAND(WX9649, I31321)
--	I31323 = NAND(WX9572, I31321)
--	WX10183 = NAND(I31322, I31323)
--	I31334 = NAND(WX9650, WX9574)
--	I31335 = NAND(WX9650, I31334)
--	I31336 = NAND(WX9574, I31334)
--	WX10190 = NAND(I31335, I31336)
--	I31347 = NAND(WX9651, WX9576)
--	I31348 = NAND(WX9651, I31347)
--	I31349 = NAND(WX9576, I31347)
--	WX10197 = NAND(I31348, I31349)
--	I31360 = NAND(WX9652, WX9578)
--	I31361 = NAND(WX9652, I31360)
--	I31362 = NAND(WX9578, I31360)
--	WX10204 = NAND(I31361, I31362)
--	I31373 = NAND(WX9653, WX9580)
--	I31374 = NAND(WX9653, I31373)
--	I31375 = NAND(WX9580, I31373)
--	WX10211 = NAND(I31374, I31375)
--	I31386 = NAND(WX9654, WX9582)
--	I31387 = NAND(WX9654, I31386)
--	I31388 = NAND(WX9582, I31386)
--	WX10218 = NAND(I31387, I31388)
--	I31399 = NAND(WX9655, WX9584)
--	I31400 = NAND(WX9655, I31399)
--	I31401 = NAND(WX9584, I31399)
--	WX10225 = NAND(I31400, I31401)
--	I31412 = NAND(WX9656, WX9586)
--	I31413 = NAND(WX9656, I31412)
--	I31414 = NAND(WX9586, I31412)
--	WX10232 = NAND(I31413, I31414)
--	I31425 = NAND(WX9657, WX9588)
--	I31426 = NAND(WX9657, I31425)
--	I31427 = NAND(WX9588, I31425)
--	WX10239 = NAND(I31426, I31427)
--	I31438 = NAND(WX9658, WX9590)
--	I31439 = NAND(WX9658, I31438)
--	I31440 = NAND(WX9590, I31438)
--	WX10246 = NAND(I31439, I31440)
--	I31451 = NAND(WX9659, WX9592)
--	I31452 = NAND(WX9659, I31451)
--	I31453 = NAND(WX9592, I31451)
--	WX10253 = NAND(I31452, I31453)
--	I31464 = NAND(WX9660, WX9594)
--	I31465 = NAND(WX9660, I31464)
--	I31466 = NAND(WX9594, I31464)
--	WX10260 = NAND(I31465, I31466)
--	I31477 = NAND(WX9661, WX9596)
--	I31478 = NAND(WX9661, I31477)
--	I31479 = NAND(WX9596, I31477)
--	WX10267 = NAND(I31478, I31479)
--	I31490 = NAND(WX9662, WX9598)
--	I31491 = NAND(WX9662, I31490)
--	I31492 = NAND(WX9598, I31490)
--	WX10274 = NAND(I31491, I31492)
--	I31505 = NAND(WX9678, CRC_OUT_2_31)
--	I31506 = NAND(WX9678, I31505)
--	I31507 = NAND(CRC_OUT_2_31, I31505)
--	I31504 = NAND(I31506, I31507)
--	I31512 = NAND(CRC_OUT_2_15, I31504)
--	I31513 = NAND(CRC_OUT_2_15, I31512)
--	I31514 = NAND(I31504, I31512)
--	WX10282 = NAND(I31513, I31514)
--	I31520 = NAND(WX9683, CRC_OUT_2_31)
--	I31521 = NAND(WX9683, I31520)
--	I31522 = NAND(CRC_OUT_2_31, I31520)
--	I31519 = NAND(I31521, I31522)
--	I31527 = NAND(CRC_OUT_2_10, I31519)
--	I31528 = NAND(CRC_OUT_2_10, I31527)
--	I31529 = NAND(I31519, I31527)
--	WX10283 = NAND(I31528, I31529)
--	I31535 = NAND(WX9690, CRC_OUT_2_31)
--	I31536 = NAND(WX9690, I31535)
--	I31537 = NAND(CRC_OUT_2_31, I31535)
--	I31534 = NAND(I31536, I31537)
--	I31542 = NAND(CRC_OUT_2_3, I31534)
--	I31543 = NAND(CRC_OUT_2_3, I31542)
--	I31544 = NAND(I31534, I31542)
--	WX10284 = NAND(I31543, I31544)
--	I31549 = NAND(WX9694, CRC_OUT_2_31)
--	I31550 = NAND(WX9694, I31549)
--	I31551 = NAND(CRC_OUT_2_31, I31549)
--	WX10285 = NAND(I31550, I31551)
--	I31556 = NAND(WX9663, CRC_OUT_2_30)
--	I31557 = NAND(WX9663, I31556)
--	I31558 = NAND(CRC_OUT_2_30, I31556)
--	WX10286 = NAND(I31557, I31558)
--	I31563 = NAND(WX9664, CRC_OUT_2_29)
--	I31564 = NAND(WX9664, I31563)
--	I31565 = NAND(CRC_OUT_2_29, I31563)
--	WX10287 = NAND(I31564, I31565)
--	I31570 = NAND(WX9665, CRC_OUT_2_28)
--	I31571 = NAND(WX9665, I31570)
--	I31572 = NAND(CRC_OUT_2_28, I31570)
--	WX10288 = NAND(I31571, I31572)
--	I31577 = NAND(WX9666, CRC_OUT_2_27)
--	I31578 = NAND(WX9666, I31577)
--	I31579 = NAND(CRC_OUT_2_27, I31577)
--	WX10289 = NAND(I31578, I31579)
--	I31584 = NAND(WX9667, CRC_OUT_2_26)
--	I31585 = NAND(WX9667, I31584)
--	I31586 = NAND(CRC_OUT_2_26, I31584)
--	WX10290 = NAND(I31585, I31586)
--	I31591 = NAND(WX9668, CRC_OUT_2_25)
--	I31592 = NAND(WX9668, I31591)
--	I31593 = NAND(CRC_OUT_2_25, I31591)
--	WX10291 = NAND(I31592, I31593)
--	I31598 = NAND(WX9669, CRC_OUT_2_24)
--	I31599 = NAND(WX9669, I31598)
--	I31600 = NAND(CRC_OUT_2_24, I31598)
--	WX10292 = NAND(I31599, I31600)
--	I31605 = NAND(WX9670, CRC_OUT_2_23)
--	I31606 = NAND(WX9670, I31605)
--	I31607 = NAND(CRC_OUT_2_23, I31605)
--	WX10293 = NAND(I31606, I31607)
--	I31612 = NAND(WX9671, CRC_OUT_2_22)
--	I31613 = NAND(WX9671, I31612)
--	I31614 = NAND(CRC_OUT_2_22, I31612)
--	WX10294 = NAND(I31613, I31614)
--	I31619 = NAND(WX9672, CRC_OUT_2_21)
--	I31620 = NAND(WX9672, I31619)
--	I31621 = NAND(CRC_OUT_2_21, I31619)
--	WX10295 = NAND(I31620, I31621)
--	I31626 = NAND(WX9673, CRC_OUT_2_20)
--	I31627 = NAND(WX9673, I31626)
--	I31628 = NAND(CRC_OUT_2_20, I31626)
--	WX10296 = NAND(I31627, I31628)
--	I31633 = NAND(WX9674, CRC_OUT_2_19)
--	I31634 = NAND(WX9674, I31633)
--	I31635 = NAND(CRC_OUT_2_19, I31633)
--	WX10297 = NAND(I31634, I31635)
--	I31640 = NAND(WX9675, CRC_OUT_2_18)
--	I31641 = NAND(WX9675, I31640)
--	I31642 = NAND(CRC_OUT_2_18, I31640)
--	WX10298 = NAND(I31641, I31642)
--	I31647 = NAND(WX9676, CRC_OUT_2_17)
--	I31648 = NAND(WX9676, I31647)
--	I31649 = NAND(CRC_OUT_2_17, I31647)
--	WX10299 = NAND(I31648, I31649)
--	I31654 = NAND(WX9677, CRC_OUT_2_16)
--	I31655 = NAND(WX9677, I31654)
--	I31656 = NAND(CRC_OUT_2_16, I31654)
--	WX10300 = NAND(I31655, I31656)
--	I31661 = NAND(WX9679, CRC_OUT_2_14)
--	I31662 = NAND(WX9679, I31661)
--	I31663 = NAND(CRC_OUT_2_14, I31661)
--	WX10301 = NAND(I31662, I31663)
--	I31668 = NAND(WX9680, CRC_OUT_2_13)
--	I31669 = NAND(WX9680, I31668)
--	I31670 = NAND(CRC_OUT_2_13, I31668)
--	WX10302 = NAND(I31669, I31670)
--	I31675 = NAND(WX9681, CRC_OUT_2_12)
--	I31676 = NAND(WX9681, I31675)
--	I31677 = NAND(CRC_OUT_2_12, I31675)
--	WX10303 = NAND(I31676, I31677)
--	I31682 = NAND(WX9682, CRC_OUT_2_11)
--	I31683 = NAND(WX9682, I31682)
--	I31684 = NAND(CRC_OUT_2_11, I31682)
--	WX10304 = NAND(I31683, I31684)
--	I31689 = NAND(WX9684, CRC_OUT_2_9)
--	I31690 = NAND(WX9684, I31689)
--	I31691 = NAND(CRC_OUT_2_9, I31689)
--	WX10305 = NAND(I31690, I31691)
--	I31696 = NAND(WX9685, CRC_OUT_2_8)
--	I31697 = NAND(WX9685, I31696)
--	I31698 = NAND(CRC_OUT_2_8, I31696)
--	WX10306 = NAND(I31697, I31698)
--	I31703 = NAND(WX9686, CRC_OUT_2_7)
--	I31704 = NAND(WX9686, I31703)
--	I31705 = NAND(CRC_OUT_2_7, I31703)
--	WX10307 = NAND(I31704, I31705)
--	I31710 = NAND(WX9687, CRC_OUT_2_6)
--	I31711 = NAND(WX9687, I31710)
--	I31712 = NAND(CRC_OUT_2_6, I31710)
--	WX10308 = NAND(I31711, I31712)
--	I31717 = NAND(WX9688, CRC_OUT_2_5)
--	I31718 = NAND(WX9688, I31717)
--	I31719 = NAND(CRC_OUT_2_5, I31717)
--	WX10309 = NAND(I31718, I31719)
--	I31724 = NAND(WX9689, CRC_OUT_2_4)
--	I31725 = NAND(WX9689, I31724)
--	I31726 = NAND(CRC_OUT_2_4, I31724)
--	WX10310 = NAND(I31725, I31726)
--	I31731 = NAND(WX9691, CRC_OUT_2_2)
--	I31732 = NAND(WX9691, I31731)
--	I31733 = NAND(CRC_OUT_2_2, I31731)
--	WX10311 = NAND(I31732, I31733)
--	I31738 = NAND(WX9692, CRC_OUT_2_1)
--	I31739 = NAND(WX9692, I31738)
--	I31740 = NAND(CRC_OUT_2_1, I31738)
--	WX10312 = NAND(I31739, I31740)
--	I31745 = NAND(WX9693, CRC_OUT_2_0)
--	I31746 = NAND(WX9693, I31745)
--	I31747 = NAND(CRC_OUT_2_0, I31745)
--	WX10313 = NAND(I31746, I31747)
--	I34028 = NAND(WX11345, WX10989)
--	I34029 = NAND(WX11345, I34028)
--	I34030 = NAND(WX10989, I34028)
--	I34027 = NAND(I34029, I34030)
--	I34035 = NAND(WX11053, I34027)
--	I34036 = NAND(WX11053, I34035)
--	I34037 = NAND(I34027, I34035)
--	I34026 = NAND(I34036, I34037)
--	I34043 = NAND(WX11117, WX11181)
--	I34044 = NAND(WX11117, I34043)
--	I34045 = NAND(WX11181, I34043)
--	I34042 = NAND(I34044, I34045)
--	I34050 = NAND(I34026, I34042)
--	I34051 = NAND(I34026, I34050)
--	I34052 = NAND(I34042, I34050)
--	WX11244 = NAND(I34051, I34052)
--	I34059 = NAND(WX11345, WX10991)
--	I34060 = NAND(WX11345, I34059)
--	I34061 = NAND(WX10991, I34059)
--	I34058 = NAND(I34060, I34061)
--	I34066 = NAND(WX11055, I34058)
--	I34067 = NAND(WX11055, I34066)
--	I34068 = NAND(I34058, I34066)
--	I34057 = NAND(I34067, I34068)
--	I34074 = NAND(WX11119, WX11183)
--	I34075 = NAND(WX11119, I34074)
--	I34076 = NAND(WX11183, I34074)
--	I34073 = NAND(I34075, I34076)
--	I34081 = NAND(I34057, I34073)
--	I34082 = NAND(I34057, I34081)
--	I34083 = NAND(I34073, I34081)
--	WX11245 = NAND(I34082, I34083)
--	I34090 = NAND(WX11345, WX10993)
--	I34091 = NAND(WX11345, I34090)
--	I34092 = NAND(WX10993, I34090)
--	I34089 = NAND(I34091, I34092)
--	I34097 = NAND(WX11057, I34089)
--	I34098 = NAND(WX11057, I34097)
--	I34099 = NAND(I34089, I34097)
--	I34088 = NAND(I34098, I34099)
--	I34105 = NAND(WX11121, WX11185)
--	I34106 = NAND(WX11121, I34105)
--	I34107 = NAND(WX11185, I34105)
--	I34104 = NAND(I34106, I34107)
--	I34112 = NAND(I34088, I34104)
--	I34113 = NAND(I34088, I34112)
--	I34114 = NAND(I34104, I34112)
--	WX11246 = NAND(I34113, I34114)
--	I34121 = NAND(WX11345, WX10995)
--	I34122 = NAND(WX11345, I34121)
--	I34123 = NAND(WX10995, I34121)
--	I34120 = NAND(I34122, I34123)
--	I34128 = NAND(WX11059, I34120)
--	I34129 = NAND(WX11059, I34128)
--	I34130 = NAND(I34120, I34128)
--	I34119 = NAND(I34129, I34130)
--	I34136 = NAND(WX11123, WX11187)
--	I34137 = NAND(WX11123, I34136)
--	I34138 = NAND(WX11187, I34136)
--	I34135 = NAND(I34137, I34138)
--	I34143 = NAND(I34119, I34135)
--	I34144 = NAND(I34119, I34143)
--	I34145 = NAND(I34135, I34143)
--	WX11247 = NAND(I34144, I34145)
--	I34152 = NAND(WX11345, WX10997)
--	I34153 = NAND(WX11345, I34152)
--	I34154 = NAND(WX10997, I34152)
--	I34151 = NAND(I34153, I34154)
--	I34159 = NAND(WX11061, I34151)
--	I34160 = NAND(WX11061, I34159)
--	I34161 = NAND(I34151, I34159)
--	I34150 = NAND(I34160, I34161)
--	I34167 = NAND(WX11125, WX11189)
--	I34168 = NAND(WX11125, I34167)
--	I34169 = NAND(WX11189, I34167)
--	I34166 = NAND(I34168, I34169)
--	I34174 = NAND(I34150, I34166)
--	I34175 = NAND(I34150, I34174)
--	I34176 = NAND(I34166, I34174)
--	WX11248 = NAND(I34175, I34176)
--	I34183 = NAND(WX11345, WX10999)
--	I34184 = NAND(WX11345, I34183)
--	I34185 = NAND(WX10999, I34183)
--	I34182 = NAND(I34184, I34185)
--	I34190 = NAND(WX11063, I34182)
--	I34191 = NAND(WX11063, I34190)
--	I34192 = NAND(I34182, I34190)
--	I34181 = NAND(I34191, I34192)
--	I34198 = NAND(WX11127, WX11191)
--	I34199 = NAND(WX11127, I34198)
--	I34200 = NAND(WX11191, I34198)
--	I34197 = NAND(I34199, I34200)
--	I34205 = NAND(I34181, I34197)
--	I34206 = NAND(I34181, I34205)
--	I34207 = NAND(I34197, I34205)
--	WX11249 = NAND(I34206, I34207)
--	I34214 = NAND(WX11345, WX11001)
--	I34215 = NAND(WX11345, I34214)
--	I34216 = NAND(WX11001, I34214)
--	I34213 = NAND(I34215, I34216)
--	I34221 = NAND(WX11065, I34213)
--	I34222 = NAND(WX11065, I34221)
--	I34223 = NAND(I34213, I34221)
--	I34212 = NAND(I34222, I34223)
--	I34229 = NAND(WX11129, WX11193)
--	I34230 = NAND(WX11129, I34229)
--	I34231 = NAND(WX11193, I34229)
--	I34228 = NAND(I34230, I34231)
--	I34236 = NAND(I34212, I34228)
--	I34237 = NAND(I34212, I34236)
--	I34238 = NAND(I34228, I34236)
--	WX11250 = NAND(I34237, I34238)
--	I34245 = NAND(WX11345, WX11003)
--	I34246 = NAND(WX11345, I34245)
--	I34247 = NAND(WX11003, I34245)
--	I34244 = NAND(I34246, I34247)
--	I34252 = NAND(WX11067, I34244)
--	I34253 = NAND(WX11067, I34252)
--	I34254 = NAND(I34244, I34252)
--	I34243 = NAND(I34253, I34254)
--	I34260 = NAND(WX11131, WX11195)
--	I34261 = NAND(WX11131, I34260)
--	I34262 = NAND(WX11195, I34260)
--	I34259 = NAND(I34261, I34262)
--	I34267 = NAND(I34243, I34259)
--	I34268 = NAND(I34243, I34267)
--	I34269 = NAND(I34259, I34267)
--	WX11251 = NAND(I34268, I34269)
--	I34276 = NAND(WX11345, WX11005)
--	I34277 = NAND(WX11345, I34276)
--	I34278 = NAND(WX11005, I34276)
--	I34275 = NAND(I34277, I34278)
--	I34283 = NAND(WX11069, I34275)
--	I34284 = NAND(WX11069, I34283)
--	I34285 = NAND(I34275, I34283)
--	I34274 = NAND(I34284, I34285)
--	I34291 = NAND(WX11133, WX11197)
--	I34292 = NAND(WX11133, I34291)
--	I34293 = NAND(WX11197, I34291)
--	I34290 = NAND(I34292, I34293)
--	I34298 = NAND(I34274, I34290)
--	I34299 = NAND(I34274, I34298)
--	I34300 = NAND(I34290, I34298)
--	WX11252 = NAND(I34299, I34300)
--	I34307 = NAND(WX11345, WX11007)
--	I34308 = NAND(WX11345, I34307)
--	I34309 = NAND(WX11007, I34307)
--	I34306 = NAND(I34308, I34309)
--	I34314 = NAND(WX11071, I34306)
--	I34315 = NAND(WX11071, I34314)
--	I34316 = NAND(I34306, I34314)
--	I34305 = NAND(I34315, I34316)
--	I34322 = NAND(WX11135, WX11199)
--	I34323 = NAND(WX11135, I34322)
--	I34324 = NAND(WX11199, I34322)
--	I34321 = NAND(I34323, I34324)
--	I34329 = NAND(I34305, I34321)
--	I34330 = NAND(I34305, I34329)
--	I34331 = NAND(I34321, I34329)
--	WX11253 = NAND(I34330, I34331)
--	I34338 = NAND(WX11345, WX11009)
--	I34339 = NAND(WX11345, I34338)
--	I34340 = NAND(WX11009, I34338)
--	I34337 = NAND(I34339, I34340)
--	I34345 = NAND(WX11073, I34337)
--	I34346 = NAND(WX11073, I34345)
--	I34347 = NAND(I34337, I34345)
--	I34336 = NAND(I34346, I34347)
--	I34353 = NAND(WX11137, WX11201)
--	I34354 = NAND(WX11137, I34353)
--	I34355 = NAND(WX11201, I34353)
--	I34352 = NAND(I34354, I34355)
--	I34360 = NAND(I34336, I34352)
--	I34361 = NAND(I34336, I34360)
--	I34362 = NAND(I34352, I34360)
--	WX11254 = NAND(I34361, I34362)
--	I34369 = NAND(WX11345, WX11011)
--	I34370 = NAND(WX11345, I34369)
--	I34371 = NAND(WX11011, I34369)
--	I34368 = NAND(I34370, I34371)
--	I34376 = NAND(WX11075, I34368)
--	I34377 = NAND(WX11075, I34376)
--	I34378 = NAND(I34368, I34376)
--	I34367 = NAND(I34377, I34378)
--	I34384 = NAND(WX11139, WX11203)
--	I34385 = NAND(WX11139, I34384)
--	I34386 = NAND(WX11203, I34384)
--	I34383 = NAND(I34385, I34386)
--	I34391 = NAND(I34367, I34383)
--	I34392 = NAND(I34367, I34391)
--	I34393 = NAND(I34383, I34391)
--	WX11255 = NAND(I34392, I34393)
--	I34400 = NAND(WX11345, WX11013)
--	I34401 = NAND(WX11345, I34400)
--	I34402 = NAND(WX11013, I34400)
--	I34399 = NAND(I34401, I34402)
--	I34407 = NAND(WX11077, I34399)
--	I34408 = NAND(WX11077, I34407)
--	I34409 = NAND(I34399, I34407)
--	I34398 = NAND(I34408, I34409)
--	I34415 = NAND(WX11141, WX11205)
--	I34416 = NAND(WX11141, I34415)
--	I34417 = NAND(WX11205, I34415)
--	I34414 = NAND(I34416, I34417)
--	I34422 = NAND(I34398, I34414)
--	I34423 = NAND(I34398, I34422)
--	I34424 = NAND(I34414, I34422)
--	WX11256 = NAND(I34423, I34424)
--	I34431 = NAND(WX11345, WX11015)
--	I34432 = NAND(WX11345, I34431)
--	I34433 = NAND(WX11015, I34431)
--	I34430 = NAND(I34432, I34433)
--	I34438 = NAND(WX11079, I34430)
--	I34439 = NAND(WX11079, I34438)
--	I34440 = NAND(I34430, I34438)
--	I34429 = NAND(I34439, I34440)
--	I34446 = NAND(WX11143, WX11207)
--	I34447 = NAND(WX11143, I34446)
--	I34448 = NAND(WX11207, I34446)
--	I34445 = NAND(I34447, I34448)
--	I34453 = NAND(I34429, I34445)
--	I34454 = NAND(I34429, I34453)
--	I34455 = NAND(I34445, I34453)
--	WX11257 = NAND(I34454, I34455)
--	I34462 = NAND(WX11345, WX11017)
--	I34463 = NAND(WX11345, I34462)
--	I34464 = NAND(WX11017, I34462)
--	I34461 = NAND(I34463, I34464)
--	I34469 = NAND(WX11081, I34461)
--	I34470 = NAND(WX11081, I34469)
--	I34471 = NAND(I34461, I34469)
--	I34460 = NAND(I34470, I34471)
--	I34477 = NAND(WX11145, WX11209)
--	I34478 = NAND(WX11145, I34477)
--	I34479 = NAND(WX11209, I34477)
--	I34476 = NAND(I34478, I34479)
--	I34484 = NAND(I34460, I34476)
--	I34485 = NAND(I34460, I34484)
--	I34486 = NAND(I34476, I34484)
--	WX11258 = NAND(I34485, I34486)
--	I34493 = NAND(WX11345, WX11019)
--	I34494 = NAND(WX11345, I34493)
--	I34495 = NAND(WX11019, I34493)
--	I34492 = NAND(I34494, I34495)
--	I34500 = NAND(WX11083, I34492)
--	I34501 = NAND(WX11083, I34500)
--	I34502 = NAND(I34492, I34500)
--	I34491 = NAND(I34501, I34502)
--	I34508 = NAND(WX11147, WX11211)
--	I34509 = NAND(WX11147, I34508)
--	I34510 = NAND(WX11211, I34508)
--	I34507 = NAND(I34509, I34510)
--	I34515 = NAND(I34491, I34507)
--	I34516 = NAND(I34491, I34515)
--	I34517 = NAND(I34507, I34515)
--	WX11259 = NAND(I34516, I34517)
--	I34524 = NAND(WX11346, WX11021)
--	I34525 = NAND(WX11346, I34524)
--	I34526 = NAND(WX11021, I34524)
--	I34523 = NAND(I34525, I34526)
--	I34531 = NAND(WX11085, I34523)
--	I34532 = NAND(WX11085, I34531)
--	I34533 = NAND(I34523, I34531)
--	I34522 = NAND(I34532, I34533)
--	I34539 = NAND(WX11149, WX11213)
--	I34540 = NAND(WX11149, I34539)
--	I34541 = NAND(WX11213, I34539)
--	I34538 = NAND(I34540, I34541)
--	I34546 = NAND(I34522, I34538)
--	I34547 = NAND(I34522, I34546)
--	I34548 = NAND(I34538, I34546)
--	WX11260 = NAND(I34547, I34548)
--	I34555 = NAND(WX11346, WX11023)
--	I34556 = NAND(WX11346, I34555)
--	I34557 = NAND(WX11023, I34555)
--	I34554 = NAND(I34556, I34557)
--	I34562 = NAND(WX11087, I34554)
--	I34563 = NAND(WX11087, I34562)
--	I34564 = NAND(I34554, I34562)
--	I34553 = NAND(I34563, I34564)
--	I34570 = NAND(WX11151, WX11215)
--	I34571 = NAND(WX11151, I34570)
--	I34572 = NAND(WX11215, I34570)
--	I34569 = NAND(I34571, I34572)
--	I34577 = NAND(I34553, I34569)
--	I34578 = NAND(I34553, I34577)
--	I34579 = NAND(I34569, I34577)
--	WX11261 = NAND(I34578, I34579)
--	I34586 = NAND(WX11346, WX11025)
--	I34587 = NAND(WX11346, I34586)
--	I34588 = NAND(WX11025, I34586)
--	I34585 = NAND(I34587, I34588)
--	I34593 = NAND(WX11089, I34585)
--	I34594 = NAND(WX11089, I34593)
--	I34595 = NAND(I34585, I34593)
--	I34584 = NAND(I34594, I34595)
--	I34601 = NAND(WX11153, WX11217)
--	I34602 = NAND(WX11153, I34601)
--	I34603 = NAND(WX11217, I34601)
--	I34600 = NAND(I34602, I34603)
--	I34608 = NAND(I34584, I34600)
--	I34609 = NAND(I34584, I34608)
--	I34610 = NAND(I34600, I34608)
--	WX11262 = NAND(I34609, I34610)
--	I34617 = NAND(WX11346, WX11027)
--	I34618 = NAND(WX11346, I34617)
--	I34619 = NAND(WX11027, I34617)
--	I34616 = NAND(I34618, I34619)
--	I34624 = NAND(WX11091, I34616)
--	I34625 = NAND(WX11091, I34624)
--	I34626 = NAND(I34616, I34624)
--	I34615 = NAND(I34625, I34626)
--	I34632 = NAND(WX11155, WX11219)
--	I34633 = NAND(WX11155, I34632)
--	I34634 = NAND(WX11219, I34632)
--	I34631 = NAND(I34633, I34634)
--	I34639 = NAND(I34615, I34631)
--	I34640 = NAND(I34615, I34639)
--	I34641 = NAND(I34631, I34639)
--	WX11263 = NAND(I34640, I34641)
--	I34648 = NAND(WX11346, WX11029)
--	I34649 = NAND(WX11346, I34648)
--	I34650 = NAND(WX11029, I34648)
--	I34647 = NAND(I34649, I34650)
--	I34655 = NAND(WX11093, I34647)
--	I34656 = NAND(WX11093, I34655)
--	I34657 = NAND(I34647, I34655)
--	I34646 = NAND(I34656, I34657)
--	I34663 = NAND(WX11157, WX11221)
--	I34664 = NAND(WX11157, I34663)
--	I34665 = NAND(WX11221, I34663)
--	I34662 = NAND(I34664, I34665)
--	I34670 = NAND(I34646, I34662)
--	I34671 = NAND(I34646, I34670)
--	I34672 = NAND(I34662, I34670)
--	WX11264 = NAND(I34671, I34672)
--	I34679 = NAND(WX11346, WX11031)
--	I34680 = NAND(WX11346, I34679)
--	I34681 = NAND(WX11031, I34679)
--	I34678 = NAND(I34680, I34681)
--	I34686 = NAND(WX11095, I34678)
--	I34687 = NAND(WX11095, I34686)
--	I34688 = NAND(I34678, I34686)
--	I34677 = NAND(I34687, I34688)
--	I34694 = NAND(WX11159, WX11223)
--	I34695 = NAND(WX11159, I34694)
--	I34696 = NAND(WX11223, I34694)
--	I34693 = NAND(I34695, I34696)
--	I34701 = NAND(I34677, I34693)
--	I34702 = NAND(I34677, I34701)
--	I34703 = NAND(I34693, I34701)
--	WX11265 = NAND(I34702, I34703)
--	I34710 = NAND(WX11346, WX11033)
--	I34711 = NAND(WX11346, I34710)
--	I34712 = NAND(WX11033, I34710)
--	I34709 = NAND(I34711, I34712)
--	I34717 = NAND(WX11097, I34709)
--	I34718 = NAND(WX11097, I34717)
--	I34719 = NAND(I34709, I34717)
--	I34708 = NAND(I34718, I34719)
--	I34725 = NAND(WX11161, WX11225)
--	I34726 = NAND(WX11161, I34725)
--	I34727 = NAND(WX11225, I34725)
--	I34724 = NAND(I34726, I34727)
--	I34732 = NAND(I34708, I34724)
--	I34733 = NAND(I34708, I34732)
--	I34734 = NAND(I34724, I34732)
--	WX11266 = NAND(I34733, I34734)
--	I34741 = NAND(WX11346, WX11035)
--	I34742 = NAND(WX11346, I34741)
--	I34743 = NAND(WX11035, I34741)
--	I34740 = NAND(I34742, I34743)
--	I34748 = NAND(WX11099, I34740)
--	I34749 = NAND(WX11099, I34748)
--	I34750 = NAND(I34740, I34748)
--	I34739 = NAND(I34749, I34750)
--	I34756 = NAND(WX11163, WX11227)
--	I34757 = NAND(WX11163, I34756)
--	I34758 = NAND(WX11227, I34756)
--	I34755 = NAND(I34757, I34758)
--	I34763 = NAND(I34739, I34755)
--	I34764 = NAND(I34739, I34763)
--	I34765 = NAND(I34755, I34763)
--	WX11267 = NAND(I34764, I34765)
--	I34772 = NAND(WX11346, WX11037)
--	I34773 = NAND(WX11346, I34772)
--	I34774 = NAND(WX11037, I34772)
--	I34771 = NAND(I34773, I34774)
--	I34779 = NAND(WX11101, I34771)
--	I34780 = NAND(WX11101, I34779)
--	I34781 = NAND(I34771, I34779)
--	I34770 = NAND(I34780, I34781)
--	I34787 = NAND(WX11165, WX11229)
--	I34788 = NAND(WX11165, I34787)
--	I34789 = NAND(WX11229, I34787)
--	I34786 = NAND(I34788, I34789)
--	I34794 = NAND(I34770, I34786)
--	I34795 = NAND(I34770, I34794)
--	I34796 = NAND(I34786, I34794)
--	WX11268 = NAND(I34795, I34796)
--	I34803 = NAND(WX11346, WX11039)
--	I34804 = NAND(WX11346, I34803)
--	I34805 = NAND(WX11039, I34803)
--	I34802 = NAND(I34804, I34805)
--	I34810 = NAND(WX11103, I34802)
--	I34811 = NAND(WX11103, I34810)
--	I34812 = NAND(I34802, I34810)
--	I34801 = NAND(I34811, I34812)
--	I34818 = NAND(WX11167, WX11231)
--	I34819 = NAND(WX11167, I34818)
--	I34820 = NAND(WX11231, I34818)
--	I34817 = NAND(I34819, I34820)
--	I34825 = NAND(I34801, I34817)
--	I34826 = NAND(I34801, I34825)
--	I34827 = NAND(I34817, I34825)
--	WX11269 = NAND(I34826, I34827)
--	I34834 = NAND(WX11346, WX11041)
--	I34835 = NAND(WX11346, I34834)
--	I34836 = NAND(WX11041, I34834)
--	I34833 = NAND(I34835, I34836)
--	I34841 = NAND(WX11105, I34833)
--	I34842 = NAND(WX11105, I34841)
--	I34843 = NAND(I34833, I34841)
--	I34832 = NAND(I34842, I34843)
--	I34849 = NAND(WX11169, WX11233)
--	I34850 = NAND(WX11169, I34849)
--	I34851 = NAND(WX11233, I34849)
--	I34848 = NAND(I34850, I34851)
--	I34856 = NAND(I34832, I34848)
--	I34857 = NAND(I34832, I34856)
--	I34858 = NAND(I34848, I34856)
--	WX11270 = NAND(I34857, I34858)
--	I34865 = NAND(WX11346, WX11043)
--	I34866 = NAND(WX11346, I34865)
--	I34867 = NAND(WX11043, I34865)
--	I34864 = NAND(I34866, I34867)
--	I34872 = NAND(WX11107, I34864)
--	I34873 = NAND(WX11107, I34872)
--	I34874 = NAND(I34864, I34872)
--	I34863 = NAND(I34873, I34874)
--	I34880 = NAND(WX11171, WX11235)
--	I34881 = NAND(WX11171, I34880)
--	I34882 = NAND(WX11235, I34880)
--	I34879 = NAND(I34881, I34882)
--	I34887 = NAND(I34863, I34879)
--	I34888 = NAND(I34863, I34887)
--	I34889 = NAND(I34879, I34887)
--	WX11271 = NAND(I34888, I34889)
--	I34896 = NAND(WX11346, WX11045)
--	I34897 = NAND(WX11346, I34896)
--	I34898 = NAND(WX11045, I34896)
--	I34895 = NAND(I34897, I34898)
--	I34903 = NAND(WX11109, I34895)
--	I34904 = NAND(WX11109, I34903)
--	I34905 = NAND(I34895, I34903)
--	I34894 = NAND(I34904, I34905)
--	I34911 = NAND(WX11173, WX11237)
--	I34912 = NAND(WX11173, I34911)
--	I34913 = NAND(WX11237, I34911)
--	I34910 = NAND(I34912, I34913)
--	I34918 = NAND(I34894, I34910)
--	I34919 = NAND(I34894, I34918)
--	I34920 = NAND(I34910, I34918)
--	WX11272 = NAND(I34919, I34920)
--	I34927 = NAND(WX11346, WX11047)
--	I34928 = NAND(WX11346, I34927)
--	I34929 = NAND(WX11047, I34927)
--	I34926 = NAND(I34928, I34929)
--	I34934 = NAND(WX11111, I34926)
--	I34935 = NAND(WX11111, I34934)
--	I34936 = NAND(I34926, I34934)
--	I34925 = NAND(I34935, I34936)
--	I34942 = NAND(WX11175, WX11239)
--	I34943 = NAND(WX11175, I34942)
--	I34944 = NAND(WX11239, I34942)
--	I34941 = NAND(I34943, I34944)
--	I34949 = NAND(I34925, I34941)
--	I34950 = NAND(I34925, I34949)
--	I34951 = NAND(I34941, I34949)
--	WX11273 = NAND(I34950, I34951)
--	I34958 = NAND(WX11346, WX11049)
--	I34959 = NAND(WX11346, I34958)
--	I34960 = NAND(WX11049, I34958)
--	I34957 = NAND(I34959, I34960)
--	I34965 = NAND(WX11113, I34957)
--	I34966 = NAND(WX11113, I34965)
--	I34967 = NAND(I34957, I34965)
--	I34956 = NAND(I34966, I34967)
--	I34973 = NAND(WX11177, WX11241)
--	I34974 = NAND(WX11177, I34973)
--	I34975 = NAND(WX11241, I34973)
--	I34972 = NAND(I34974, I34975)
--	I34980 = NAND(I34956, I34972)
--	I34981 = NAND(I34956, I34980)
--	I34982 = NAND(I34972, I34980)
--	WX11274 = NAND(I34981, I34982)
--	I34989 = NAND(WX11346, WX11051)
--	I34990 = NAND(WX11346, I34989)
--	I34991 = NAND(WX11051, I34989)
--	I34988 = NAND(I34990, I34991)
--	I34996 = NAND(WX11115, I34988)
--	I34997 = NAND(WX11115, I34996)
--	I34998 = NAND(I34988, I34996)
--	I34987 = NAND(I34997, I34998)
--	I35004 = NAND(WX11179, WX11243)
--	I35005 = NAND(WX11179, I35004)
--	I35006 = NAND(WX11243, I35004)
--	I35003 = NAND(I35005, I35006)
--	I35011 = NAND(I34987, I35003)
--	I35012 = NAND(I34987, I35011)
--	I35013 = NAND(I35003, I35011)
--	WX11275 = NAND(I35012, I35013)
--	I35092 = NAND(WX10924, WX10829)
--	I35093 = NAND(WX10924, I35092)
--	I35094 = NAND(WX10829, I35092)
--	WX11350 = NAND(I35093, I35094)
--	I35105 = NAND(WX10925, WX10831)
--	I35106 = NAND(WX10925, I35105)
--	I35107 = NAND(WX10831, I35105)
--	WX11357 = NAND(I35106, I35107)
--	I35118 = NAND(WX10926, WX10833)
--	I35119 = NAND(WX10926, I35118)
--	I35120 = NAND(WX10833, I35118)
--	WX11364 = NAND(I35119, I35120)
--	I35131 = NAND(WX10927, WX10835)
--	I35132 = NAND(WX10927, I35131)
--	I35133 = NAND(WX10835, I35131)
--	WX11371 = NAND(I35132, I35133)
--	I35144 = NAND(WX10928, WX10837)
--	I35145 = NAND(WX10928, I35144)
--	I35146 = NAND(WX10837, I35144)
--	WX11378 = NAND(I35145, I35146)
--	I35157 = NAND(WX10929, WX10839)
--	I35158 = NAND(WX10929, I35157)
--	I35159 = NAND(WX10839, I35157)
--	WX11385 = NAND(I35158, I35159)
--	I35170 = NAND(WX10930, WX10841)
--	I35171 = NAND(WX10930, I35170)
--	I35172 = NAND(WX10841, I35170)
--	WX11392 = NAND(I35171, I35172)
--	I35183 = NAND(WX10931, WX10843)
--	I35184 = NAND(WX10931, I35183)
--	I35185 = NAND(WX10843, I35183)
--	WX11399 = NAND(I35184, I35185)
--	I35196 = NAND(WX10932, WX10845)
--	I35197 = NAND(WX10932, I35196)
--	I35198 = NAND(WX10845, I35196)
--	WX11406 = NAND(I35197, I35198)
--	I35209 = NAND(WX10933, WX10847)
--	I35210 = NAND(WX10933, I35209)
--	I35211 = NAND(WX10847, I35209)
--	WX11413 = NAND(I35210, I35211)
--	I35222 = NAND(WX10934, WX10849)
--	I35223 = NAND(WX10934, I35222)
--	I35224 = NAND(WX10849, I35222)
--	WX11420 = NAND(I35223, I35224)
--	I35235 = NAND(WX10935, WX10851)
--	I35236 = NAND(WX10935, I35235)
--	I35237 = NAND(WX10851, I35235)
--	WX11427 = NAND(I35236, I35237)
--	I35248 = NAND(WX10936, WX10853)
--	I35249 = NAND(WX10936, I35248)
--	I35250 = NAND(WX10853, I35248)
--	WX11434 = NAND(I35249, I35250)
--	I35261 = NAND(WX10937, WX10855)
--	I35262 = NAND(WX10937, I35261)
--	I35263 = NAND(WX10855, I35261)
--	WX11441 = NAND(I35262, I35263)
--	I35274 = NAND(WX10938, WX10857)
--	I35275 = NAND(WX10938, I35274)
--	I35276 = NAND(WX10857, I35274)
--	WX11448 = NAND(I35275, I35276)
--	I35287 = NAND(WX10939, WX10859)
--	I35288 = NAND(WX10939, I35287)
--	I35289 = NAND(WX10859, I35287)
--	WX11455 = NAND(I35288, I35289)
--	I35300 = NAND(WX10940, WX10861)
--	I35301 = NAND(WX10940, I35300)
--	I35302 = NAND(WX10861, I35300)
--	WX11462 = NAND(I35301, I35302)
--	I35313 = NAND(WX10941, WX10863)
--	I35314 = NAND(WX10941, I35313)
--	I35315 = NAND(WX10863, I35313)
--	WX11469 = NAND(I35314, I35315)
--	I35326 = NAND(WX10942, WX10865)
--	I35327 = NAND(WX10942, I35326)
--	I35328 = NAND(WX10865, I35326)
--	WX11476 = NAND(I35327, I35328)
--	I35339 = NAND(WX10943, WX10867)
--	I35340 = NAND(WX10943, I35339)
--	I35341 = NAND(WX10867, I35339)
--	WX11483 = NAND(I35340, I35341)
--	I35352 = NAND(WX10944, WX10869)
--	I35353 = NAND(WX10944, I35352)
--	I35354 = NAND(WX10869, I35352)
--	WX11490 = NAND(I35353, I35354)
--	I35365 = NAND(WX10945, WX10871)
--	I35366 = NAND(WX10945, I35365)
--	I35367 = NAND(WX10871, I35365)
--	WX11497 = NAND(I35366, I35367)
--	I35378 = NAND(WX10946, WX10873)
--	I35379 = NAND(WX10946, I35378)
--	I35380 = NAND(WX10873, I35378)
--	WX11504 = NAND(I35379, I35380)
--	I35391 = NAND(WX10947, WX10875)
--	I35392 = NAND(WX10947, I35391)
--	I35393 = NAND(WX10875, I35391)
--	WX11511 = NAND(I35392, I35393)
--	I35404 = NAND(WX10948, WX10877)
--	I35405 = NAND(WX10948, I35404)
--	I35406 = NAND(WX10877, I35404)
--	WX11518 = NAND(I35405, I35406)
--	I35417 = NAND(WX10949, WX10879)
--	I35418 = NAND(WX10949, I35417)
--	I35419 = NAND(WX10879, I35417)
--	WX11525 = NAND(I35418, I35419)
--	I35430 = NAND(WX10950, WX10881)
--	I35431 = NAND(WX10950, I35430)
--	I35432 = NAND(WX10881, I35430)
--	WX11532 = NAND(I35431, I35432)
--	I35443 = NAND(WX10951, WX10883)
--	I35444 = NAND(WX10951, I35443)
--	I35445 = NAND(WX10883, I35443)
--	WX11539 = NAND(I35444, I35445)
--	I35456 = NAND(WX10952, WX10885)
--	I35457 = NAND(WX10952, I35456)
--	I35458 = NAND(WX10885, I35456)
--	WX11546 = NAND(I35457, I35458)
--	I35469 = NAND(WX10953, WX10887)
--	I35470 = NAND(WX10953, I35469)
--	I35471 = NAND(WX10887, I35469)
--	WX11553 = NAND(I35470, I35471)
--	I35482 = NAND(WX10954, WX10889)
--	I35483 = NAND(WX10954, I35482)
--	I35484 = NAND(WX10889, I35482)
--	WX11560 = NAND(I35483, I35484)
--	I35495 = NAND(WX10955, WX10891)
--	I35496 = NAND(WX10955, I35495)
--	I35497 = NAND(WX10891, I35495)
--	WX11567 = NAND(I35496, I35497)
--	I35510 = NAND(WX10971, CRC_OUT_1_31)
--	I35511 = NAND(WX10971, I35510)
--	I35512 = NAND(CRC_OUT_1_31, I35510)
--	I35509 = NAND(I35511, I35512)
--	I35517 = NAND(CRC_OUT_1_15, I35509)
--	I35518 = NAND(CRC_OUT_1_15, I35517)
--	I35519 = NAND(I35509, I35517)
--	WX11575 = NAND(I35518, I35519)
--	I35525 = NAND(WX10976, CRC_OUT_1_31)
--	I35526 = NAND(WX10976, I35525)
--	I35527 = NAND(CRC_OUT_1_31, I35525)
--	I35524 = NAND(I35526, I35527)
--	I35532 = NAND(CRC_OUT_1_10, I35524)
--	I35533 = NAND(CRC_OUT_1_10, I35532)
--	I35534 = NAND(I35524, I35532)
--	WX11576 = NAND(I35533, I35534)
--	I35540 = NAND(WX10983, CRC_OUT_1_31)
--	I35541 = NAND(WX10983, I35540)
--	I35542 = NAND(CRC_OUT_1_31, I35540)
--	I35539 = NAND(I35541, I35542)
--	I35547 = NAND(CRC_OUT_1_3, I35539)
--	I35548 = NAND(CRC_OUT_1_3, I35547)
--	I35549 = NAND(I35539, I35547)
--	WX11577 = NAND(I35548, I35549)
--	I35554 = NAND(WX10987, CRC_OUT_1_31)
--	I35555 = NAND(WX10987, I35554)
--	I35556 = NAND(CRC_OUT_1_31, I35554)
--	WX11578 = NAND(I35555, I35556)
--	I35561 = NAND(WX10956, CRC_OUT_1_30)
--	I35562 = NAND(WX10956, I35561)
--	I35563 = NAND(CRC_OUT_1_30, I35561)
--	WX11579 = NAND(I35562, I35563)
--	I35568 = NAND(WX10957, CRC_OUT_1_29)
--	I35569 = NAND(WX10957, I35568)
--	I35570 = NAND(CRC_OUT_1_29, I35568)
--	WX11580 = NAND(I35569, I35570)
--	I35575 = NAND(WX10958, CRC_OUT_1_28)
--	I35576 = NAND(WX10958, I35575)
--	I35577 = NAND(CRC_OUT_1_28, I35575)
--	WX11581 = NAND(I35576, I35577)
--	I35582 = NAND(WX10959, CRC_OUT_1_27)
--	I35583 = NAND(WX10959, I35582)
--	I35584 = NAND(CRC_OUT_1_27, I35582)
--	WX11582 = NAND(I35583, I35584)
--	I35589 = NAND(WX10960, CRC_OUT_1_26)
--	I35590 = NAND(WX10960, I35589)
--	I35591 = NAND(CRC_OUT_1_26, I35589)
--	WX11583 = NAND(I35590, I35591)
--	I35596 = NAND(WX10961, CRC_OUT_1_25)
--	I35597 = NAND(WX10961, I35596)
--	I35598 = NAND(CRC_OUT_1_25, I35596)
--	WX11584 = NAND(I35597, I35598)
--	I35603 = NAND(WX10962, CRC_OUT_1_24)
--	I35604 = NAND(WX10962, I35603)
--	I35605 = NAND(CRC_OUT_1_24, I35603)
--	WX11585 = NAND(I35604, I35605)
--	I35610 = NAND(WX10963, CRC_OUT_1_23)
--	I35611 = NAND(WX10963, I35610)
--	I35612 = NAND(CRC_OUT_1_23, I35610)
--	WX11586 = NAND(I35611, I35612)
--	I35617 = NAND(WX10964, CRC_OUT_1_22)
--	I35618 = NAND(WX10964, I35617)
--	I35619 = NAND(CRC_OUT_1_22, I35617)
--	WX11587 = NAND(I35618, I35619)
--	I35624 = NAND(WX10965, CRC_OUT_1_21)
--	I35625 = NAND(WX10965, I35624)
--	I35626 = NAND(CRC_OUT_1_21, I35624)
--	WX11588 = NAND(I35625, I35626)
--	I35631 = NAND(WX10966, CRC_OUT_1_20)
--	I35632 = NAND(WX10966, I35631)
--	I35633 = NAND(CRC_OUT_1_20, I35631)
--	WX11589 = NAND(I35632, I35633)
--	I35638 = NAND(WX10967, CRC_OUT_1_19)
--	I35639 = NAND(WX10967, I35638)
--	I35640 = NAND(CRC_OUT_1_19, I35638)
--	WX11590 = NAND(I35639, I35640)
--	I35645 = NAND(WX10968, CRC_OUT_1_18)
--	I35646 = NAND(WX10968, I35645)
--	I35647 = NAND(CRC_OUT_1_18, I35645)
--	WX11591 = NAND(I35646, I35647)
--	I35652 = NAND(WX10969, CRC_OUT_1_17)
--	I35653 = NAND(WX10969, I35652)
--	I35654 = NAND(CRC_OUT_1_17, I35652)
--	WX11592 = NAND(I35653, I35654)
--	I35659 = NAND(WX10970, CRC_OUT_1_16)
--	I35660 = NAND(WX10970, I35659)
--	I35661 = NAND(CRC_OUT_1_16, I35659)
--	WX11593 = NAND(I35660, I35661)
--	I35666 = NAND(WX10972, CRC_OUT_1_14)
--	I35667 = NAND(WX10972, I35666)
--	I35668 = NAND(CRC_OUT_1_14, I35666)
--	WX11594 = NAND(I35667, I35668)
--	I35673 = NAND(WX10973, CRC_OUT_1_13)
--	I35674 = NAND(WX10973, I35673)
--	I35675 = NAND(CRC_OUT_1_13, I35673)
--	WX11595 = NAND(I35674, I35675)
--	I35680 = NAND(WX10974, CRC_OUT_1_12)
--	I35681 = NAND(WX10974, I35680)
--	I35682 = NAND(CRC_OUT_1_12, I35680)
--	WX11596 = NAND(I35681, I35682)
--	I35687 = NAND(WX10975, CRC_OUT_1_11)
--	I35688 = NAND(WX10975, I35687)
--	I35689 = NAND(CRC_OUT_1_11, I35687)
--	WX11597 = NAND(I35688, I35689)
--	I35694 = NAND(WX10977, CRC_OUT_1_9)
--	I35695 = NAND(WX10977, I35694)
--	I35696 = NAND(CRC_OUT_1_9, I35694)
--	WX11598 = NAND(I35695, I35696)
--	I35701 = NAND(WX10978, CRC_OUT_1_8)
--	I35702 = NAND(WX10978, I35701)
--	I35703 = NAND(CRC_OUT_1_8, I35701)
--	WX11599 = NAND(I35702, I35703)
--	I35708 = NAND(WX10979, CRC_OUT_1_7)
--	I35709 = NAND(WX10979, I35708)
--	I35710 = NAND(CRC_OUT_1_7, I35708)
--	WX11600 = NAND(I35709, I35710)
--	I35715 = NAND(WX10980, CRC_OUT_1_6)
--	I35716 = NAND(WX10980, I35715)
--	I35717 = NAND(CRC_OUT_1_6, I35715)
--	WX11601 = NAND(I35716, I35717)
--	I35722 = NAND(WX10981, CRC_OUT_1_5)
--	I35723 = NAND(WX10981, I35722)
--	I35724 = NAND(CRC_OUT_1_5, I35722)
--	WX11602 = NAND(I35723, I35724)
--	I35729 = NAND(WX10982, CRC_OUT_1_4)
--	I35730 = NAND(WX10982, I35729)
--	I35731 = NAND(CRC_OUT_1_4, I35729)
--	WX11603 = NAND(I35730, I35731)
--	I35736 = NAND(WX10984, CRC_OUT_1_2)
--	I35737 = NAND(WX10984, I35736)
--	I35738 = NAND(CRC_OUT_1_2, I35736)
--	WX11604 = NAND(I35737, I35738)
--	I35743 = NAND(WX10985, CRC_OUT_1_1)
--	I35744 = NAND(WX10985, I35743)
--	I35745 = NAND(CRC_OUT_1_1, I35743)
--	WX11605 = NAND(I35744, I35745)
--	I35750 = NAND(WX10986, CRC_OUT_1_0)
--	I35751 = NAND(WX10986, I35750)
--	I35752 = NAND(CRC_OUT_1_0, I35750)
--	WX11606 = NAND(I35751, I35752)
--
-- VHDL Output
-- =============
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.MATH_REAL.ALL;

entity s35932 is
	port (
		CLK: in std_logic;
		DATA_0_0: in std_logic;
		DATA_0_1: in std_logic;
		DATA_0_2: in std_logic;
		DATA_0_3: in std_logic;
		DATA_0_4: in std_logic;
		DATA_0_5: in std_logic;
		DATA_0_6: in std_logic;
		DATA_0_7: in std_logic;
		DATA_0_8: in std_logic;
		DATA_0_9: in std_logic;
		DATA_0_10: in std_logic;
		DATA_0_11: in std_logic;
		DATA_0_12: in std_logic;
		DATA_0_13: in std_logic;
		DATA_0_14: in std_logic;
		DATA_0_15: in std_logic;
		DATA_0_16: in std_logic;
		DATA_0_17: in std_logic;
		DATA_0_18: in std_logic;
		DATA_0_19: in std_logic;
		DATA_0_20: in std_logic;
		DATA_0_21: in std_logic;
		DATA_0_22: in std_logic;
		DATA_0_23: in std_logic;
		DATA_0_24: in std_logic;
		DATA_0_25: in std_logic;
		DATA_0_26: in std_logic;
		DATA_0_27: in std_logic;
		DATA_0_28: in std_logic;
		DATA_0_29: in std_logic;
		DATA_0_30: in std_logic;
		DATA_0_31: in std_logic;
		RESET: in std_logic;
		TM0: in std_logic;
		TM1: in std_logic;
		CRC_OUT_1_0: out std_logic;
		CRC_OUT_1_1: out std_logic;
		CRC_OUT_1_2: out std_logic;
		CRC_OUT_1_3: out std_logic;
		CRC_OUT_1_4: out std_logic;
		CRC_OUT_1_5: out std_logic;
		CRC_OUT_1_6: out std_logic;
		CRC_OUT_1_7: out std_logic;
		CRC_OUT_1_8: out std_logic;
		CRC_OUT_1_9: out std_logic;
		CRC_OUT_1_10: out std_logic;
		CRC_OUT_1_11: out std_logic;
		CRC_OUT_1_12: out std_logic;
		CRC_OUT_1_13: out std_logic;
		CRC_OUT_1_14: out std_logic;
		CRC_OUT_1_15: out std_logic;
		CRC_OUT_1_16: out std_logic;
		CRC_OUT_1_17: out std_logic;
		CRC_OUT_1_18: out std_logic;
		CRC_OUT_1_19: out std_logic;
		CRC_OUT_1_20: out std_logic;
		CRC_OUT_1_21: out std_logic;
		CRC_OUT_1_22: out std_logic;
		CRC_OUT_1_23: out std_logic;
		CRC_OUT_1_24: out std_logic;
		CRC_OUT_1_25: out std_logic;
		CRC_OUT_1_26: out std_logic;
		CRC_OUT_1_27: out std_logic;
		CRC_OUT_1_28: out std_logic;
		CRC_OUT_1_29: out std_logic;
		CRC_OUT_1_30: out std_logic;
		CRC_OUT_1_31: out std_logic;
		CRC_OUT_2_0: out std_logic;
		CRC_OUT_2_1: out std_logic;
		CRC_OUT_2_2: out std_logic;
		CRC_OUT_2_3: out std_logic;
		CRC_OUT_2_4: out std_logic;
		CRC_OUT_2_5: out std_logic;
		CRC_OUT_2_6: out std_logic;
		CRC_OUT_2_7: out std_logic;
		CRC_OUT_2_8: out std_logic;
		CRC_OUT_2_9: out std_logic;
		CRC_OUT_2_10: out std_logic;
		CRC_OUT_2_11: out std_logic;
		CRC_OUT_2_12: out std_logic;
		CRC_OUT_2_13: out std_logic;
		CRC_OUT_2_14: out std_logic;
		CRC_OUT_2_15: out std_logic;
		CRC_OUT_2_16: out std_logic;
		CRC_OUT_2_17: out std_logic;
		CRC_OUT_2_18: out std_logic;
		CRC_OUT_2_19: out std_logic;
		CRC_OUT_2_20: out std_logic;
		CRC_OUT_2_21: out std_logic;
		CRC_OUT_2_22: out std_logic;
		CRC_OUT_2_23: out std_logic;
		CRC_OUT_2_24: out std_logic;
		CRC_OUT_2_25: out std_logic;
		CRC_OUT_2_26: out std_logic;
		CRC_OUT_2_27: out std_logic;
		CRC_OUT_2_28: out std_logic;
		CRC_OUT_2_29: out std_logic;
		CRC_OUT_2_30: out std_logic;
		CRC_OUT_2_31: out std_logic;
		CRC_OUT_3_0: out std_logic;
		CRC_OUT_3_1: out std_logic;
		CRC_OUT_3_2: out std_logic;
		CRC_OUT_3_3: out std_logic;
		CRC_OUT_3_4: out std_logic;
		CRC_OUT_3_5: out std_logic;
		CRC_OUT_3_6: out std_logic;
		CRC_OUT_3_7: out std_logic;
		CRC_OUT_3_8: out std_logic;
		CRC_OUT_3_9: out std_logic;
		CRC_OUT_3_10: out std_logic;
		CRC_OUT_3_11: out std_logic;
		CRC_OUT_3_12: out std_logic;
		CRC_OUT_3_13: out std_logic;
		CRC_OUT_3_14: out std_logic;
		CRC_OUT_3_15: out std_logic;
		CRC_OUT_3_16: out std_logic;
		CRC_OUT_3_17: out std_logic;
		CRC_OUT_3_18: out std_logic;
		CRC_OUT_3_19: out std_logic;
		CRC_OUT_3_20: out std_logic;
		CRC_OUT_3_21: out std_logic;
		CRC_OUT_3_22: out std_logic;
		CRC_OUT_3_23: out std_logic;
		CRC_OUT_3_24: out std_logic;
		CRC_OUT_3_25: out std_logic;
		CRC_OUT_3_26: out std_logic;
		CRC_OUT_3_27: out std_logic;
		CRC_OUT_3_28: out std_logic;
		CRC_OUT_3_29: out std_logic;
		CRC_OUT_3_30: out std_logic;
		CRC_OUT_3_31: out std_logic;
		CRC_OUT_4_0: out std_logic;
		CRC_OUT_4_1: out std_logic;
		CRC_OUT_4_2: out std_logic;
		CRC_OUT_4_3: out std_logic;
		CRC_OUT_4_4: out std_logic;
		CRC_OUT_4_5: out std_logic;
		CRC_OUT_4_6: out std_logic;
		CRC_OUT_4_7: out std_logic;
		CRC_OUT_4_8: out std_logic;
		CRC_OUT_4_9: out std_logic;
		CRC_OUT_4_10: out std_logic;
		CRC_OUT_4_11: out std_logic;
		CRC_OUT_4_12: out std_logic;
		CRC_OUT_4_13: out std_logic;
		CRC_OUT_4_14: out std_logic;
		CRC_OUT_4_15: out std_logic;
		CRC_OUT_4_16: out std_logic;
		CRC_OUT_4_17: out std_logic;
		CRC_OUT_4_18: out std_logic;
		CRC_OUT_4_19: out std_logic;
		CRC_OUT_4_20: out std_logic;
		CRC_OUT_4_21: out std_logic;
		CRC_OUT_4_22: out std_logic;
		CRC_OUT_4_23: out std_logic;
		CRC_OUT_4_24: out std_logic;
		CRC_OUT_4_25: out std_logic;
		CRC_OUT_4_26: out std_logic;
		CRC_OUT_4_27: out std_logic;
		CRC_OUT_4_28: out std_logic;
		CRC_OUT_4_29: out std_logic;
		CRC_OUT_4_30: out std_logic;
		CRC_OUT_4_31: out std_logic;
		CRC_OUT_5_0: out std_logic;
		CRC_OUT_5_1: out std_logic;
		CRC_OUT_5_2: out std_logic;
		CRC_OUT_5_3: out std_logic;
		CRC_OUT_5_4: out std_logic;
		CRC_OUT_5_5: out std_logic;
		CRC_OUT_5_6: out std_logic;
		CRC_OUT_5_7: out std_logic;
		CRC_OUT_5_8: out std_logic;
		CRC_OUT_5_9: out std_logic;
		CRC_OUT_5_10: out std_logic;
		CRC_OUT_5_11: out std_logic;
		CRC_OUT_5_12: out std_logic;
		CRC_OUT_5_13: out std_logic;
		CRC_OUT_5_14: out std_logic;
		CRC_OUT_5_15: out std_logic;
		CRC_OUT_5_16: out std_logic;
		CRC_OUT_5_17: out std_logic;
		CRC_OUT_5_18: out std_logic;
		CRC_OUT_5_19: out std_logic;
		CRC_OUT_5_20: out std_logic;
		CRC_OUT_5_21: out std_logic;
		CRC_OUT_5_22: out std_logic;
		CRC_OUT_5_23: out std_logic;
		CRC_OUT_5_24: out std_logic;
		CRC_OUT_5_25: out std_logic;
		CRC_OUT_5_26: out std_logic;
		CRC_OUT_5_27: out std_logic;
		CRC_OUT_5_28: out std_logic;
		CRC_OUT_5_29: out std_logic;
		CRC_OUT_5_30: out std_logic;
		CRC_OUT_5_31: out std_logic;
		CRC_OUT_6_0: out std_logic;
		CRC_OUT_6_1: out std_logic;
		CRC_OUT_6_2: out std_logic;
		CRC_OUT_6_3: out std_logic;
		CRC_OUT_6_4: out std_logic;
		CRC_OUT_6_5: out std_logic;
		CRC_OUT_6_6: out std_logic;
		CRC_OUT_6_7: out std_logic;
		CRC_OUT_6_8: out std_logic;
		CRC_OUT_6_9: out std_logic;
		CRC_OUT_6_10: out std_logic;
		CRC_OUT_6_11: out std_logic;
		CRC_OUT_6_12: out std_logic;
		CRC_OUT_6_13: out std_logic;
		CRC_OUT_6_14: out std_logic;
		CRC_OUT_6_15: out std_logic;
		CRC_OUT_6_16: out std_logic;
		CRC_OUT_6_17: out std_logic;
		CRC_OUT_6_18: out std_logic;
		CRC_OUT_6_19: out std_logic;
		CRC_OUT_6_20: out std_logic;
		CRC_OUT_6_21: out std_logic;
		CRC_OUT_6_22: out std_logic;
		CRC_OUT_6_23: out std_logic;
		CRC_OUT_6_24: out std_logic;
		CRC_OUT_6_25: out std_logic;
		CRC_OUT_6_26: out std_logic;
		CRC_OUT_6_27: out std_logic;
		CRC_OUT_6_28: out std_logic;
		CRC_OUT_6_29: out std_logic;
		CRC_OUT_6_30: out std_logic;
		CRC_OUT_6_31: out std_logic;
		CRC_OUT_7_0: out std_logic;
		CRC_OUT_7_1: out std_logic;
		CRC_OUT_7_2: out std_logic;
		CRC_OUT_7_3: out std_logic;
		CRC_OUT_7_4: out std_logic;
		CRC_OUT_7_5: out std_logic;
		CRC_OUT_7_6: out std_logic;
		CRC_OUT_7_7: out std_logic;
		CRC_OUT_7_8: out std_logic;
		CRC_OUT_7_9: out std_logic;
		CRC_OUT_7_10: out std_logic;
		CRC_OUT_7_11: out std_logic;
		CRC_OUT_7_12: out std_logic;
		CRC_OUT_7_13: out std_logic;
		CRC_OUT_7_14: out std_logic;
		CRC_OUT_7_15: out std_logic;
		CRC_OUT_7_16: out std_logic;
		CRC_OUT_7_17: out std_logic;
		CRC_OUT_7_18: out std_logic;
		CRC_OUT_7_19: out std_logic;
		CRC_OUT_7_20: out std_logic;
		CRC_OUT_7_21: out std_logic;
		CRC_OUT_7_22: out std_logic;
		CRC_OUT_7_23: out std_logic;
		CRC_OUT_7_24: out std_logic;
		CRC_OUT_7_25: out std_logic;
		CRC_OUT_7_26: out std_logic;
		CRC_OUT_7_27: out std_logic;
		CRC_OUT_7_28: out std_logic;
		CRC_OUT_7_29: out std_logic;
		CRC_OUT_7_30: out std_logic;
		CRC_OUT_7_31: out std_logic;
		CRC_OUT_8_0: out std_logic;
		CRC_OUT_8_1: out std_logic;
		CRC_OUT_8_2: out std_logic;
		CRC_OUT_8_3: out std_logic;
		CRC_OUT_8_4: out std_logic;
		CRC_OUT_8_5: out std_logic;
		CRC_OUT_8_6: out std_logic;
		CRC_OUT_8_7: out std_logic;
		CRC_OUT_8_8: out std_logic;
		CRC_OUT_8_9: out std_logic;
		CRC_OUT_8_10: out std_logic;
		CRC_OUT_8_11: out std_logic;
		CRC_OUT_8_12: out std_logic;
		CRC_OUT_8_13: out std_logic;
		CRC_OUT_8_14: out std_logic;
		CRC_OUT_8_15: out std_logic;
		CRC_OUT_8_16: out std_logic;
		CRC_OUT_8_17: out std_logic;
		CRC_OUT_8_18: out std_logic;
		CRC_OUT_8_19: out std_logic;
		CRC_OUT_8_20: out std_logic;
		CRC_OUT_8_21: out std_logic;
		CRC_OUT_8_22: out std_logic;
		CRC_OUT_8_23: out std_logic;
		CRC_OUT_8_24: out std_logic;
		CRC_OUT_8_25: out std_logic;
		CRC_OUT_8_26: out std_logic;
		CRC_OUT_8_27: out std_logic;
		CRC_OUT_8_28: out std_logic;
		CRC_OUT_8_29: out std_logic;
		CRC_OUT_8_30: out std_logic;
		CRC_OUT_8_31: out std_logic;
		CRC_OUT_9_0: out std_logic;
		CRC_OUT_9_1: out std_logic;
		CRC_OUT_9_2: out std_logic;
		CRC_OUT_9_3: out std_logic;
		CRC_OUT_9_4: out std_logic;
		CRC_OUT_9_5: out std_logic;
		CRC_OUT_9_6: out std_logic;
		CRC_OUT_9_7: out std_logic;
		CRC_OUT_9_8: out std_logic;
		CRC_OUT_9_9: out std_logic;
		CRC_OUT_9_10: out std_logic;
		CRC_OUT_9_11: out std_logic;
		CRC_OUT_9_12: out std_logic;
		CRC_OUT_9_13: out std_logic;
		CRC_OUT_9_14: out std_logic;
		CRC_OUT_9_15: out std_logic;
		CRC_OUT_9_16: out std_logic;
		CRC_OUT_9_17: out std_logic;
		CRC_OUT_9_18: out std_logic;
		CRC_OUT_9_19: out std_logic;
		CRC_OUT_9_20: out std_logic;
		CRC_OUT_9_21: out std_logic;
		CRC_OUT_9_22: out std_logic;
		CRC_OUT_9_23: out std_logic;
		CRC_OUT_9_24: out std_logic;
		CRC_OUT_9_25: out std_logic;
		CRC_OUT_9_26: out std_logic;
		CRC_OUT_9_27: out std_logic;
		CRC_OUT_9_28: out std_logic;
		CRC_OUT_9_29: out std_logic;
		CRC_OUT_9_30: out std_logic;
		CRC_OUT_9_31: out std_logic;
		DATA_9_0: out std_logic;
		DATA_9_1: out std_logic;
		DATA_9_2: out std_logic;
		DATA_9_3: out std_logic;
		DATA_9_4: out std_logic;
		DATA_9_5: out std_logic;
		DATA_9_6: out std_logic;
		DATA_9_7: out std_logic;
		DATA_9_8: out std_logic;
		DATA_9_9: out std_logic;
		DATA_9_10: out std_logic;
		DATA_9_11: out std_logic;
		DATA_9_12: out std_logic;
		DATA_9_13: out std_logic;
		DATA_9_14: out std_logic;
		DATA_9_15: out std_logic;
		DATA_9_16: out std_logic;
		DATA_9_17: out std_logic;
		DATA_9_18: out std_logic;
		DATA_9_19: out std_logic;
		DATA_9_20: out std_logic;
		DATA_9_21: out std_logic;
		DATA_9_22: out std_logic;
		DATA_9_23: out std_logic;
		DATA_9_24: out std_logic;
		DATA_9_25: out std_logic;
		DATA_9_26: out std_logic;
		DATA_9_27: out std_logic;
		DATA_9_28: out std_logic;
		DATA_9_29: out std_logic;
		DATA_9_30: out std_logic;
		DATA_9_31: out std_logic
	);
end entity;

architecture RTL of s35932 is
	attribute dont_touch: boolean;

	signal I1986: std_logic; attribute dont_touch of I1986: signal is true;
	signal I1987: std_logic; attribute dont_touch of I1987: signal is true;
	signal I1988: std_logic; attribute dont_touch of I1988: signal is true;
	signal I1989: std_logic; attribute dont_touch of I1989: signal is true;
	signal I1990: std_logic; attribute dont_touch of I1990: signal is true;
	signal I1995: std_logic; attribute dont_touch of I1995: signal is true;
	signal I1996: std_logic; attribute dont_touch of I1996: signal is true;
	signal I1997: std_logic; attribute dont_touch of I1997: signal is true;
	signal I2002: std_logic; attribute dont_touch of I2002: signal is true;
	signal I2003: std_logic; attribute dont_touch of I2003: signal is true;
	signal I2004: std_logic; attribute dont_touch of I2004: signal is true;
	signal I2005: std_logic; attribute dont_touch of I2005: signal is true;
	signal I2010: std_logic; attribute dont_touch of I2010: signal is true;
	signal I2011: std_logic; attribute dont_touch of I2011: signal is true;
	signal I2012: std_logic; attribute dont_touch of I2012: signal is true;
	signal I2017: std_logic; attribute dont_touch of I2017: signal is true;
	signal I2018: std_logic; attribute dont_touch of I2018: signal is true;
	signal I2019: std_logic; attribute dont_touch of I2019: signal is true;
	signal I2020: std_logic; attribute dont_touch of I2020: signal is true;
	signal I2021: std_logic; attribute dont_touch of I2021: signal is true;
	signal I2026: std_logic; attribute dont_touch of I2026: signal is true;
	signal I2027: std_logic; attribute dont_touch of I2027: signal is true;
	signal I2028: std_logic; attribute dont_touch of I2028: signal is true;
	signal I2033: std_logic; attribute dont_touch of I2033: signal is true;
	signal I2034: std_logic; attribute dont_touch of I2034: signal is true;
	signal I2035: std_logic; attribute dont_touch of I2035: signal is true;
	signal I2036: std_logic; attribute dont_touch of I2036: signal is true;
	signal I2041: std_logic; attribute dont_touch of I2041: signal is true;
	signal I2042: std_logic; attribute dont_touch of I2042: signal is true;
	signal I2043: std_logic; attribute dont_touch of I2043: signal is true;
	signal I2048: std_logic; attribute dont_touch of I2048: signal is true;
	signal I2049: std_logic; attribute dont_touch of I2049: signal is true;
	signal I2050: std_logic; attribute dont_touch of I2050: signal is true;
	signal I2051: std_logic; attribute dont_touch of I2051: signal is true;
	signal I2052: std_logic; attribute dont_touch of I2052: signal is true;
	signal I2057: std_logic; attribute dont_touch of I2057: signal is true;
	signal I2058: std_logic; attribute dont_touch of I2058: signal is true;
	signal I2059: std_logic; attribute dont_touch of I2059: signal is true;
	signal I2064: std_logic; attribute dont_touch of I2064: signal is true;
	signal I2065: std_logic; attribute dont_touch of I2065: signal is true;
	signal I2066: std_logic; attribute dont_touch of I2066: signal is true;
	signal I2067: std_logic; attribute dont_touch of I2067: signal is true;
	signal I2072: std_logic; attribute dont_touch of I2072: signal is true;
	signal I2073: std_logic; attribute dont_touch of I2073: signal is true;
	signal I2074: std_logic; attribute dont_touch of I2074: signal is true;
	signal I2079: std_logic; attribute dont_touch of I2079: signal is true;
	signal I2080: std_logic; attribute dont_touch of I2080: signal is true;
	signal I2081: std_logic; attribute dont_touch of I2081: signal is true;
	signal I2082: std_logic; attribute dont_touch of I2082: signal is true;
	signal I2083: std_logic; attribute dont_touch of I2083: signal is true;
	signal I2088: std_logic; attribute dont_touch of I2088: signal is true;
	signal I2089: std_logic; attribute dont_touch of I2089: signal is true;
	signal I2090: std_logic; attribute dont_touch of I2090: signal is true;
	signal I2095: std_logic; attribute dont_touch of I2095: signal is true;
	signal I2096: std_logic; attribute dont_touch of I2096: signal is true;
	signal I2097: std_logic; attribute dont_touch of I2097: signal is true;
	signal I2098: std_logic; attribute dont_touch of I2098: signal is true;
	signal I2103: std_logic; attribute dont_touch of I2103: signal is true;
	signal I2104: std_logic; attribute dont_touch of I2104: signal is true;
	signal I2105: std_logic; attribute dont_touch of I2105: signal is true;
	signal I2110: std_logic; attribute dont_touch of I2110: signal is true;
	signal I2111: std_logic; attribute dont_touch of I2111: signal is true;
	signal I2112: std_logic; attribute dont_touch of I2112: signal is true;
	signal I2113: std_logic; attribute dont_touch of I2113: signal is true;
	signal I2114: std_logic; attribute dont_touch of I2114: signal is true;
	signal I2119: std_logic; attribute dont_touch of I2119: signal is true;
	signal I2120: std_logic; attribute dont_touch of I2120: signal is true;
	signal I2121: std_logic; attribute dont_touch of I2121: signal is true;
	signal I2126: std_logic; attribute dont_touch of I2126: signal is true;
	signal I2127: std_logic; attribute dont_touch of I2127: signal is true;
	signal I2128: std_logic; attribute dont_touch of I2128: signal is true;
	signal I2129: std_logic; attribute dont_touch of I2129: signal is true;
	signal I2134: std_logic; attribute dont_touch of I2134: signal is true;
	signal I2135: std_logic; attribute dont_touch of I2135: signal is true;
	signal I2136: std_logic; attribute dont_touch of I2136: signal is true;
	signal I2141: std_logic; attribute dont_touch of I2141: signal is true;
	signal I2142: std_logic; attribute dont_touch of I2142: signal is true;
	signal I2143: std_logic; attribute dont_touch of I2143: signal is true;
	signal I2144: std_logic; attribute dont_touch of I2144: signal is true;
	signal I2145: std_logic; attribute dont_touch of I2145: signal is true;
	signal I2150: std_logic; attribute dont_touch of I2150: signal is true;
	signal I2151: std_logic; attribute dont_touch of I2151: signal is true;
	signal I2152: std_logic; attribute dont_touch of I2152: signal is true;
	signal I2157: std_logic; attribute dont_touch of I2157: signal is true;
	signal I2158: std_logic; attribute dont_touch of I2158: signal is true;
	signal I2159: std_logic; attribute dont_touch of I2159: signal is true;
	signal I2160: std_logic; attribute dont_touch of I2160: signal is true;
	signal I2165: std_logic; attribute dont_touch of I2165: signal is true;
	signal I2166: std_logic; attribute dont_touch of I2166: signal is true;
	signal I2167: std_logic; attribute dont_touch of I2167: signal is true;
	signal I2172: std_logic; attribute dont_touch of I2172: signal is true;
	signal I2173: std_logic; attribute dont_touch of I2173: signal is true;
	signal I2174: std_logic; attribute dont_touch of I2174: signal is true;
	signal I2175: std_logic; attribute dont_touch of I2175: signal is true;
	signal I2176: std_logic; attribute dont_touch of I2176: signal is true;
	signal I2181: std_logic; attribute dont_touch of I2181: signal is true;
	signal I2182: std_logic; attribute dont_touch of I2182: signal is true;
	signal I2183: std_logic; attribute dont_touch of I2183: signal is true;
	signal I2188: std_logic; attribute dont_touch of I2188: signal is true;
	signal I2189: std_logic; attribute dont_touch of I2189: signal is true;
	signal I2190: std_logic; attribute dont_touch of I2190: signal is true;
	signal I2191: std_logic; attribute dont_touch of I2191: signal is true;
	signal I2196: std_logic; attribute dont_touch of I2196: signal is true;
	signal I2197: std_logic; attribute dont_touch of I2197: signal is true;
	signal I2198: std_logic; attribute dont_touch of I2198: signal is true;
	signal I2203: std_logic; attribute dont_touch of I2203: signal is true;
	signal I2204: std_logic; attribute dont_touch of I2204: signal is true;
	signal I2205: std_logic; attribute dont_touch of I2205: signal is true;
	signal I2206: std_logic; attribute dont_touch of I2206: signal is true;
	signal I2207: std_logic; attribute dont_touch of I2207: signal is true;
	signal I2212: std_logic; attribute dont_touch of I2212: signal is true;
	signal I2213: std_logic; attribute dont_touch of I2213: signal is true;
	signal I2214: std_logic; attribute dont_touch of I2214: signal is true;
	signal I2219: std_logic; attribute dont_touch of I2219: signal is true;
	signal I2220: std_logic; attribute dont_touch of I2220: signal is true;
	signal I2221: std_logic; attribute dont_touch of I2221: signal is true;
	signal I2222: std_logic; attribute dont_touch of I2222: signal is true;
	signal I2227: std_logic; attribute dont_touch of I2227: signal is true;
	signal I2228: std_logic; attribute dont_touch of I2228: signal is true;
	signal I2229: std_logic; attribute dont_touch of I2229: signal is true;
	signal I2234: std_logic; attribute dont_touch of I2234: signal is true;
	signal I2235: std_logic; attribute dont_touch of I2235: signal is true;
	signal I2236: std_logic; attribute dont_touch of I2236: signal is true;
	signal I2237: std_logic; attribute dont_touch of I2237: signal is true;
	signal I2238: std_logic; attribute dont_touch of I2238: signal is true;
	signal I2243: std_logic; attribute dont_touch of I2243: signal is true;
	signal I2244: std_logic; attribute dont_touch of I2244: signal is true;
	signal I2245: std_logic; attribute dont_touch of I2245: signal is true;
	signal I2250: std_logic; attribute dont_touch of I2250: signal is true;
	signal I2251: std_logic; attribute dont_touch of I2251: signal is true;
	signal I2252: std_logic; attribute dont_touch of I2252: signal is true;
	signal I2253: std_logic; attribute dont_touch of I2253: signal is true;
	signal I2258: std_logic; attribute dont_touch of I2258: signal is true;
	signal I2259: std_logic; attribute dont_touch of I2259: signal is true;
	signal I2260: std_logic; attribute dont_touch of I2260: signal is true;
	signal I2265: std_logic; attribute dont_touch of I2265: signal is true;
	signal I2266: std_logic; attribute dont_touch of I2266: signal is true;
	signal I2267: std_logic; attribute dont_touch of I2267: signal is true;
	signal I2268: std_logic; attribute dont_touch of I2268: signal is true;
	signal I2269: std_logic; attribute dont_touch of I2269: signal is true;
	signal I2274: std_logic; attribute dont_touch of I2274: signal is true;
	signal I2275: std_logic; attribute dont_touch of I2275: signal is true;
	signal I2276: std_logic; attribute dont_touch of I2276: signal is true;
	signal I2281: std_logic; attribute dont_touch of I2281: signal is true;
	signal I2282: std_logic; attribute dont_touch of I2282: signal is true;
	signal I2283: std_logic; attribute dont_touch of I2283: signal is true;
	signal I2284: std_logic; attribute dont_touch of I2284: signal is true;
	signal I2289: std_logic; attribute dont_touch of I2289: signal is true;
	signal I2290: std_logic; attribute dont_touch of I2290: signal is true;
	signal I2291: std_logic; attribute dont_touch of I2291: signal is true;
	signal I2296: std_logic; attribute dont_touch of I2296: signal is true;
	signal I2297: std_logic; attribute dont_touch of I2297: signal is true;
	signal I2298: std_logic; attribute dont_touch of I2298: signal is true;
	signal I2299: std_logic; attribute dont_touch of I2299: signal is true;
	signal I2300: std_logic; attribute dont_touch of I2300: signal is true;
	signal I2305: std_logic; attribute dont_touch of I2305: signal is true;
	signal I2306: std_logic; attribute dont_touch of I2306: signal is true;
	signal I2307: std_logic; attribute dont_touch of I2307: signal is true;
	signal I2312: std_logic; attribute dont_touch of I2312: signal is true;
	signal I2313: std_logic; attribute dont_touch of I2313: signal is true;
	signal I2314: std_logic; attribute dont_touch of I2314: signal is true;
	signal I2315: std_logic; attribute dont_touch of I2315: signal is true;
	signal I2320: std_logic; attribute dont_touch of I2320: signal is true;
	signal I2321: std_logic; attribute dont_touch of I2321: signal is true;
	signal I2322: std_logic; attribute dont_touch of I2322: signal is true;
	signal I2327: std_logic; attribute dont_touch of I2327: signal is true;
	signal I2328: std_logic; attribute dont_touch of I2328: signal is true;
	signal I2329: std_logic; attribute dont_touch of I2329: signal is true;
	signal I2330: std_logic; attribute dont_touch of I2330: signal is true;
	signal I2331: std_logic; attribute dont_touch of I2331: signal is true;
	signal I2336: std_logic; attribute dont_touch of I2336: signal is true;
	signal I2337: std_logic; attribute dont_touch of I2337: signal is true;
	signal I2338: std_logic; attribute dont_touch of I2338: signal is true;
	signal I2343: std_logic; attribute dont_touch of I2343: signal is true;
	signal I2344: std_logic; attribute dont_touch of I2344: signal is true;
	signal I2345: std_logic; attribute dont_touch of I2345: signal is true;
	signal I2346: std_logic; attribute dont_touch of I2346: signal is true;
	signal I2351: std_logic; attribute dont_touch of I2351: signal is true;
	signal I2352: std_logic; attribute dont_touch of I2352: signal is true;
	signal I2353: std_logic; attribute dont_touch of I2353: signal is true;
	signal I2358: std_logic; attribute dont_touch of I2358: signal is true;
	signal I2359: std_logic; attribute dont_touch of I2359: signal is true;
	signal I2360: std_logic; attribute dont_touch of I2360: signal is true;
	signal I2361: std_logic; attribute dont_touch of I2361: signal is true;
	signal I2362: std_logic; attribute dont_touch of I2362: signal is true;
	signal I2367: std_logic; attribute dont_touch of I2367: signal is true;
	signal I2368: std_logic; attribute dont_touch of I2368: signal is true;
	signal I2369: std_logic; attribute dont_touch of I2369: signal is true;
	signal I2374: std_logic; attribute dont_touch of I2374: signal is true;
	signal I2375: std_logic; attribute dont_touch of I2375: signal is true;
	signal I2376: std_logic; attribute dont_touch of I2376: signal is true;
	signal I2377: std_logic; attribute dont_touch of I2377: signal is true;
	signal I2382: std_logic; attribute dont_touch of I2382: signal is true;
	signal I2383: std_logic; attribute dont_touch of I2383: signal is true;
	signal I2384: std_logic; attribute dont_touch of I2384: signal is true;
	signal I2389: std_logic; attribute dont_touch of I2389: signal is true;
	signal I2390: std_logic; attribute dont_touch of I2390: signal is true;
	signal I2391: std_logic; attribute dont_touch of I2391: signal is true;
	signal I2392: std_logic; attribute dont_touch of I2392: signal is true;
	signal I2393: std_logic; attribute dont_touch of I2393: signal is true;
	signal I2398: std_logic; attribute dont_touch of I2398: signal is true;
	signal I2399: std_logic; attribute dont_touch of I2399: signal is true;
	signal I2400: std_logic; attribute dont_touch of I2400: signal is true;
	signal I2405: std_logic; attribute dont_touch of I2405: signal is true;
	signal I2406: std_logic; attribute dont_touch of I2406: signal is true;
	signal I2407: std_logic; attribute dont_touch of I2407: signal is true;
	signal I2408: std_logic; attribute dont_touch of I2408: signal is true;
	signal I2413: std_logic; attribute dont_touch of I2413: signal is true;
	signal I2414: std_logic; attribute dont_touch of I2414: signal is true;
	signal I2415: std_logic; attribute dont_touch of I2415: signal is true;
	signal I2420: std_logic; attribute dont_touch of I2420: signal is true;
	signal I2421: std_logic; attribute dont_touch of I2421: signal is true;
	signal I2422: std_logic; attribute dont_touch of I2422: signal is true;
	signal I2423: std_logic; attribute dont_touch of I2423: signal is true;
	signal I2424: std_logic; attribute dont_touch of I2424: signal is true;
	signal I2429: std_logic; attribute dont_touch of I2429: signal is true;
	signal I2430: std_logic; attribute dont_touch of I2430: signal is true;
	signal I2431: std_logic; attribute dont_touch of I2431: signal is true;
	signal I2436: std_logic; attribute dont_touch of I2436: signal is true;
	signal I2437: std_logic; attribute dont_touch of I2437: signal is true;
	signal I2438: std_logic; attribute dont_touch of I2438: signal is true;
	signal I2439: std_logic; attribute dont_touch of I2439: signal is true;
	signal I2444: std_logic; attribute dont_touch of I2444: signal is true;
	signal I2445: std_logic; attribute dont_touch of I2445: signal is true;
	signal I2446: std_logic; attribute dont_touch of I2446: signal is true;
	signal I2451: std_logic; attribute dont_touch of I2451: signal is true;
	signal I2452: std_logic; attribute dont_touch of I2452: signal is true;
	signal I2453: std_logic; attribute dont_touch of I2453: signal is true;
	signal I2454: std_logic; attribute dont_touch of I2454: signal is true;
	signal I2455: std_logic; attribute dont_touch of I2455: signal is true;
	signal I2460: std_logic; attribute dont_touch of I2460: signal is true;
	signal I2461: std_logic; attribute dont_touch of I2461: signal is true;
	signal I2462: std_logic; attribute dont_touch of I2462: signal is true;
	signal I2467: std_logic; attribute dont_touch of I2467: signal is true;
	signal I2468: std_logic; attribute dont_touch of I2468: signal is true;
	signal I2469: std_logic; attribute dont_touch of I2469: signal is true;
	signal I2470: std_logic; attribute dont_touch of I2470: signal is true;
	signal I2475: std_logic; attribute dont_touch of I2475: signal is true;
	signal I2476: std_logic; attribute dont_touch of I2476: signal is true;
	signal I2477: std_logic; attribute dont_touch of I2477: signal is true;
	signal I2482: std_logic; attribute dont_touch of I2482: signal is true;
	signal I2483: std_logic; attribute dont_touch of I2483: signal is true;
	signal I2484: std_logic; attribute dont_touch of I2484: signal is true;
	signal I2485: std_logic; attribute dont_touch of I2485: signal is true;
	signal I2486: std_logic; attribute dont_touch of I2486: signal is true;
	signal I2491: std_logic; attribute dont_touch of I2491: signal is true;
	signal I2492: std_logic; attribute dont_touch of I2492: signal is true;
	signal I2493: std_logic; attribute dont_touch of I2493: signal is true;
	signal I2498: std_logic; attribute dont_touch of I2498: signal is true;
	signal I2499: std_logic; attribute dont_touch of I2499: signal is true;
	signal I2500: std_logic; attribute dont_touch of I2500: signal is true;
	signal I2501: std_logic; attribute dont_touch of I2501: signal is true;
	signal I2506: std_logic; attribute dont_touch of I2506: signal is true;
	signal I2507: std_logic; attribute dont_touch of I2507: signal is true;
	signal I2508: std_logic; attribute dont_touch of I2508: signal is true;
	signal I2513: std_logic; attribute dont_touch of I2513: signal is true;
	signal I2514: std_logic; attribute dont_touch of I2514: signal is true;
	signal I2515: std_logic; attribute dont_touch of I2515: signal is true;
	signal I2516: std_logic; attribute dont_touch of I2516: signal is true;
	signal I2517: std_logic; attribute dont_touch of I2517: signal is true;
	signal I2522: std_logic; attribute dont_touch of I2522: signal is true;
	signal I2523: std_logic; attribute dont_touch of I2523: signal is true;
	signal I2524: std_logic; attribute dont_touch of I2524: signal is true;
	signal I2529: std_logic; attribute dont_touch of I2529: signal is true;
	signal I2530: std_logic; attribute dont_touch of I2530: signal is true;
	signal I2531: std_logic; attribute dont_touch of I2531: signal is true;
	signal I2532: std_logic; attribute dont_touch of I2532: signal is true;
	signal I2537: std_logic; attribute dont_touch of I2537: signal is true;
	signal I2538: std_logic; attribute dont_touch of I2538: signal is true;
	signal I2539: std_logic; attribute dont_touch of I2539: signal is true;
	signal I2544: std_logic; attribute dont_touch of I2544: signal is true;
	signal I2545: std_logic; attribute dont_touch of I2545: signal is true;
	signal I2546: std_logic; attribute dont_touch of I2546: signal is true;
	signal I2547: std_logic; attribute dont_touch of I2547: signal is true;
	signal I2548: std_logic; attribute dont_touch of I2548: signal is true;
	signal I2553: std_logic; attribute dont_touch of I2553: signal is true;
	signal I2554: std_logic; attribute dont_touch of I2554: signal is true;
	signal I2555: std_logic; attribute dont_touch of I2555: signal is true;
	signal I2560: std_logic; attribute dont_touch of I2560: signal is true;
	signal I2561: std_logic; attribute dont_touch of I2561: signal is true;
	signal I2562: std_logic; attribute dont_touch of I2562: signal is true;
	signal I2563: std_logic; attribute dont_touch of I2563: signal is true;
	signal I2568: std_logic; attribute dont_touch of I2568: signal is true;
	signal I2569: std_logic; attribute dont_touch of I2569: signal is true;
	signal I2570: std_logic; attribute dont_touch of I2570: signal is true;
	signal I2575: std_logic; attribute dont_touch of I2575: signal is true;
	signal I2576: std_logic; attribute dont_touch of I2576: signal is true;
	signal I2577: std_logic; attribute dont_touch of I2577: signal is true;
	signal I2578: std_logic; attribute dont_touch of I2578: signal is true;
	signal I2579: std_logic; attribute dont_touch of I2579: signal is true;
	signal I2584: std_logic; attribute dont_touch of I2584: signal is true;
	signal I2585: std_logic; attribute dont_touch of I2585: signal is true;
	signal I2586: std_logic; attribute dont_touch of I2586: signal is true;
	signal I2591: std_logic; attribute dont_touch of I2591: signal is true;
	signal I2592: std_logic; attribute dont_touch of I2592: signal is true;
	signal I2593: std_logic; attribute dont_touch of I2593: signal is true;
	signal I2594: std_logic; attribute dont_touch of I2594: signal is true;
	signal I2599: std_logic; attribute dont_touch of I2599: signal is true;
	signal I2600: std_logic; attribute dont_touch of I2600: signal is true;
	signal I2601: std_logic; attribute dont_touch of I2601: signal is true;
	signal I2606: std_logic; attribute dont_touch of I2606: signal is true;
	signal I2607: std_logic; attribute dont_touch of I2607: signal is true;
	signal I2608: std_logic; attribute dont_touch of I2608: signal is true;
	signal I2609: std_logic; attribute dont_touch of I2609: signal is true;
	signal I2610: std_logic; attribute dont_touch of I2610: signal is true;
	signal I2615: std_logic; attribute dont_touch of I2615: signal is true;
	signal I2616: std_logic; attribute dont_touch of I2616: signal is true;
	signal I2617: std_logic; attribute dont_touch of I2617: signal is true;
	signal I2622: std_logic; attribute dont_touch of I2622: signal is true;
	signal I2623: std_logic; attribute dont_touch of I2623: signal is true;
	signal I2624: std_logic; attribute dont_touch of I2624: signal is true;
	signal I2625: std_logic; attribute dont_touch of I2625: signal is true;
	signal I2630: std_logic; attribute dont_touch of I2630: signal is true;
	signal I2631: std_logic; attribute dont_touch of I2631: signal is true;
	signal I2632: std_logic; attribute dont_touch of I2632: signal is true;
	signal I2637: std_logic; attribute dont_touch of I2637: signal is true;
	signal I2638: std_logic; attribute dont_touch of I2638: signal is true;
	signal I2639: std_logic; attribute dont_touch of I2639: signal is true;
	signal I2640: std_logic; attribute dont_touch of I2640: signal is true;
	signal I2641: std_logic; attribute dont_touch of I2641: signal is true;
	signal I2646: std_logic; attribute dont_touch of I2646: signal is true;
	signal I2647: std_logic; attribute dont_touch of I2647: signal is true;
	signal I2648: std_logic; attribute dont_touch of I2648: signal is true;
	signal I2653: std_logic; attribute dont_touch of I2653: signal is true;
	signal I2654: std_logic; attribute dont_touch of I2654: signal is true;
	signal I2655: std_logic; attribute dont_touch of I2655: signal is true;
	signal I2656: std_logic; attribute dont_touch of I2656: signal is true;
	signal I2661: std_logic; attribute dont_touch of I2661: signal is true;
	signal I2662: std_logic; attribute dont_touch of I2662: signal is true;
	signal I2663: std_logic; attribute dont_touch of I2663: signal is true;
	signal I2668: std_logic; attribute dont_touch of I2668: signal is true;
	signal I2669: std_logic; attribute dont_touch of I2669: signal is true;
	signal I2670: std_logic; attribute dont_touch of I2670: signal is true;
	signal I2671: std_logic; attribute dont_touch of I2671: signal is true;
	signal I2672: std_logic; attribute dont_touch of I2672: signal is true;
	signal I2677: std_logic; attribute dont_touch of I2677: signal is true;
	signal I2678: std_logic; attribute dont_touch of I2678: signal is true;
	signal I2679: std_logic; attribute dont_touch of I2679: signal is true;
	signal I2684: std_logic; attribute dont_touch of I2684: signal is true;
	signal I2685: std_logic; attribute dont_touch of I2685: signal is true;
	signal I2686: std_logic; attribute dont_touch of I2686: signal is true;
	signal I2687: std_logic; attribute dont_touch of I2687: signal is true;
	signal I2692: std_logic; attribute dont_touch of I2692: signal is true;
	signal I2693: std_logic; attribute dont_touch of I2693: signal is true;
	signal I2694: std_logic; attribute dont_touch of I2694: signal is true;
	signal I2699: std_logic; attribute dont_touch of I2699: signal is true;
	signal I2700: std_logic; attribute dont_touch of I2700: signal is true;
	signal I2701: std_logic; attribute dont_touch of I2701: signal is true;
	signal I2702: std_logic; attribute dont_touch of I2702: signal is true;
	signal I2703: std_logic; attribute dont_touch of I2703: signal is true;
	signal I2708: std_logic; attribute dont_touch of I2708: signal is true;
	signal I2709: std_logic; attribute dont_touch of I2709: signal is true;
	signal I2710: std_logic; attribute dont_touch of I2710: signal is true;
	signal I2715: std_logic; attribute dont_touch of I2715: signal is true;
	signal I2716: std_logic; attribute dont_touch of I2716: signal is true;
	signal I2717: std_logic; attribute dont_touch of I2717: signal is true;
	signal I2718: std_logic; attribute dont_touch of I2718: signal is true;
	signal I2723: std_logic; attribute dont_touch of I2723: signal is true;
	signal I2724: std_logic; attribute dont_touch of I2724: signal is true;
	signal I2725: std_logic; attribute dont_touch of I2725: signal is true;
	signal I2730: std_logic; attribute dont_touch of I2730: signal is true;
	signal I2731: std_logic; attribute dont_touch of I2731: signal is true;
	signal I2732: std_logic; attribute dont_touch of I2732: signal is true;
	signal I2733: std_logic; attribute dont_touch of I2733: signal is true;
	signal I2734: std_logic; attribute dont_touch of I2734: signal is true;
	signal I2739: std_logic; attribute dont_touch of I2739: signal is true;
	signal I2740: std_logic; attribute dont_touch of I2740: signal is true;
	signal I2741: std_logic; attribute dont_touch of I2741: signal is true;
	signal I2746: std_logic; attribute dont_touch of I2746: signal is true;
	signal I2747: std_logic; attribute dont_touch of I2747: signal is true;
	signal I2748: std_logic; attribute dont_touch of I2748: signal is true;
	signal I2749: std_logic; attribute dont_touch of I2749: signal is true;
	signal I2754: std_logic; attribute dont_touch of I2754: signal is true;
	signal I2755: std_logic; attribute dont_touch of I2755: signal is true;
	signal I2756: std_logic; attribute dont_touch of I2756: signal is true;
	signal I2761: std_logic; attribute dont_touch of I2761: signal is true;
	signal I2762: std_logic; attribute dont_touch of I2762: signal is true;
	signal I2763: std_logic; attribute dont_touch of I2763: signal is true;
	signal I2764: std_logic; attribute dont_touch of I2764: signal is true;
	signal I2765: std_logic; attribute dont_touch of I2765: signal is true;
	signal I2770: std_logic; attribute dont_touch of I2770: signal is true;
	signal I2771: std_logic; attribute dont_touch of I2771: signal is true;
	signal I2772: std_logic; attribute dont_touch of I2772: signal is true;
	signal I2777: std_logic; attribute dont_touch of I2777: signal is true;
	signal I2778: std_logic; attribute dont_touch of I2778: signal is true;
	signal I2779: std_logic; attribute dont_touch of I2779: signal is true;
	signal I2780: std_logic; attribute dont_touch of I2780: signal is true;
	signal I2785: std_logic; attribute dont_touch of I2785: signal is true;
	signal I2786: std_logic; attribute dont_touch of I2786: signal is true;
	signal I2787: std_logic; attribute dont_touch of I2787: signal is true;
	signal I2792: std_logic; attribute dont_touch of I2792: signal is true;
	signal I2793: std_logic; attribute dont_touch of I2793: signal is true;
	signal I2794: std_logic; attribute dont_touch of I2794: signal is true;
	signal I2795: std_logic; attribute dont_touch of I2795: signal is true;
	signal I2796: std_logic; attribute dont_touch of I2796: signal is true;
	signal I2801: std_logic; attribute dont_touch of I2801: signal is true;
	signal I2802: std_logic; attribute dont_touch of I2802: signal is true;
	signal I2803: std_logic; attribute dont_touch of I2803: signal is true;
	signal I2808: std_logic; attribute dont_touch of I2808: signal is true;
	signal I2809: std_logic; attribute dont_touch of I2809: signal is true;
	signal I2810: std_logic; attribute dont_touch of I2810: signal is true;
	signal I2811: std_logic; attribute dont_touch of I2811: signal is true;
	signal I2816: std_logic; attribute dont_touch of I2816: signal is true;
	signal I2817: std_logic; attribute dont_touch of I2817: signal is true;
	signal I2818: std_logic; attribute dont_touch of I2818: signal is true;
	signal I2823: std_logic; attribute dont_touch of I2823: signal is true;
	signal I2824: std_logic; attribute dont_touch of I2824: signal is true;
	signal I2825: std_logic; attribute dont_touch of I2825: signal is true;
	signal I2826: std_logic; attribute dont_touch of I2826: signal is true;
	signal I2827: std_logic; attribute dont_touch of I2827: signal is true;
	signal I2832: std_logic; attribute dont_touch of I2832: signal is true;
	signal I2833: std_logic; attribute dont_touch of I2833: signal is true;
	signal I2834: std_logic; attribute dont_touch of I2834: signal is true;
	signal I2839: std_logic; attribute dont_touch of I2839: signal is true;
	signal I2840: std_logic; attribute dont_touch of I2840: signal is true;
	signal I2841: std_logic; attribute dont_touch of I2841: signal is true;
	signal I2842: std_logic; attribute dont_touch of I2842: signal is true;
	signal I2847: std_logic; attribute dont_touch of I2847: signal is true;
	signal I2848: std_logic; attribute dont_touch of I2848: signal is true;
	signal I2849: std_logic; attribute dont_touch of I2849: signal is true;
	signal I2854: std_logic; attribute dont_touch of I2854: signal is true;
	signal I2855: std_logic; attribute dont_touch of I2855: signal is true;
	signal I2856: std_logic; attribute dont_touch of I2856: signal is true;
	signal I2857: std_logic; attribute dont_touch of I2857: signal is true;
	signal I2858: std_logic; attribute dont_touch of I2858: signal is true;
	signal I2863: std_logic; attribute dont_touch of I2863: signal is true;
	signal I2864: std_logic; attribute dont_touch of I2864: signal is true;
	signal I2865: std_logic; attribute dont_touch of I2865: signal is true;
	signal I2870: std_logic; attribute dont_touch of I2870: signal is true;
	signal I2871: std_logic; attribute dont_touch of I2871: signal is true;
	signal I2872: std_logic; attribute dont_touch of I2872: signal is true;
	signal I2873: std_logic; attribute dont_touch of I2873: signal is true;
	signal I2878: std_logic; attribute dont_touch of I2878: signal is true;
	signal I2879: std_logic; attribute dont_touch of I2879: signal is true;
	signal I2880: std_logic; attribute dont_touch of I2880: signal is true;
	signal I2885: std_logic; attribute dont_touch of I2885: signal is true;
	signal I2886: std_logic; attribute dont_touch of I2886: signal is true;
	signal I2887: std_logic; attribute dont_touch of I2887: signal is true;
	signal I2888: std_logic; attribute dont_touch of I2888: signal is true;
	signal I2889: std_logic; attribute dont_touch of I2889: signal is true;
	signal I2894: std_logic; attribute dont_touch of I2894: signal is true;
	signal I2895: std_logic; attribute dont_touch of I2895: signal is true;
	signal I2896: std_logic; attribute dont_touch of I2896: signal is true;
	signal I2901: std_logic; attribute dont_touch of I2901: signal is true;
	signal I2902: std_logic; attribute dont_touch of I2902: signal is true;
	signal I2903: std_logic; attribute dont_touch of I2903: signal is true;
	signal I2904: std_logic; attribute dont_touch of I2904: signal is true;
	signal I2909: std_logic; attribute dont_touch of I2909: signal is true;
	signal I2910: std_logic; attribute dont_touch of I2910: signal is true;
	signal I2911: std_logic; attribute dont_touch of I2911: signal is true;
	signal I2916: std_logic; attribute dont_touch of I2916: signal is true;
	signal I2917: std_logic; attribute dont_touch of I2917: signal is true;
	signal I2918: std_logic; attribute dont_touch of I2918: signal is true;
	signal I2919: std_logic; attribute dont_touch of I2919: signal is true;
	signal I2920: std_logic; attribute dont_touch of I2920: signal is true;
	signal I2925: std_logic; attribute dont_touch of I2925: signal is true;
	signal I2926: std_logic; attribute dont_touch of I2926: signal is true;
	signal I2927: std_logic; attribute dont_touch of I2927: signal is true;
	signal I2932: std_logic; attribute dont_touch of I2932: signal is true;
	signal I2933: std_logic; attribute dont_touch of I2933: signal is true;
	signal I2934: std_logic; attribute dont_touch of I2934: signal is true;
	signal I2935: std_logic; attribute dont_touch of I2935: signal is true;
	signal I2940: std_logic; attribute dont_touch of I2940: signal is true;
	signal I2941: std_logic; attribute dont_touch of I2941: signal is true;
	signal I2942: std_logic; attribute dont_touch of I2942: signal is true;
	signal I2947: std_logic; attribute dont_touch of I2947: signal is true;
	signal I2948: std_logic; attribute dont_touch of I2948: signal is true;
	signal I2949: std_logic; attribute dont_touch of I2949: signal is true;
	signal I2950: std_logic; attribute dont_touch of I2950: signal is true;
	signal I2951: std_logic; attribute dont_touch of I2951: signal is true;
	signal I2956: std_logic; attribute dont_touch of I2956: signal is true;
	signal I2957: std_logic; attribute dont_touch of I2957: signal is true;
	signal I2958: std_logic; attribute dont_touch of I2958: signal is true;
	signal I2963: std_logic; attribute dont_touch of I2963: signal is true;
	signal I2964: std_logic; attribute dont_touch of I2964: signal is true;
	signal I2965: std_logic; attribute dont_touch of I2965: signal is true;
	signal I2966: std_logic; attribute dont_touch of I2966: signal is true;
	signal I2971: std_logic; attribute dont_touch of I2971: signal is true;
	signal I2972: std_logic; attribute dont_touch of I2972: signal is true;
	signal I2973: std_logic; attribute dont_touch of I2973: signal is true;
	signal I3052: std_logic; attribute dont_touch of I3052: signal is true;
	signal I3053: std_logic; attribute dont_touch of I3053: signal is true;
	signal I3054: std_logic; attribute dont_touch of I3054: signal is true;
	signal I3065: std_logic; attribute dont_touch of I3065: signal is true;
	signal I3066: std_logic; attribute dont_touch of I3066: signal is true;
	signal I3067: std_logic; attribute dont_touch of I3067: signal is true;
	signal I3078: std_logic; attribute dont_touch of I3078: signal is true;
	signal I3079: std_logic; attribute dont_touch of I3079: signal is true;
	signal I3080: std_logic; attribute dont_touch of I3080: signal is true;
	signal I3091: std_logic; attribute dont_touch of I3091: signal is true;
	signal I3092: std_logic; attribute dont_touch of I3092: signal is true;
	signal I3093: std_logic; attribute dont_touch of I3093: signal is true;
	signal I3104: std_logic; attribute dont_touch of I3104: signal is true;
	signal I3105: std_logic; attribute dont_touch of I3105: signal is true;
	signal I3106: std_logic; attribute dont_touch of I3106: signal is true;
	signal I3117: std_logic; attribute dont_touch of I3117: signal is true;
	signal I3118: std_logic; attribute dont_touch of I3118: signal is true;
	signal I3119: std_logic; attribute dont_touch of I3119: signal is true;
	signal I3130: std_logic; attribute dont_touch of I3130: signal is true;
	signal I3131: std_logic; attribute dont_touch of I3131: signal is true;
	signal I3132: std_logic; attribute dont_touch of I3132: signal is true;
	signal I3143: std_logic; attribute dont_touch of I3143: signal is true;
	signal I3144: std_logic; attribute dont_touch of I3144: signal is true;
	signal I3145: std_logic; attribute dont_touch of I3145: signal is true;
	signal I3156: std_logic; attribute dont_touch of I3156: signal is true;
	signal I3157: std_logic; attribute dont_touch of I3157: signal is true;
	signal I3158: std_logic; attribute dont_touch of I3158: signal is true;
	signal I3169: std_logic; attribute dont_touch of I3169: signal is true;
	signal I3170: std_logic; attribute dont_touch of I3170: signal is true;
	signal I3171: std_logic; attribute dont_touch of I3171: signal is true;
	signal I3182: std_logic; attribute dont_touch of I3182: signal is true;
	signal I3183: std_logic; attribute dont_touch of I3183: signal is true;
	signal I3184: std_logic; attribute dont_touch of I3184: signal is true;
	signal I3195: std_logic; attribute dont_touch of I3195: signal is true;
	signal I3196: std_logic; attribute dont_touch of I3196: signal is true;
	signal I3197: std_logic; attribute dont_touch of I3197: signal is true;
	signal I3208: std_logic; attribute dont_touch of I3208: signal is true;
	signal I3209: std_logic; attribute dont_touch of I3209: signal is true;
	signal I3210: std_logic; attribute dont_touch of I3210: signal is true;
	signal I3221: std_logic; attribute dont_touch of I3221: signal is true;
	signal I3222: std_logic; attribute dont_touch of I3222: signal is true;
	signal I3223: std_logic; attribute dont_touch of I3223: signal is true;
	signal I3234: std_logic; attribute dont_touch of I3234: signal is true;
	signal I3235: std_logic; attribute dont_touch of I3235: signal is true;
	signal I3236: std_logic; attribute dont_touch of I3236: signal is true;
	signal I3247: std_logic; attribute dont_touch of I3247: signal is true;
	signal I3248: std_logic; attribute dont_touch of I3248: signal is true;
	signal I3249: std_logic; attribute dont_touch of I3249: signal is true;
	signal I3260: std_logic; attribute dont_touch of I3260: signal is true;
	signal I3261: std_logic; attribute dont_touch of I3261: signal is true;
	signal I3262: std_logic; attribute dont_touch of I3262: signal is true;
	signal I3273: std_logic; attribute dont_touch of I3273: signal is true;
	signal I3274: std_logic; attribute dont_touch of I3274: signal is true;
	signal I3275: std_logic; attribute dont_touch of I3275: signal is true;
	signal I3286: std_logic; attribute dont_touch of I3286: signal is true;
	signal I3287: std_logic; attribute dont_touch of I3287: signal is true;
	signal I3288: std_logic; attribute dont_touch of I3288: signal is true;
	signal I3299: std_logic; attribute dont_touch of I3299: signal is true;
	signal I3300: std_logic; attribute dont_touch of I3300: signal is true;
	signal I3301: std_logic; attribute dont_touch of I3301: signal is true;
	signal I3312: std_logic; attribute dont_touch of I3312: signal is true;
	signal I3313: std_logic; attribute dont_touch of I3313: signal is true;
	signal I3314: std_logic; attribute dont_touch of I3314: signal is true;
	signal I3325: std_logic; attribute dont_touch of I3325: signal is true;
	signal I3326: std_logic; attribute dont_touch of I3326: signal is true;
	signal I3327: std_logic; attribute dont_touch of I3327: signal is true;
	signal I3338: std_logic; attribute dont_touch of I3338: signal is true;
	signal I3339: std_logic; attribute dont_touch of I3339: signal is true;
	signal I3340: std_logic; attribute dont_touch of I3340: signal is true;
	signal I3351: std_logic; attribute dont_touch of I3351: signal is true;
	signal I3352: std_logic; attribute dont_touch of I3352: signal is true;
	signal I3353: std_logic; attribute dont_touch of I3353: signal is true;
	signal I3364: std_logic; attribute dont_touch of I3364: signal is true;
	signal I3365: std_logic; attribute dont_touch of I3365: signal is true;
	signal I3366: std_logic; attribute dont_touch of I3366: signal is true;
	signal I3377: std_logic; attribute dont_touch of I3377: signal is true;
	signal I3378: std_logic; attribute dont_touch of I3378: signal is true;
	signal I3379: std_logic; attribute dont_touch of I3379: signal is true;
	signal I3390: std_logic; attribute dont_touch of I3390: signal is true;
	signal I3391: std_logic; attribute dont_touch of I3391: signal is true;
	signal I3392: std_logic; attribute dont_touch of I3392: signal is true;
	signal I3403: std_logic; attribute dont_touch of I3403: signal is true;
	signal I3404: std_logic; attribute dont_touch of I3404: signal is true;
	signal I3405: std_logic; attribute dont_touch of I3405: signal is true;
	signal I3416: std_logic; attribute dont_touch of I3416: signal is true;
	signal I3417: std_logic; attribute dont_touch of I3417: signal is true;
	signal I3418: std_logic; attribute dont_touch of I3418: signal is true;
	signal I3429: std_logic; attribute dont_touch of I3429: signal is true;
	signal I3430: std_logic; attribute dont_touch of I3430: signal is true;
	signal I3431: std_logic; attribute dont_touch of I3431: signal is true;
	signal I3442: std_logic; attribute dont_touch of I3442: signal is true;
	signal I3443: std_logic; attribute dont_touch of I3443: signal is true;
	signal I3444: std_logic; attribute dont_touch of I3444: signal is true;
	signal I3455: std_logic; attribute dont_touch of I3455: signal is true;
	signal I3456: std_logic; attribute dont_touch of I3456: signal is true;
	signal I3457: std_logic; attribute dont_touch of I3457: signal is true;
	signal I3469: std_logic; attribute dont_touch of I3469: signal is true;
	signal I3470: std_logic; attribute dont_touch of I3470: signal is true;
	signal I3471: std_logic; attribute dont_touch of I3471: signal is true;
	signal I3472: std_logic; attribute dont_touch of I3472: signal is true;
	signal I3477: std_logic; attribute dont_touch of I3477: signal is true;
	signal I3478: std_logic; attribute dont_touch of I3478: signal is true;
	signal I3479: std_logic; attribute dont_touch of I3479: signal is true;
	signal I3484: std_logic; attribute dont_touch of I3484: signal is true;
	signal I3485: std_logic; attribute dont_touch of I3485: signal is true;
	signal I3486: std_logic; attribute dont_touch of I3486: signal is true;
	signal I3487: std_logic; attribute dont_touch of I3487: signal is true;
	signal I3492: std_logic; attribute dont_touch of I3492: signal is true;
	signal I3493: std_logic; attribute dont_touch of I3493: signal is true;
	signal I3494: std_logic; attribute dont_touch of I3494: signal is true;
	signal I3499: std_logic; attribute dont_touch of I3499: signal is true;
	signal I3500: std_logic; attribute dont_touch of I3500: signal is true;
	signal I3501: std_logic; attribute dont_touch of I3501: signal is true;
	signal I3502: std_logic; attribute dont_touch of I3502: signal is true;
	signal I3507: std_logic; attribute dont_touch of I3507: signal is true;
	signal I3508: std_logic; attribute dont_touch of I3508: signal is true;
	signal I3509: std_logic; attribute dont_touch of I3509: signal is true;
	signal I3514: std_logic; attribute dont_touch of I3514: signal is true;
	signal I3515: std_logic; attribute dont_touch of I3515: signal is true;
	signal I3516: std_logic; attribute dont_touch of I3516: signal is true;
	signal I3521: std_logic; attribute dont_touch of I3521: signal is true;
	signal I3522: std_logic; attribute dont_touch of I3522: signal is true;
	signal I3523: std_logic; attribute dont_touch of I3523: signal is true;
	signal I3528: std_logic; attribute dont_touch of I3528: signal is true;
	signal I3529: std_logic; attribute dont_touch of I3529: signal is true;
	signal I3530: std_logic; attribute dont_touch of I3530: signal is true;
	signal I3535: std_logic; attribute dont_touch of I3535: signal is true;
	signal I3536: std_logic; attribute dont_touch of I3536: signal is true;
	signal I3537: std_logic; attribute dont_touch of I3537: signal is true;
	signal I3542: std_logic; attribute dont_touch of I3542: signal is true;
	signal I3543: std_logic; attribute dont_touch of I3543: signal is true;
	signal I3544: std_logic; attribute dont_touch of I3544: signal is true;
	signal I3549: std_logic; attribute dont_touch of I3549: signal is true;
	signal I3550: std_logic; attribute dont_touch of I3550: signal is true;
	signal I3551: std_logic; attribute dont_touch of I3551: signal is true;
	signal I3556: std_logic; attribute dont_touch of I3556: signal is true;
	signal I3557: std_logic; attribute dont_touch of I3557: signal is true;
	signal I3558: std_logic; attribute dont_touch of I3558: signal is true;
	signal I3563: std_logic; attribute dont_touch of I3563: signal is true;
	signal I3564: std_logic; attribute dont_touch of I3564: signal is true;
	signal I3565: std_logic; attribute dont_touch of I3565: signal is true;
	signal I3570: std_logic; attribute dont_touch of I3570: signal is true;
	signal I3571: std_logic; attribute dont_touch of I3571: signal is true;
	signal I3572: std_logic; attribute dont_touch of I3572: signal is true;
	signal I3577: std_logic; attribute dont_touch of I3577: signal is true;
	signal I3578: std_logic; attribute dont_touch of I3578: signal is true;
	signal I3579: std_logic; attribute dont_touch of I3579: signal is true;
	signal I3584: std_logic; attribute dont_touch of I3584: signal is true;
	signal I3585: std_logic; attribute dont_touch of I3585: signal is true;
	signal I3586: std_logic; attribute dont_touch of I3586: signal is true;
	signal I3591: std_logic; attribute dont_touch of I3591: signal is true;
	signal I3592: std_logic; attribute dont_touch of I3592: signal is true;
	signal I3593: std_logic; attribute dont_touch of I3593: signal is true;
	signal I3598: std_logic; attribute dont_touch of I3598: signal is true;
	signal I3599: std_logic; attribute dont_touch of I3599: signal is true;
	signal I3600: std_logic; attribute dont_touch of I3600: signal is true;
	signal I3605: std_logic; attribute dont_touch of I3605: signal is true;
	signal I3606: std_logic; attribute dont_touch of I3606: signal is true;
	signal I3607: std_logic; attribute dont_touch of I3607: signal is true;
	signal I3612: std_logic; attribute dont_touch of I3612: signal is true;
	signal I3613: std_logic; attribute dont_touch of I3613: signal is true;
	signal I3614: std_logic; attribute dont_touch of I3614: signal is true;
	signal I3619: std_logic; attribute dont_touch of I3619: signal is true;
	signal I3620: std_logic; attribute dont_touch of I3620: signal is true;
	signal I3621: std_logic; attribute dont_touch of I3621: signal is true;
	signal I3626: std_logic; attribute dont_touch of I3626: signal is true;
	signal I3627: std_logic; attribute dont_touch of I3627: signal is true;
	signal I3628: std_logic; attribute dont_touch of I3628: signal is true;
	signal I3633: std_logic; attribute dont_touch of I3633: signal is true;
	signal I3634: std_logic; attribute dont_touch of I3634: signal is true;
	signal I3635: std_logic; attribute dont_touch of I3635: signal is true;
	signal I3640: std_logic; attribute dont_touch of I3640: signal is true;
	signal I3641: std_logic; attribute dont_touch of I3641: signal is true;
	signal I3642: std_logic; attribute dont_touch of I3642: signal is true;
	signal I3647: std_logic; attribute dont_touch of I3647: signal is true;
	signal I3648: std_logic; attribute dont_touch of I3648: signal is true;
	signal I3649: std_logic; attribute dont_touch of I3649: signal is true;
	signal I3654: std_logic; attribute dont_touch of I3654: signal is true;
	signal I3655: std_logic; attribute dont_touch of I3655: signal is true;
	signal I3656: std_logic; attribute dont_touch of I3656: signal is true;
	signal I3661: std_logic; attribute dont_touch of I3661: signal is true;
	signal I3662: std_logic; attribute dont_touch of I3662: signal is true;
	signal I3663: std_logic; attribute dont_touch of I3663: signal is true;
	signal I3668: std_logic; attribute dont_touch of I3668: signal is true;
	signal I3669: std_logic; attribute dont_touch of I3669: signal is true;
	signal I3670: std_logic; attribute dont_touch of I3670: signal is true;
	signal I3675: std_logic; attribute dont_touch of I3675: signal is true;
	signal I3676: std_logic; attribute dont_touch of I3676: signal is true;
	signal I3677: std_logic; attribute dont_touch of I3677: signal is true;
	signal I3682: std_logic; attribute dont_touch of I3682: signal is true;
	signal I3683: std_logic; attribute dont_touch of I3683: signal is true;
	signal I3684: std_logic; attribute dont_touch of I3684: signal is true;
	signal I3689: std_logic; attribute dont_touch of I3689: signal is true;
	signal I3690: std_logic; attribute dont_touch of I3690: signal is true;
	signal I3691: std_logic; attribute dont_touch of I3691: signal is true;
	signal I3696: std_logic; attribute dont_touch of I3696: signal is true;
	signal I3697: std_logic; attribute dont_touch of I3697: signal is true;
	signal I3698: std_logic; attribute dont_touch of I3698: signal is true;
	signal I3703: std_logic; attribute dont_touch of I3703: signal is true;
	signal I3704: std_logic; attribute dont_touch of I3704: signal is true;
	signal I3705: std_logic; attribute dont_touch of I3705: signal is true;
	signal I3710: std_logic; attribute dont_touch of I3710: signal is true;
	signal I3711: std_logic; attribute dont_touch of I3711: signal is true;
	signal I3712: std_logic; attribute dont_touch of I3712: signal is true;
	signal I5991: std_logic; attribute dont_touch of I5991: signal is true;
	signal I5992: std_logic; attribute dont_touch of I5992: signal is true;
	signal I5993: std_logic; attribute dont_touch of I5993: signal is true;
	signal I5994: std_logic; attribute dont_touch of I5994: signal is true;
	signal I5995: std_logic; attribute dont_touch of I5995: signal is true;
	signal I6000: std_logic; attribute dont_touch of I6000: signal is true;
	signal I6001: std_logic; attribute dont_touch of I6001: signal is true;
	signal I6002: std_logic; attribute dont_touch of I6002: signal is true;
	signal I6007: std_logic; attribute dont_touch of I6007: signal is true;
	signal I6008: std_logic; attribute dont_touch of I6008: signal is true;
	signal I6009: std_logic; attribute dont_touch of I6009: signal is true;
	signal I6010: std_logic; attribute dont_touch of I6010: signal is true;
	signal I6015: std_logic; attribute dont_touch of I6015: signal is true;
	signal I6016: std_logic; attribute dont_touch of I6016: signal is true;
	signal I6017: std_logic; attribute dont_touch of I6017: signal is true;
	signal I6022: std_logic; attribute dont_touch of I6022: signal is true;
	signal I6023: std_logic; attribute dont_touch of I6023: signal is true;
	signal I6024: std_logic; attribute dont_touch of I6024: signal is true;
	signal I6025: std_logic; attribute dont_touch of I6025: signal is true;
	signal I6026: std_logic; attribute dont_touch of I6026: signal is true;
	signal I6031: std_logic; attribute dont_touch of I6031: signal is true;
	signal I6032: std_logic; attribute dont_touch of I6032: signal is true;
	signal I6033: std_logic; attribute dont_touch of I6033: signal is true;
	signal I6038: std_logic; attribute dont_touch of I6038: signal is true;
	signal I6039: std_logic; attribute dont_touch of I6039: signal is true;
	signal I6040: std_logic; attribute dont_touch of I6040: signal is true;
	signal I6041: std_logic; attribute dont_touch of I6041: signal is true;
	signal I6046: std_logic; attribute dont_touch of I6046: signal is true;
	signal I6047: std_logic; attribute dont_touch of I6047: signal is true;
	signal I6048: std_logic; attribute dont_touch of I6048: signal is true;
	signal I6053: std_logic; attribute dont_touch of I6053: signal is true;
	signal I6054: std_logic; attribute dont_touch of I6054: signal is true;
	signal I6055: std_logic; attribute dont_touch of I6055: signal is true;
	signal I6056: std_logic; attribute dont_touch of I6056: signal is true;
	signal I6057: std_logic; attribute dont_touch of I6057: signal is true;
	signal I6062: std_logic; attribute dont_touch of I6062: signal is true;
	signal I6063: std_logic; attribute dont_touch of I6063: signal is true;
	signal I6064: std_logic; attribute dont_touch of I6064: signal is true;
	signal I6069: std_logic; attribute dont_touch of I6069: signal is true;
	signal I6070: std_logic; attribute dont_touch of I6070: signal is true;
	signal I6071: std_logic; attribute dont_touch of I6071: signal is true;
	signal I6072: std_logic; attribute dont_touch of I6072: signal is true;
	signal I6077: std_logic; attribute dont_touch of I6077: signal is true;
	signal I6078: std_logic; attribute dont_touch of I6078: signal is true;
	signal I6079: std_logic; attribute dont_touch of I6079: signal is true;
	signal I6084: std_logic; attribute dont_touch of I6084: signal is true;
	signal I6085: std_logic; attribute dont_touch of I6085: signal is true;
	signal I6086: std_logic; attribute dont_touch of I6086: signal is true;
	signal I6087: std_logic; attribute dont_touch of I6087: signal is true;
	signal I6088: std_logic; attribute dont_touch of I6088: signal is true;
	signal I6093: std_logic; attribute dont_touch of I6093: signal is true;
	signal I6094: std_logic; attribute dont_touch of I6094: signal is true;
	signal I6095: std_logic; attribute dont_touch of I6095: signal is true;
	signal I6100: std_logic; attribute dont_touch of I6100: signal is true;
	signal I6101: std_logic; attribute dont_touch of I6101: signal is true;
	signal I6102: std_logic; attribute dont_touch of I6102: signal is true;
	signal I6103: std_logic; attribute dont_touch of I6103: signal is true;
	signal I6108: std_logic; attribute dont_touch of I6108: signal is true;
	signal I6109: std_logic; attribute dont_touch of I6109: signal is true;
	signal I6110: std_logic; attribute dont_touch of I6110: signal is true;
	signal I6115: std_logic; attribute dont_touch of I6115: signal is true;
	signal I6116: std_logic; attribute dont_touch of I6116: signal is true;
	signal I6117: std_logic; attribute dont_touch of I6117: signal is true;
	signal I6118: std_logic; attribute dont_touch of I6118: signal is true;
	signal I6119: std_logic; attribute dont_touch of I6119: signal is true;
	signal I6124: std_logic; attribute dont_touch of I6124: signal is true;
	signal I6125: std_logic; attribute dont_touch of I6125: signal is true;
	signal I6126: std_logic; attribute dont_touch of I6126: signal is true;
	signal I6131: std_logic; attribute dont_touch of I6131: signal is true;
	signal I6132: std_logic; attribute dont_touch of I6132: signal is true;
	signal I6133: std_logic; attribute dont_touch of I6133: signal is true;
	signal I6134: std_logic; attribute dont_touch of I6134: signal is true;
	signal I6139: std_logic; attribute dont_touch of I6139: signal is true;
	signal I6140: std_logic; attribute dont_touch of I6140: signal is true;
	signal I6141: std_logic; attribute dont_touch of I6141: signal is true;
	signal I6146: std_logic; attribute dont_touch of I6146: signal is true;
	signal I6147: std_logic; attribute dont_touch of I6147: signal is true;
	signal I6148: std_logic; attribute dont_touch of I6148: signal is true;
	signal I6149: std_logic; attribute dont_touch of I6149: signal is true;
	signal I6150: std_logic; attribute dont_touch of I6150: signal is true;
	signal I6155: std_logic; attribute dont_touch of I6155: signal is true;
	signal I6156: std_logic; attribute dont_touch of I6156: signal is true;
	signal I6157: std_logic; attribute dont_touch of I6157: signal is true;
	signal I6162: std_logic; attribute dont_touch of I6162: signal is true;
	signal I6163: std_logic; attribute dont_touch of I6163: signal is true;
	signal I6164: std_logic; attribute dont_touch of I6164: signal is true;
	signal I6165: std_logic; attribute dont_touch of I6165: signal is true;
	signal I6170: std_logic; attribute dont_touch of I6170: signal is true;
	signal I6171: std_logic; attribute dont_touch of I6171: signal is true;
	signal I6172: std_logic; attribute dont_touch of I6172: signal is true;
	signal I6177: std_logic; attribute dont_touch of I6177: signal is true;
	signal I6178: std_logic; attribute dont_touch of I6178: signal is true;
	signal I6179: std_logic; attribute dont_touch of I6179: signal is true;
	signal I6180: std_logic; attribute dont_touch of I6180: signal is true;
	signal I6181: std_logic; attribute dont_touch of I6181: signal is true;
	signal I6186: std_logic; attribute dont_touch of I6186: signal is true;
	signal I6187: std_logic; attribute dont_touch of I6187: signal is true;
	signal I6188: std_logic; attribute dont_touch of I6188: signal is true;
	signal I6193: std_logic; attribute dont_touch of I6193: signal is true;
	signal I6194: std_logic; attribute dont_touch of I6194: signal is true;
	signal I6195: std_logic; attribute dont_touch of I6195: signal is true;
	signal I6196: std_logic; attribute dont_touch of I6196: signal is true;
	signal I6201: std_logic; attribute dont_touch of I6201: signal is true;
	signal I6202: std_logic; attribute dont_touch of I6202: signal is true;
	signal I6203: std_logic; attribute dont_touch of I6203: signal is true;
	signal I6208: std_logic; attribute dont_touch of I6208: signal is true;
	signal I6209: std_logic; attribute dont_touch of I6209: signal is true;
	signal I6210: std_logic; attribute dont_touch of I6210: signal is true;
	signal I6211: std_logic; attribute dont_touch of I6211: signal is true;
	signal I6212: std_logic; attribute dont_touch of I6212: signal is true;
	signal I6217: std_logic; attribute dont_touch of I6217: signal is true;
	signal I6218: std_logic; attribute dont_touch of I6218: signal is true;
	signal I6219: std_logic; attribute dont_touch of I6219: signal is true;
	signal I6224: std_logic; attribute dont_touch of I6224: signal is true;
	signal I6225: std_logic; attribute dont_touch of I6225: signal is true;
	signal I6226: std_logic; attribute dont_touch of I6226: signal is true;
	signal I6227: std_logic; attribute dont_touch of I6227: signal is true;
	signal I6232: std_logic; attribute dont_touch of I6232: signal is true;
	signal I6233: std_logic; attribute dont_touch of I6233: signal is true;
	signal I6234: std_logic; attribute dont_touch of I6234: signal is true;
	signal I6239: std_logic; attribute dont_touch of I6239: signal is true;
	signal I6240: std_logic; attribute dont_touch of I6240: signal is true;
	signal I6241: std_logic; attribute dont_touch of I6241: signal is true;
	signal I6242: std_logic; attribute dont_touch of I6242: signal is true;
	signal I6243: std_logic; attribute dont_touch of I6243: signal is true;
	signal I6248: std_logic; attribute dont_touch of I6248: signal is true;
	signal I6249: std_logic; attribute dont_touch of I6249: signal is true;
	signal I6250: std_logic; attribute dont_touch of I6250: signal is true;
	signal I6255: std_logic; attribute dont_touch of I6255: signal is true;
	signal I6256: std_logic; attribute dont_touch of I6256: signal is true;
	signal I6257: std_logic; attribute dont_touch of I6257: signal is true;
	signal I6258: std_logic; attribute dont_touch of I6258: signal is true;
	signal I6263: std_logic; attribute dont_touch of I6263: signal is true;
	signal I6264: std_logic; attribute dont_touch of I6264: signal is true;
	signal I6265: std_logic; attribute dont_touch of I6265: signal is true;
	signal I6270: std_logic; attribute dont_touch of I6270: signal is true;
	signal I6271: std_logic; attribute dont_touch of I6271: signal is true;
	signal I6272: std_logic; attribute dont_touch of I6272: signal is true;
	signal I6273: std_logic; attribute dont_touch of I6273: signal is true;
	signal I6274: std_logic; attribute dont_touch of I6274: signal is true;
	signal I6279: std_logic; attribute dont_touch of I6279: signal is true;
	signal I6280: std_logic; attribute dont_touch of I6280: signal is true;
	signal I6281: std_logic; attribute dont_touch of I6281: signal is true;
	signal I6286: std_logic; attribute dont_touch of I6286: signal is true;
	signal I6287: std_logic; attribute dont_touch of I6287: signal is true;
	signal I6288: std_logic; attribute dont_touch of I6288: signal is true;
	signal I6289: std_logic; attribute dont_touch of I6289: signal is true;
	signal I6294: std_logic; attribute dont_touch of I6294: signal is true;
	signal I6295: std_logic; attribute dont_touch of I6295: signal is true;
	signal I6296: std_logic; attribute dont_touch of I6296: signal is true;
	signal I6301: std_logic; attribute dont_touch of I6301: signal is true;
	signal I6302: std_logic; attribute dont_touch of I6302: signal is true;
	signal I6303: std_logic; attribute dont_touch of I6303: signal is true;
	signal I6304: std_logic; attribute dont_touch of I6304: signal is true;
	signal I6305: std_logic; attribute dont_touch of I6305: signal is true;
	signal I6310: std_logic; attribute dont_touch of I6310: signal is true;
	signal I6311: std_logic; attribute dont_touch of I6311: signal is true;
	signal I6312: std_logic; attribute dont_touch of I6312: signal is true;
	signal I6317: std_logic; attribute dont_touch of I6317: signal is true;
	signal I6318: std_logic; attribute dont_touch of I6318: signal is true;
	signal I6319: std_logic; attribute dont_touch of I6319: signal is true;
	signal I6320: std_logic; attribute dont_touch of I6320: signal is true;
	signal I6325: std_logic; attribute dont_touch of I6325: signal is true;
	signal I6326: std_logic; attribute dont_touch of I6326: signal is true;
	signal I6327: std_logic; attribute dont_touch of I6327: signal is true;
	signal I6332: std_logic; attribute dont_touch of I6332: signal is true;
	signal I6333: std_logic; attribute dont_touch of I6333: signal is true;
	signal I6334: std_logic; attribute dont_touch of I6334: signal is true;
	signal I6335: std_logic; attribute dont_touch of I6335: signal is true;
	signal I6336: std_logic; attribute dont_touch of I6336: signal is true;
	signal I6341: std_logic; attribute dont_touch of I6341: signal is true;
	signal I6342: std_logic; attribute dont_touch of I6342: signal is true;
	signal I6343: std_logic; attribute dont_touch of I6343: signal is true;
	signal I6348: std_logic; attribute dont_touch of I6348: signal is true;
	signal I6349: std_logic; attribute dont_touch of I6349: signal is true;
	signal I6350: std_logic; attribute dont_touch of I6350: signal is true;
	signal I6351: std_logic; attribute dont_touch of I6351: signal is true;
	signal I6356: std_logic; attribute dont_touch of I6356: signal is true;
	signal I6357: std_logic; attribute dont_touch of I6357: signal is true;
	signal I6358: std_logic; attribute dont_touch of I6358: signal is true;
	signal I6363: std_logic; attribute dont_touch of I6363: signal is true;
	signal I6364: std_logic; attribute dont_touch of I6364: signal is true;
	signal I6365: std_logic; attribute dont_touch of I6365: signal is true;
	signal I6366: std_logic; attribute dont_touch of I6366: signal is true;
	signal I6367: std_logic; attribute dont_touch of I6367: signal is true;
	signal I6372: std_logic; attribute dont_touch of I6372: signal is true;
	signal I6373: std_logic; attribute dont_touch of I6373: signal is true;
	signal I6374: std_logic; attribute dont_touch of I6374: signal is true;
	signal I6379: std_logic; attribute dont_touch of I6379: signal is true;
	signal I6380: std_logic; attribute dont_touch of I6380: signal is true;
	signal I6381: std_logic; attribute dont_touch of I6381: signal is true;
	signal I6382: std_logic; attribute dont_touch of I6382: signal is true;
	signal I6387: std_logic; attribute dont_touch of I6387: signal is true;
	signal I6388: std_logic; attribute dont_touch of I6388: signal is true;
	signal I6389: std_logic; attribute dont_touch of I6389: signal is true;
	signal I6394: std_logic; attribute dont_touch of I6394: signal is true;
	signal I6395: std_logic; attribute dont_touch of I6395: signal is true;
	signal I6396: std_logic; attribute dont_touch of I6396: signal is true;
	signal I6397: std_logic; attribute dont_touch of I6397: signal is true;
	signal I6398: std_logic; attribute dont_touch of I6398: signal is true;
	signal I6403: std_logic; attribute dont_touch of I6403: signal is true;
	signal I6404: std_logic; attribute dont_touch of I6404: signal is true;
	signal I6405: std_logic; attribute dont_touch of I6405: signal is true;
	signal I6410: std_logic; attribute dont_touch of I6410: signal is true;
	signal I6411: std_logic; attribute dont_touch of I6411: signal is true;
	signal I6412: std_logic; attribute dont_touch of I6412: signal is true;
	signal I6413: std_logic; attribute dont_touch of I6413: signal is true;
	signal I6418: std_logic; attribute dont_touch of I6418: signal is true;
	signal I6419: std_logic; attribute dont_touch of I6419: signal is true;
	signal I6420: std_logic; attribute dont_touch of I6420: signal is true;
	signal I6425: std_logic; attribute dont_touch of I6425: signal is true;
	signal I6426: std_logic; attribute dont_touch of I6426: signal is true;
	signal I6427: std_logic; attribute dont_touch of I6427: signal is true;
	signal I6428: std_logic; attribute dont_touch of I6428: signal is true;
	signal I6429: std_logic; attribute dont_touch of I6429: signal is true;
	signal I6434: std_logic; attribute dont_touch of I6434: signal is true;
	signal I6435: std_logic; attribute dont_touch of I6435: signal is true;
	signal I6436: std_logic; attribute dont_touch of I6436: signal is true;
	signal I6441: std_logic; attribute dont_touch of I6441: signal is true;
	signal I6442: std_logic; attribute dont_touch of I6442: signal is true;
	signal I6443: std_logic; attribute dont_touch of I6443: signal is true;
	signal I6444: std_logic; attribute dont_touch of I6444: signal is true;
	signal I6449: std_logic; attribute dont_touch of I6449: signal is true;
	signal I6450: std_logic; attribute dont_touch of I6450: signal is true;
	signal I6451: std_logic; attribute dont_touch of I6451: signal is true;
	signal I6456: std_logic; attribute dont_touch of I6456: signal is true;
	signal I6457: std_logic; attribute dont_touch of I6457: signal is true;
	signal I6458: std_logic; attribute dont_touch of I6458: signal is true;
	signal I6459: std_logic; attribute dont_touch of I6459: signal is true;
	signal I6460: std_logic; attribute dont_touch of I6460: signal is true;
	signal I6465: std_logic; attribute dont_touch of I6465: signal is true;
	signal I6466: std_logic; attribute dont_touch of I6466: signal is true;
	signal I6467: std_logic; attribute dont_touch of I6467: signal is true;
	signal I6472: std_logic; attribute dont_touch of I6472: signal is true;
	signal I6473: std_logic; attribute dont_touch of I6473: signal is true;
	signal I6474: std_logic; attribute dont_touch of I6474: signal is true;
	signal I6475: std_logic; attribute dont_touch of I6475: signal is true;
	signal I6480: std_logic; attribute dont_touch of I6480: signal is true;
	signal I6481: std_logic; attribute dont_touch of I6481: signal is true;
	signal I6482: std_logic; attribute dont_touch of I6482: signal is true;
	signal I6487: std_logic; attribute dont_touch of I6487: signal is true;
	signal I6488: std_logic; attribute dont_touch of I6488: signal is true;
	signal I6489: std_logic; attribute dont_touch of I6489: signal is true;
	signal I6490: std_logic; attribute dont_touch of I6490: signal is true;
	signal I6491: std_logic; attribute dont_touch of I6491: signal is true;
	signal I6496: std_logic; attribute dont_touch of I6496: signal is true;
	signal I6497: std_logic; attribute dont_touch of I6497: signal is true;
	signal I6498: std_logic; attribute dont_touch of I6498: signal is true;
	signal I6503: std_logic; attribute dont_touch of I6503: signal is true;
	signal I6504: std_logic; attribute dont_touch of I6504: signal is true;
	signal I6505: std_logic; attribute dont_touch of I6505: signal is true;
	signal I6506: std_logic; attribute dont_touch of I6506: signal is true;
	signal I6511: std_logic; attribute dont_touch of I6511: signal is true;
	signal I6512: std_logic; attribute dont_touch of I6512: signal is true;
	signal I6513: std_logic; attribute dont_touch of I6513: signal is true;
	signal I6518: std_logic; attribute dont_touch of I6518: signal is true;
	signal I6519: std_logic; attribute dont_touch of I6519: signal is true;
	signal I6520: std_logic; attribute dont_touch of I6520: signal is true;
	signal I6521: std_logic; attribute dont_touch of I6521: signal is true;
	signal I6522: std_logic; attribute dont_touch of I6522: signal is true;
	signal I6527: std_logic; attribute dont_touch of I6527: signal is true;
	signal I6528: std_logic; attribute dont_touch of I6528: signal is true;
	signal I6529: std_logic; attribute dont_touch of I6529: signal is true;
	signal I6534: std_logic; attribute dont_touch of I6534: signal is true;
	signal I6535: std_logic; attribute dont_touch of I6535: signal is true;
	signal I6536: std_logic; attribute dont_touch of I6536: signal is true;
	signal I6537: std_logic; attribute dont_touch of I6537: signal is true;
	signal I6542: std_logic; attribute dont_touch of I6542: signal is true;
	signal I6543: std_logic; attribute dont_touch of I6543: signal is true;
	signal I6544: std_logic; attribute dont_touch of I6544: signal is true;
	signal I6549: std_logic; attribute dont_touch of I6549: signal is true;
	signal I6550: std_logic; attribute dont_touch of I6550: signal is true;
	signal I6551: std_logic; attribute dont_touch of I6551: signal is true;
	signal I6552: std_logic; attribute dont_touch of I6552: signal is true;
	signal I6553: std_logic; attribute dont_touch of I6553: signal is true;
	signal I6558: std_logic; attribute dont_touch of I6558: signal is true;
	signal I6559: std_logic; attribute dont_touch of I6559: signal is true;
	signal I6560: std_logic; attribute dont_touch of I6560: signal is true;
	signal I6565: std_logic; attribute dont_touch of I6565: signal is true;
	signal I6566: std_logic; attribute dont_touch of I6566: signal is true;
	signal I6567: std_logic; attribute dont_touch of I6567: signal is true;
	signal I6568: std_logic; attribute dont_touch of I6568: signal is true;
	signal I6573: std_logic; attribute dont_touch of I6573: signal is true;
	signal I6574: std_logic; attribute dont_touch of I6574: signal is true;
	signal I6575: std_logic; attribute dont_touch of I6575: signal is true;
	signal I6580: std_logic; attribute dont_touch of I6580: signal is true;
	signal I6581: std_logic; attribute dont_touch of I6581: signal is true;
	signal I6582: std_logic; attribute dont_touch of I6582: signal is true;
	signal I6583: std_logic; attribute dont_touch of I6583: signal is true;
	signal I6584: std_logic; attribute dont_touch of I6584: signal is true;
	signal I6589: std_logic; attribute dont_touch of I6589: signal is true;
	signal I6590: std_logic; attribute dont_touch of I6590: signal is true;
	signal I6591: std_logic; attribute dont_touch of I6591: signal is true;
	signal I6596: std_logic; attribute dont_touch of I6596: signal is true;
	signal I6597: std_logic; attribute dont_touch of I6597: signal is true;
	signal I6598: std_logic; attribute dont_touch of I6598: signal is true;
	signal I6599: std_logic; attribute dont_touch of I6599: signal is true;
	signal I6604: std_logic; attribute dont_touch of I6604: signal is true;
	signal I6605: std_logic; attribute dont_touch of I6605: signal is true;
	signal I6606: std_logic; attribute dont_touch of I6606: signal is true;
	signal I6611: std_logic; attribute dont_touch of I6611: signal is true;
	signal I6612: std_logic; attribute dont_touch of I6612: signal is true;
	signal I6613: std_logic; attribute dont_touch of I6613: signal is true;
	signal I6614: std_logic; attribute dont_touch of I6614: signal is true;
	signal I6615: std_logic; attribute dont_touch of I6615: signal is true;
	signal I6620: std_logic; attribute dont_touch of I6620: signal is true;
	signal I6621: std_logic; attribute dont_touch of I6621: signal is true;
	signal I6622: std_logic; attribute dont_touch of I6622: signal is true;
	signal I6627: std_logic; attribute dont_touch of I6627: signal is true;
	signal I6628: std_logic; attribute dont_touch of I6628: signal is true;
	signal I6629: std_logic; attribute dont_touch of I6629: signal is true;
	signal I6630: std_logic; attribute dont_touch of I6630: signal is true;
	signal I6635: std_logic; attribute dont_touch of I6635: signal is true;
	signal I6636: std_logic; attribute dont_touch of I6636: signal is true;
	signal I6637: std_logic; attribute dont_touch of I6637: signal is true;
	signal I6642: std_logic; attribute dont_touch of I6642: signal is true;
	signal I6643: std_logic; attribute dont_touch of I6643: signal is true;
	signal I6644: std_logic; attribute dont_touch of I6644: signal is true;
	signal I6645: std_logic; attribute dont_touch of I6645: signal is true;
	signal I6646: std_logic; attribute dont_touch of I6646: signal is true;
	signal I6651: std_logic; attribute dont_touch of I6651: signal is true;
	signal I6652: std_logic; attribute dont_touch of I6652: signal is true;
	signal I6653: std_logic; attribute dont_touch of I6653: signal is true;
	signal I6658: std_logic; attribute dont_touch of I6658: signal is true;
	signal I6659: std_logic; attribute dont_touch of I6659: signal is true;
	signal I6660: std_logic; attribute dont_touch of I6660: signal is true;
	signal I6661: std_logic; attribute dont_touch of I6661: signal is true;
	signal I6666: std_logic; attribute dont_touch of I6666: signal is true;
	signal I6667: std_logic; attribute dont_touch of I6667: signal is true;
	signal I6668: std_logic; attribute dont_touch of I6668: signal is true;
	signal I6673: std_logic; attribute dont_touch of I6673: signal is true;
	signal I6674: std_logic; attribute dont_touch of I6674: signal is true;
	signal I6675: std_logic; attribute dont_touch of I6675: signal is true;
	signal I6676: std_logic; attribute dont_touch of I6676: signal is true;
	signal I6677: std_logic; attribute dont_touch of I6677: signal is true;
	signal I6682: std_logic; attribute dont_touch of I6682: signal is true;
	signal I6683: std_logic; attribute dont_touch of I6683: signal is true;
	signal I6684: std_logic; attribute dont_touch of I6684: signal is true;
	signal I6689: std_logic; attribute dont_touch of I6689: signal is true;
	signal I6690: std_logic; attribute dont_touch of I6690: signal is true;
	signal I6691: std_logic; attribute dont_touch of I6691: signal is true;
	signal I6692: std_logic; attribute dont_touch of I6692: signal is true;
	signal I6697: std_logic; attribute dont_touch of I6697: signal is true;
	signal I6698: std_logic; attribute dont_touch of I6698: signal is true;
	signal I6699: std_logic; attribute dont_touch of I6699: signal is true;
	signal I6704: std_logic; attribute dont_touch of I6704: signal is true;
	signal I6705: std_logic; attribute dont_touch of I6705: signal is true;
	signal I6706: std_logic; attribute dont_touch of I6706: signal is true;
	signal I6707: std_logic; attribute dont_touch of I6707: signal is true;
	signal I6708: std_logic; attribute dont_touch of I6708: signal is true;
	signal I6713: std_logic; attribute dont_touch of I6713: signal is true;
	signal I6714: std_logic; attribute dont_touch of I6714: signal is true;
	signal I6715: std_logic; attribute dont_touch of I6715: signal is true;
	signal I6720: std_logic; attribute dont_touch of I6720: signal is true;
	signal I6721: std_logic; attribute dont_touch of I6721: signal is true;
	signal I6722: std_logic; attribute dont_touch of I6722: signal is true;
	signal I6723: std_logic; attribute dont_touch of I6723: signal is true;
	signal I6728: std_logic; attribute dont_touch of I6728: signal is true;
	signal I6729: std_logic; attribute dont_touch of I6729: signal is true;
	signal I6730: std_logic; attribute dont_touch of I6730: signal is true;
	signal I6735: std_logic; attribute dont_touch of I6735: signal is true;
	signal I6736: std_logic; attribute dont_touch of I6736: signal is true;
	signal I6737: std_logic; attribute dont_touch of I6737: signal is true;
	signal I6738: std_logic; attribute dont_touch of I6738: signal is true;
	signal I6739: std_logic; attribute dont_touch of I6739: signal is true;
	signal I6744: std_logic; attribute dont_touch of I6744: signal is true;
	signal I6745: std_logic; attribute dont_touch of I6745: signal is true;
	signal I6746: std_logic; attribute dont_touch of I6746: signal is true;
	signal I6751: std_logic; attribute dont_touch of I6751: signal is true;
	signal I6752: std_logic; attribute dont_touch of I6752: signal is true;
	signal I6753: std_logic; attribute dont_touch of I6753: signal is true;
	signal I6754: std_logic; attribute dont_touch of I6754: signal is true;
	signal I6759: std_logic; attribute dont_touch of I6759: signal is true;
	signal I6760: std_logic; attribute dont_touch of I6760: signal is true;
	signal I6761: std_logic; attribute dont_touch of I6761: signal is true;
	signal I6766: std_logic; attribute dont_touch of I6766: signal is true;
	signal I6767: std_logic; attribute dont_touch of I6767: signal is true;
	signal I6768: std_logic; attribute dont_touch of I6768: signal is true;
	signal I6769: std_logic; attribute dont_touch of I6769: signal is true;
	signal I6770: std_logic; attribute dont_touch of I6770: signal is true;
	signal I6775: std_logic; attribute dont_touch of I6775: signal is true;
	signal I6776: std_logic; attribute dont_touch of I6776: signal is true;
	signal I6777: std_logic; attribute dont_touch of I6777: signal is true;
	signal I6782: std_logic; attribute dont_touch of I6782: signal is true;
	signal I6783: std_logic; attribute dont_touch of I6783: signal is true;
	signal I6784: std_logic; attribute dont_touch of I6784: signal is true;
	signal I6785: std_logic; attribute dont_touch of I6785: signal is true;
	signal I6790: std_logic; attribute dont_touch of I6790: signal is true;
	signal I6791: std_logic; attribute dont_touch of I6791: signal is true;
	signal I6792: std_logic; attribute dont_touch of I6792: signal is true;
	signal I6797: std_logic; attribute dont_touch of I6797: signal is true;
	signal I6798: std_logic; attribute dont_touch of I6798: signal is true;
	signal I6799: std_logic; attribute dont_touch of I6799: signal is true;
	signal I6800: std_logic; attribute dont_touch of I6800: signal is true;
	signal I6801: std_logic; attribute dont_touch of I6801: signal is true;
	signal I6806: std_logic; attribute dont_touch of I6806: signal is true;
	signal I6807: std_logic; attribute dont_touch of I6807: signal is true;
	signal I6808: std_logic; attribute dont_touch of I6808: signal is true;
	signal I6813: std_logic; attribute dont_touch of I6813: signal is true;
	signal I6814: std_logic; attribute dont_touch of I6814: signal is true;
	signal I6815: std_logic; attribute dont_touch of I6815: signal is true;
	signal I6816: std_logic; attribute dont_touch of I6816: signal is true;
	signal I6821: std_logic; attribute dont_touch of I6821: signal is true;
	signal I6822: std_logic; attribute dont_touch of I6822: signal is true;
	signal I6823: std_logic; attribute dont_touch of I6823: signal is true;
	signal I6828: std_logic; attribute dont_touch of I6828: signal is true;
	signal I6829: std_logic; attribute dont_touch of I6829: signal is true;
	signal I6830: std_logic; attribute dont_touch of I6830: signal is true;
	signal I6831: std_logic; attribute dont_touch of I6831: signal is true;
	signal I6832: std_logic; attribute dont_touch of I6832: signal is true;
	signal I6837: std_logic; attribute dont_touch of I6837: signal is true;
	signal I6838: std_logic; attribute dont_touch of I6838: signal is true;
	signal I6839: std_logic; attribute dont_touch of I6839: signal is true;
	signal I6844: std_logic; attribute dont_touch of I6844: signal is true;
	signal I6845: std_logic; attribute dont_touch of I6845: signal is true;
	signal I6846: std_logic; attribute dont_touch of I6846: signal is true;
	signal I6847: std_logic; attribute dont_touch of I6847: signal is true;
	signal I6852: std_logic; attribute dont_touch of I6852: signal is true;
	signal I6853: std_logic; attribute dont_touch of I6853: signal is true;
	signal I6854: std_logic; attribute dont_touch of I6854: signal is true;
	signal I6859: std_logic; attribute dont_touch of I6859: signal is true;
	signal I6860: std_logic; attribute dont_touch of I6860: signal is true;
	signal I6861: std_logic; attribute dont_touch of I6861: signal is true;
	signal I6862: std_logic; attribute dont_touch of I6862: signal is true;
	signal I6863: std_logic; attribute dont_touch of I6863: signal is true;
	signal I6868: std_logic; attribute dont_touch of I6868: signal is true;
	signal I6869: std_logic; attribute dont_touch of I6869: signal is true;
	signal I6870: std_logic; attribute dont_touch of I6870: signal is true;
	signal I6875: std_logic; attribute dont_touch of I6875: signal is true;
	signal I6876: std_logic; attribute dont_touch of I6876: signal is true;
	signal I6877: std_logic; attribute dont_touch of I6877: signal is true;
	signal I6878: std_logic; attribute dont_touch of I6878: signal is true;
	signal I6883: std_logic; attribute dont_touch of I6883: signal is true;
	signal I6884: std_logic; attribute dont_touch of I6884: signal is true;
	signal I6885: std_logic; attribute dont_touch of I6885: signal is true;
	signal I6890: std_logic; attribute dont_touch of I6890: signal is true;
	signal I6891: std_logic; attribute dont_touch of I6891: signal is true;
	signal I6892: std_logic; attribute dont_touch of I6892: signal is true;
	signal I6893: std_logic; attribute dont_touch of I6893: signal is true;
	signal I6894: std_logic; attribute dont_touch of I6894: signal is true;
	signal I6899: std_logic; attribute dont_touch of I6899: signal is true;
	signal I6900: std_logic; attribute dont_touch of I6900: signal is true;
	signal I6901: std_logic; attribute dont_touch of I6901: signal is true;
	signal I6906: std_logic; attribute dont_touch of I6906: signal is true;
	signal I6907: std_logic; attribute dont_touch of I6907: signal is true;
	signal I6908: std_logic; attribute dont_touch of I6908: signal is true;
	signal I6909: std_logic; attribute dont_touch of I6909: signal is true;
	signal I6914: std_logic; attribute dont_touch of I6914: signal is true;
	signal I6915: std_logic; attribute dont_touch of I6915: signal is true;
	signal I6916: std_logic; attribute dont_touch of I6916: signal is true;
	signal I6921: std_logic; attribute dont_touch of I6921: signal is true;
	signal I6922: std_logic; attribute dont_touch of I6922: signal is true;
	signal I6923: std_logic; attribute dont_touch of I6923: signal is true;
	signal I6924: std_logic; attribute dont_touch of I6924: signal is true;
	signal I6925: std_logic; attribute dont_touch of I6925: signal is true;
	signal I6930: std_logic; attribute dont_touch of I6930: signal is true;
	signal I6931: std_logic; attribute dont_touch of I6931: signal is true;
	signal I6932: std_logic; attribute dont_touch of I6932: signal is true;
	signal I6937: std_logic; attribute dont_touch of I6937: signal is true;
	signal I6938: std_logic; attribute dont_touch of I6938: signal is true;
	signal I6939: std_logic; attribute dont_touch of I6939: signal is true;
	signal I6940: std_logic; attribute dont_touch of I6940: signal is true;
	signal I6945: std_logic; attribute dont_touch of I6945: signal is true;
	signal I6946: std_logic; attribute dont_touch of I6946: signal is true;
	signal I6947: std_logic; attribute dont_touch of I6947: signal is true;
	signal I6952: std_logic; attribute dont_touch of I6952: signal is true;
	signal I6953: std_logic; attribute dont_touch of I6953: signal is true;
	signal I6954: std_logic; attribute dont_touch of I6954: signal is true;
	signal I6955: std_logic; attribute dont_touch of I6955: signal is true;
	signal I6956: std_logic; attribute dont_touch of I6956: signal is true;
	signal I6961: std_logic; attribute dont_touch of I6961: signal is true;
	signal I6962: std_logic; attribute dont_touch of I6962: signal is true;
	signal I6963: std_logic; attribute dont_touch of I6963: signal is true;
	signal I6968: std_logic; attribute dont_touch of I6968: signal is true;
	signal I6969: std_logic; attribute dont_touch of I6969: signal is true;
	signal I6970: std_logic; attribute dont_touch of I6970: signal is true;
	signal I6971: std_logic; attribute dont_touch of I6971: signal is true;
	signal I6976: std_logic; attribute dont_touch of I6976: signal is true;
	signal I6977: std_logic; attribute dont_touch of I6977: signal is true;
	signal I6978: std_logic; attribute dont_touch of I6978: signal is true;
	signal I7057: std_logic; attribute dont_touch of I7057: signal is true;
	signal I7058: std_logic; attribute dont_touch of I7058: signal is true;
	signal I7059: std_logic; attribute dont_touch of I7059: signal is true;
	signal I7070: std_logic; attribute dont_touch of I7070: signal is true;
	signal I7071: std_logic; attribute dont_touch of I7071: signal is true;
	signal I7072: std_logic; attribute dont_touch of I7072: signal is true;
	signal I7083: std_logic; attribute dont_touch of I7083: signal is true;
	signal I7084: std_logic; attribute dont_touch of I7084: signal is true;
	signal I7085: std_logic; attribute dont_touch of I7085: signal is true;
	signal I7096: std_logic; attribute dont_touch of I7096: signal is true;
	signal I7097: std_logic; attribute dont_touch of I7097: signal is true;
	signal I7098: std_logic; attribute dont_touch of I7098: signal is true;
	signal I7109: std_logic; attribute dont_touch of I7109: signal is true;
	signal I7110: std_logic; attribute dont_touch of I7110: signal is true;
	signal I7111: std_logic; attribute dont_touch of I7111: signal is true;
	signal I7122: std_logic; attribute dont_touch of I7122: signal is true;
	signal I7123: std_logic; attribute dont_touch of I7123: signal is true;
	signal I7124: std_logic; attribute dont_touch of I7124: signal is true;
	signal I7135: std_logic; attribute dont_touch of I7135: signal is true;
	signal I7136: std_logic; attribute dont_touch of I7136: signal is true;
	signal I7137: std_logic; attribute dont_touch of I7137: signal is true;
	signal I7148: std_logic; attribute dont_touch of I7148: signal is true;
	signal I7149: std_logic; attribute dont_touch of I7149: signal is true;
	signal I7150: std_logic; attribute dont_touch of I7150: signal is true;
	signal I7161: std_logic; attribute dont_touch of I7161: signal is true;
	signal I7162: std_logic; attribute dont_touch of I7162: signal is true;
	signal I7163: std_logic; attribute dont_touch of I7163: signal is true;
	signal I7174: std_logic; attribute dont_touch of I7174: signal is true;
	signal I7175: std_logic; attribute dont_touch of I7175: signal is true;
	signal I7176: std_logic; attribute dont_touch of I7176: signal is true;
	signal I7187: std_logic; attribute dont_touch of I7187: signal is true;
	signal I7188: std_logic; attribute dont_touch of I7188: signal is true;
	signal I7189: std_logic; attribute dont_touch of I7189: signal is true;
	signal I7200: std_logic; attribute dont_touch of I7200: signal is true;
	signal I7201: std_logic; attribute dont_touch of I7201: signal is true;
	signal I7202: std_logic; attribute dont_touch of I7202: signal is true;
	signal I7213: std_logic; attribute dont_touch of I7213: signal is true;
	signal I7214: std_logic; attribute dont_touch of I7214: signal is true;
	signal I7215: std_logic; attribute dont_touch of I7215: signal is true;
	signal I7226: std_logic; attribute dont_touch of I7226: signal is true;
	signal I7227: std_logic; attribute dont_touch of I7227: signal is true;
	signal I7228: std_logic; attribute dont_touch of I7228: signal is true;
	signal I7239: std_logic; attribute dont_touch of I7239: signal is true;
	signal I7240: std_logic; attribute dont_touch of I7240: signal is true;
	signal I7241: std_logic; attribute dont_touch of I7241: signal is true;
	signal I7252: std_logic; attribute dont_touch of I7252: signal is true;
	signal I7253: std_logic; attribute dont_touch of I7253: signal is true;
	signal I7254: std_logic; attribute dont_touch of I7254: signal is true;
	signal I7265: std_logic; attribute dont_touch of I7265: signal is true;
	signal I7266: std_logic; attribute dont_touch of I7266: signal is true;
	signal I7267: std_logic; attribute dont_touch of I7267: signal is true;
	signal I7278: std_logic; attribute dont_touch of I7278: signal is true;
	signal I7279: std_logic; attribute dont_touch of I7279: signal is true;
	signal I7280: std_logic; attribute dont_touch of I7280: signal is true;
	signal I7291: std_logic; attribute dont_touch of I7291: signal is true;
	signal I7292: std_logic; attribute dont_touch of I7292: signal is true;
	signal I7293: std_logic; attribute dont_touch of I7293: signal is true;
	signal I7304: std_logic; attribute dont_touch of I7304: signal is true;
	signal I7305: std_logic; attribute dont_touch of I7305: signal is true;
	signal I7306: std_logic; attribute dont_touch of I7306: signal is true;
	signal I7317: std_logic; attribute dont_touch of I7317: signal is true;
	signal I7318: std_logic; attribute dont_touch of I7318: signal is true;
	signal I7319: std_logic; attribute dont_touch of I7319: signal is true;
	signal I7330: std_logic; attribute dont_touch of I7330: signal is true;
	signal I7331: std_logic; attribute dont_touch of I7331: signal is true;
	signal I7332: std_logic; attribute dont_touch of I7332: signal is true;
	signal I7343: std_logic; attribute dont_touch of I7343: signal is true;
	signal I7344: std_logic; attribute dont_touch of I7344: signal is true;
	signal I7345: std_logic; attribute dont_touch of I7345: signal is true;
	signal I7356: std_logic; attribute dont_touch of I7356: signal is true;
	signal I7357: std_logic; attribute dont_touch of I7357: signal is true;
	signal I7358: std_logic; attribute dont_touch of I7358: signal is true;
	signal I7369: std_logic; attribute dont_touch of I7369: signal is true;
	signal I7370: std_logic; attribute dont_touch of I7370: signal is true;
	signal I7371: std_logic; attribute dont_touch of I7371: signal is true;
	signal I7382: std_logic; attribute dont_touch of I7382: signal is true;
	signal I7383: std_logic; attribute dont_touch of I7383: signal is true;
	signal I7384: std_logic; attribute dont_touch of I7384: signal is true;
	signal I7395: std_logic; attribute dont_touch of I7395: signal is true;
	signal I7396: std_logic; attribute dont_touch of I7396: signal is true;
	signal I7397: std_logic; attribute dont_touch of I7397: signal is true;
	signal I7408: std_logic; attribute dont_touch of I7408: signal is true;
	signal I7409: std_logic; attribute dont_touch of I7409: signal is true;
	signal I7410: std_logic; attribute dont_touch of I7410: signal is true;
	signal I7421: std_logic; attribute dont_touch of I7421: signal is true;
	signal I7422: std_logic; attribute dont_touch of I7422: signal is true;
	signal I7423: std_logic; attribute dont_touch of I7423: signal is true;
	signal I7434: std_logic; attribute dont_touch of I7434: signal is true;
	signal I7435: std_logic; attribute dont_touch of I7435: signal is true;
	signal I7436: std_logic; attribute dont_touch of I7436: signal is true;
	signal I7447: std_logic; attribute dont_touch of I7447: signal is true;
	signal I7448: std_logic; attribute dont_touch of I7448: signal is true;
	signal I7449: std_logic; attribute dont_touch of I7449: signal is true;
	signal I7460: std_logic; attribute dont_touch of I7460: signal is true;
	signal I7461: std_logic; attribute dont_touch of I7461: signal is true;
	signal I7462: std_logic; attribute dont_touch of I7462: signal is true;
	signal I7474: std_logic; attribute dont_touch of I7474: signal is true;
	signal I7475: std_logic; attribute dont_touch of I7475: signal is true;
	signal I7476: std_logic; attribute dont_touch of I7476: signal is true;
	signal I7477: std_logic; attribute dont_touch of I7477: signal is true;
	signal I7482: std_logic; attribute dont_touch of I7482: signal is true;
	signal I7483: std_logic; attribute dont_touch of I7483: signal is true;
	signal I7484: std_logic; attribute dont_touch of I7484: signal is true;
	signal I7489: std_logic; attribute dont_touch of I7489: signal is true;
	signal I7490: std_logic; attribute dont_touch of I7490: signal is true;
	signal I7491: std_logic; attribute dont_touch of I7491: signal is true;
	signal I7492: std_logic; attribute dont_touch of I7492: signal is true;
	signal I7497: std_logic; attribute dont_touch of I7497: signal is true;
	signal I7498: std_logic; attribute dont_touch of I7498: signal is true;
	signal I7499: std_logic; attribute dont_touch of I7499: signal is true;
	signal I7504: std_logic; attribute dont_touch of I7504: signal is true;
	signal I7505: std_logic; attribute dont_touch of I7505: signal is true;
	signal I7506: std_logic; attribute dont_touch of I7506: signal is true;
	signal I7507: std_logic; attribute dont_touch of I7507: signal is true;
	signal I7512: std_logic; attribute dont_touch of I7512: signal is true;
	signal I7513: std_logic; attribute dont_touch of I7513: signal is true;
	signal I7514: std_logic; attribute dont_touch of I7514: signal is true;
	signal I7519: std_logic; attribute dont_touch of I7519: signal is true;
	signal I7520: std_logic; attribute dont_touch of I7520: signal is true;
	signal I7521: std_logic; attribute dont_touch of I7521: signal is true;
	signal I7526: std_logic; attribute dont_touch of I7526: signal is true;
	signal I7527: std_logic; attribute dont_touch of I7527: signal is true;
	signal I7528: std_logic; attribute dont_touch of I7528: signal is true;
	signal I7533: std_logic; attribute dont_touch of I7533: signal is true;
	signal I7534: std_logic; attribute dont_touch of I7534: signal is true;
	signal I7535: std_logic; attribute dont_touch of I7535: signal is true;
	signal I7540: std_logic; attribute dont_touch of I7540: signal is true;
	signal I7541: std_logic; attribute dont_touch of I7541: signal is true;
	signal I7542: std_logic; attribute dont_touch of I7542: signal is true;
	signal I7547: std_logic; attribute dont_touch of I7547: signal is true;
	signal I7548: std_logic; attribute dont_touch of I7548: signal is true;
	signal I7549: std_logic; attribute dont_touch of I7549: signal is true;
	signal I7554: std_logic; attribute dont_touch of I7554: signal is true;
	signal I7555: std_logic; attribute dont_touch of I7555: signal is true;
	signal I7556: std_logic; attribute dont_touch of I7556: signal is true;
	signal I7561: std_logic; attribute dont_touch of I7561: signal is true;
	signal I7562: std_logic; attribute dont_touch of I7562: signal is true;
	signal I7563: std_logic; attribute dont_touch of I7563: signal is true;
	signal I7568: std_logic; attribute dont_touch of I7568: signal is true;
	signal I7569: std_logic; attribute dont_touch of I7569: signal is true;
	signal I7570: std_logic; attribute dont_touch of I7570: signal is true;
	signal I7575: std_logic; attribute dont_touch of I7575: signal is true;
	signal I7576: std_logic; attribute dont_touch of I7576: signal is true;
	signal I7577: std_logic; attribute dont_touch of I7577: signal is true;
	signal I7582: std_logic; attribute dont_touch of I7582: signal is true;
	signal I7583: std_logic; attribute dont_touch of I7583: signal is true;
	signal I7584: std_logic; attribute dont_touch of I7584: signal is true;
	signal I7589: std_logic; attribute dont_touch of I7589: signal is true;
	signal I7590: std_logic; attribute dont_touch of I7590: signal is true;
	signal I7591: std_logic; attribute dont_touch of I7591: signal is true;
	signal I7596: std_logic; attribute dont_touch of I7596: signal is true;
	signal I7597: std_logic; attribute dont_touch of I7597: signal is true;
	signal I7598: std_logic; attribute dont_touch of I7598: signal is true;
	signal I7603: std_logic; attribute dont_touch of I7603: signal is true;
	signal I7604: std_logic; attribute dont_touch of I7604: signal is true;
	signal I7605: std_logic; attribute dont_touch of I7605: signal is true;
	signal I7610: std_logic; attribute dont_touch of I7610: signal is true;
	signal I7611: std_logic; attribute dont_touch of I7611: signal is true;
	signal I7612: std_logic; attribute dont_touch of I7612: signal is true;
	signal I7617: std_logic; attribute dont_touch of I7617: signal is true;
	signal I7618: std_logic; attribute dont_touch of I7618: signal is true;
	signal I7619: std_logic; attribute dont_touch of I7619: signal is true;
	signal I7624: std_logic; attribute dont_touch of I7624: signal is true;
	signal I7625: std_logic; attribute dont_touch of I7625: signal is true;
	signal I7626: std_logic; attribute dont_touch of I7626: signal is true;
	signal I7631: std_logic; attribute dont_touch of I7631: signal is true;
	signal I7632: std_logic; attribute dont_touch of I7632: signal is true;
	signal I7633: std_logic; attribute dont_touch of I7633: signal is true;
	signal I7638: std_logic; attribute dont_touch of I7638: signal is true;
	signal I7639: std_logic; attribute dont_touch of I7639: signal is true;
	signal I7640: std_logic; attribute dont_touch of I7640: signal is true;
	signal I7645: std_logic; attribute dont_touch of I7645: signal is true;
	signal I7646: std_logic; attribute dont_touch of I7646: signal is true;
	signal I7647: std_logic; attribute dont_touch of I7647: signal is true;
	signal I7652: std_logic; attribute dont_touch of I7652: signal is true;
	signal I7653: std_logic; attribute dont_touch of I7653: signal is true;
	signal I7654: std_logic; attribute dont_touch of I7654: signal is true;
	signal I7659: std_logic; attribute dont_touch of I7659: signal is true;
	signal I7660: std_logic; attribute dont_touch of I7660: signal is true;
	signal I7661: std_logic; attribute dont_touch of I7661: signal is true;
	signal I7666: std_logic; attribute dont_touch of I7666: signal is true;
	signal I7667: std_logic; attribute dont_touch of I7667: signal is true;
	signal I7668: std_logic; attribute dont_touch of I7668: signal is true;
	signal I7673: std_logic; attribute dont_touch of I7673: signal is true;
	signal I7674: std_logic; attribute dont_touch of I7674: signal is true;
	signal I7675: std_logic; attribute dont_touch of I7675: signal is true;
	signal I7680: std_logic; attribute dont_touch of I7680: signal is true;
	signal I7681: std_logic; attribute dont_touch of I7681: signal is true;
	signal I7682: std_logic; attribute dont_touch of I7682: signal is true;
	signal I7687: std_logic; attribute dont_touch of I7687: signal is true;
	signal I7688: std_logic; attribute dont_touch of I7688: signal is true;
	signal I7689: std_logic; attribute dont_touch of I7689: signal is true;
	signal I7694: std_logic; attribute dont_touch of I7694: signal is true;
	signal I7695: std_logic; attribute dont_touch of I7695: signal is true;
	signal I7696: std_logic; attribute dont_touch of I7696: signal is true;
	signal I7701: std_logic; attribute dont_touch of I7701: signal is true;
	signal I7702: std_logic; attribute dont_touch of I7702: signal is true;
	signal I7703: std_logic; attribute dont_touch of I7703: signal is true;
	signal I7708: std_logic; attribute dont_touch of I7708: signal is true;
	signal I7709: std_logic; attribute dont_touch of I7709: signal is true;
	signal I7710: std_logic; attribute dont_touch of I7710: signal is true;
	signal I7715: std_logic; attribute dont_touch of I7715: signal is true;
	signal I7716: std_logic; attribute dont_touch of I7716: signal is true;
	signal I7717: std_logic; attribute dont_touch of I7717: signal is true;
	signal I9996: std_logic; attribute dont_touch of I9996: signal is true;
	signal I9997: std_logic; attribute dont_touch of I9997: signal is true;
	signal I9998: std_logic; attribute dont_touch of I9998: signal is true;
	signal I9999: std_logic; attribute dont_touch of I9999: signal is true;
	signal I10000: std_logic; attribute dont_touch of I10000: signal is true;
	signal I10005: std_logic; attribute dont_touch of I10005: signal is true;
	signal I10006: std_logic; attribute dont_touch of I10006: signal is true;
	signal I10007: std_logic; attribute dont_touch of I10007: signal is true;
	signal I10012: std_logic; attribute dont_touch of I10012: signal is true;
	signal I10013: std_logic; attribute dont_touch of I10013: signal is true;
	signal I10014: std_logic; attribute dont_touch of I10014: signal is true;
	signal I10015: std_logic; attribute dont_touch of I10015: signal is true;
	signal I10020: std_logic; attribute dont_touch of I10020: signal is true;
	signal I10021: std_logic; attribute dont_touch of I10021: signal is true;
	signal I10022: std_logic; attribute dont_touch of I10022: signal is true;
	signal I10027: std_logic; attribute dont_touch of I10027: signal is true;
	signal I10028: std_logic; attribute dont_touch of I10028: signal is true;
	signal I10029: std_logic; attribute dont_touch of I10029: signal is true;
	signal I10030: std_logic; attribute dont_touch of I10030: signal is true;
	signal I10031: std_logic; attribute dont_touch of I10031: signal is true;
	signal I10036: std_logic; attribute dont_touch of I10036: signal is true;
	signal I10037: std_logic; attribute dont_touch of I10037: signal is true;
	signal I10038: std_logic; attribute dont_touch of I10038: signal is true;
	signal I10043: std_logic; attribute dont_touch of I10043: signal is true;
	signal I10044: std_logic; attribute dont_touch of I10044: signal is true;
	signal I10045: std_logic; attribute dont_touch of I10045: signal is true;
	signal I10046: std_logic; attribute dont_touch of I10046: signal is true;
	signal I10051: std_logic; attribute dont_touch of I10051: signal is true;
	signal I10052: std_logic; attribute dont_touch of I10052: signal is true;
	signal I10053: std_logic; attribute dont_touch of I10053: signal is true;
	signal I10058: std_logic; attribute dont_touch of I10058: signal is true;
	signal I10059: std_logic; attribute dont_touch of I10059: signal is true;
	signal I10060: std_logic; attribute dont_touch of I10060: signal is true;
	signal I10061: std_logic; attribute dont_touch of I10061: signal is true;
	signal I10062: std_logic; attribute dont_touch of I10062: signal is true;
	signal I10067: std_logic; attribute dont_touch of I10067: signal is true;
	signal I10068: std_logic; attribute dont_touch of I10068: signal is true;
	signal I10069: std_logic; attribute dont_touch of I10069: signal is true;
	signal I10074: std_logic; attribute dont_touch of I10074: signal is true;
	signal I10075: std_logic; attribute dont_touch of I10075: signal is true;
	signal I10076: std_logic; attribute dont_touch of I10076: signal is true;
	signal I10077: std_logic; attribute dont_touch of I10077: signal is true;
	signal I10082: std_logic; attribute dont_touch of I10082: signal is true;
	signal I10083: std_logic; attribute dont_touch of I10083: signal is true;
	signal I10084: std_logic; attribute dont_touch of I10084: signal is true;
	signal I10089: std_logic; attribute dont_touch of I10089: signal is true;
	signal I10090: std_logic; attribute dont_touch of I10090: signal is true;
	signal I10091: std_logic; attribute dont_touch of I10091: signal is true;
	signal I10092: std_logic; attribute dont_touch of I10092: signal is true;
	signal I10093: std_logic; attribute dont_touch of I10093: signal is true;
	signal I10098: std_logic; attribute dont_touch of I10098: signal is true;
	signal I10099: std_logic; attribute dont_touch of I10099: signal is true;
	signal I10100: std_logic; attribute dont_touch of I10100: signal is true;
	signal I10105: std_logic; attribute dont_touch of I10105: signal is true;
	signal I10106: std_logic; attribute dont_touch of I10106: signal is true;
	signal I10107: std_logic; attribute dont_touch of I10107: signal is true;
	signal I10108: std_logic; attribute dont_touch of I10108: signal is true;
	signal I10113: std_logic; attribute dont_touch of I10113: signal is true;
	signal I10114: std_logic; attribute dont_touch of I10114: signal is true;
	signal I10115: std_logic; attribute dont_touch of I10115: signal is true;
	signal I10120: std_logic; attribute dont_touch of I10120: signal is true;
	signal I10121: std_logic; attribute dont_touch of I10121: signal is true;
	signal I10122: std_logic; attribute dont_touch of I10122: signal is true;
	signal I10123: std_logic; attribute dont_touch of I10123: signal is true;
	signal I10124: std_logic; attribute dont_touch of I10124: signal is true;
	signal I10129: std_logic; attribute dont_touch of I10129: signal is true;
	signal I10130: std_logic; attribute dont_touch of I10130: signal is true;
	signal I10131: std_logic; attribute dont_touch of I10131: signal is true;
	signal I10136: std_logic; attribute dont_touch of I10136: signal is true;
	signal I10137: std_logic; attribute dont_touch of I10137: signal is true;
	signal I10138: std_logic; attribute dont_touch of I10138: signal is true;
	signal I10139: std_logic; attribute dont_touch of I10139: signal is true;
	signal I10144: std_logic; attribute dont_touch of I10144: signal is true;
	signal I10145: std_logic; attribute dont_touch of I10145: signal is true;
	signal I10146: std_logic; attribute dont_touch of I10146: signal is true;
	signal I10151: std_logic; attribute dont_touch of I10151: signal is true;
	signal I10152: std_logic; attribute dont_touch of I10152: signal is true;
	signal I10153: std_logic; attribute dont_touch of I10153: signal is true;
	signal I10154: std_logic; attribute dont_touch of I10154: signal is true;
	signal I10155: std_logic; attribute dont_touch of I10155: signal is true;
	signal I10160: std_logic; attribute dont_touch of I10160: signal is true;
	signal I10161: std_logic; attribute dont_touch of I10161: signal is true;
	signal I10162: std_logic; attribute dont_touch of I10162: signal is true;
	signal I10167: std_logic; attribute dont_touch of I10167: signal is true;
	signal I10168: std_logic; attribute dont_touch of I10168: signal is true;
	signal I10169: std_logic; attribute dont_touch of I10169: signal is true;
	signal I10170: std_logic; attribute dont_touch of I10170: signal is true;
	signal I10175: std_logic; attribute dont_touch of I10175: signal is true;
	signal I10176: std_logic; attribute dont_touch of I10176: signal is true;
	signal I10177: std_logic; attribute dont_touch of I10177: signal is true;
	signal I10182: std_logic; attribute dont_touch of I10182: signal is true;
	signal I10183: std_logic; attribute dont_touch of I10183: signal is true;
	signal I10184: std_logic; attribute dont_touch of I10184: signal is true;
	signal I10185: std_logic; attribute dont_touch of I10185: signal is true;
	signal I10186: std_logic; attribute dont_touch of I10186: signal is true;
	signal I10191: std_logic; attribute dont_touch of I10191: signal is true;
	signal I10192: std_logic; attribute dont_touch of I10192: signal is true;
	signal I10193: std_logic; attribute dont_touch of I10193: signal is true;
	signal I10198: std_logic; attribute dont_touch of I10198: signal is true;
	signal I10199: std_logic; attribute dont_touch of I10199: signal is true;
	signal I10200: std_logic; attribute dont_touch of I10200: signal is true;
	signal I10201: std_logic; attribute dont_touch of I10201: signal is true;
	signal I10206: std_logic; attribute dont_touch of I10206: signal is true;
	signal I10207: std_logic; attribute dont_touch of I10207: signal is true;
	signal I10208: std_logic; attribute dont_touch of I10208: signal is true;
	signal I10213: std_logic; attribute dont_touch of I10213: signal is true;
	signal I10214: std_logic; attribute dont_touch of I10214: signal is true;
	signal I10215: std_logic; attribute dont_touch of I10215: signal is true;
	signal I10216: std_logic; attribute dont_touch of I10216: signal is true;
	signal I10217: std_logic; attribute dont_touch of I10217: signal is true;
	signal I10222: std_logic; attribute dont_touch of I10222: signal is true;
	signal I10223: std_logic; attribute dont_touch of I10223: signal is true;
	signal I10224: std_logic; attribute dont_touch of I10224: signal is true;
	signal I10229: std_logic; attribute dont_touch of I10229: signal is true;
	signal I10230: std_logic; attribute dont_touch of I10230: signal is true;
	signal I10231: std_logic; attribute dont_touch of I10231: signal is true;
	signal I10232: std_logic; attribute dont_touch of I10232: signal is true;
	signal I10237: std_logic; attribute dont_touch of I10237: signal is true;
	signal I10238: std_logic; attribute dont_touch of I10238: signal is true;
	signal I10239: std_logic; attribute dont_touch of I10239: signal is true;
	signal I10244: std_logic; attribute dont_touch of I10244: signal is true;
	signal I10245: std_logic; attribute dont_touch of I10245: signal is true;
	signal I10246: std_logic; attribute dont_touch of I10246: signal is true;
	signal I10247: std_logic; attribute dont_touch of I10247: signal is true;
	signal I10248: std_logic; attribute dont_touch of I10248: signal is true;
	signal I10253: std_logic; attribute dont_touch of I10253: signal is true;
	signal I10254: std_logic; attribute dont_touch of I10254: signal is true;
	signal I10255: std_logic; attribute dont_touch of I10255: signal is true;
	signal I10260: std_logic; attribute dont_touch of I10260: signal is true;
	signal I10261: std_logic; attribute dont_touch of I10261: signal is true;
	signal I10262: std_logic; attribute dont_touch of I10262: signal is true;
	signal I10263: std_logic; attribute dont_touch of I10263: signal is true;
	signal I10268: std_logic; attribute dont_touch of I10268: signal is true;
	signal I10269: std_logic; attribute dont_touch of I10269: signal is true;
	signal I10270: std_logic; attribute dont_touch of I10270: signal is true;
	signal I10275: std_logic; attribute dont_touch of I10275: signal is true;
	signal I10276: std_logic; attribute dont_touch of I10276: signal is true;
	signal I10277: std_logic; attribute dont_touch of I10277: signal is true;
	signal I10278: std_logic; attribute dont_touch of I10278: signal is true;
	signal I10279: std_logic; attribute dont_touch of I10279: signal is true;
	signal I10284: std_logic; attribute dont_touch of I10284: signal is true;
	signal I10285: std_logic; attribute dont_touch of I10285: signal is true;
	signal I10286: std_logic; attribute dont_touch of I10286: signal is true;
	signal I10291: std_logic; attribute dont_touch of I10291: signal is true;
	signal I10292: std_logic; attribute dont_touch of I10292: signal is true;
	signal I10293: std_logic; attribute dont_touch of I10293: signal is true;
	signal I10294: std_logic; attribute dont_touch of I10294: signal is true;
	signal I10299: std_logic; attribute dont_touch of I10299: signal is true;
	signal I10300: std_logic; attribute dont_touch of I10300: signal is true;
	signal I10301: std_logic; attribute dont_touch of I10301: signal is true;
	signal I10306: std_logic; attribute dont_touch of I10306: signal is true;
	signal I10307: std_logic; attribute dont_touch of I10307: signal is true;
	signal I10308: std_logic; attribute dont_touch of I10308: signal is true;
	signal I10309: std_logic; attribute dont_touch of I10309: signal is true;
	signal I10310: std_logic; attribute dont_touch of I10310: signal is true;
	signal I10315: std_logic; attribute dont_touch of I10315: signal is true;
	signal I10316: std_logic; attribute dont_touch of I10316: signal is true;
	signal I10317: std_logic; attribute dont_touch of I10317: signal is true;
	signal I10322: std_logic; attribute dont_touch of I10322: signal is true;
	signal I10323: std_logic; attribute dont_touch of I10323: signal is true;
	signal I10324: std_logic; attribute dont_touch of I10324: signal is true;
	signal I10325: std_logic; attribute dont_touch of I10325: signal is true;
	signal I10330: std_logic; attribute dont_touch of I10330: signal is true;
	signal I10331: std_logic; attribute dont_touch of I10331: signal is true;
	signal I10332: std_logic; attribute dont_touch of I10332: signal is true;
	signal I10337: std_logic; attribute dont_touch of I10337: signal is true;
	signal I10338: std_logic; attribute dont_touch of I10338: signal is true;
	signal I10339: std_logic; attribute dont_touch of I10339: signal is true;
	signal I10340: std_logic; attribute dont_touch of I10340: signal is true;
	signal I10341: std_logic; attribute dont_touch of I10341: signal is true;
	signal I10346: std_logic; attribute dont_touch of I10346: signal is true;
	signal I10347: std_logic; attribute dont_touch of I10347: signal is true;
	signal I10348: std_logic; attribute dont_touch of I10348: signal is true;
	signal I10353: std_logic; attribute dont_touch of I10353: signal is true;
	signal I10354: std_logic; attribute dont_touch of I10354: signal is true;
	signal I10355: std_logic; attribute dont_touch of I10355: signal is true;
	signal I10356: std_logic; attribute dont_touch of I10356: signal is true;
	signal I10361: std_logic; attribute dont_touch of I10361: signal is true;
	signal I10362: std_logic; attribute dont_touch of I10362: signal is true;
	signal I10363: std_logic; attribute dont_touch of I10363: signal is true;
	signal I10368: std_logic; attribute dont_touch of I10368: signal is true;
	signal I10369: std_logic; attribute dont_touch of I10369: signal is true;
	signal I10370: std_logic; attribute dont_touch of I10370: signal is true;
	signal I10371: std_logic; attribute dont_touch of I10371: signal is true;
	signal I10372: std_logic; attribute dont_touch of I10372: signal is true;
	signal I10377: std_logic; attribute dont_touch of I10377: signal is true;
	signal I10378: std_logic; attribute dont_touch of I10378: signal is true;
	signal I10379: std_logic; attribute dont_touch of I10379: signal is true;
	signal I10384: std_logic; attribute dont_touch of I10384: signal is true;
	signal I10385: std_logic; attribute dont_touch of I10385: signal is true;
	signal I10386: std_logic; attribute dont_touch of I10386: signal is true;
	signal I10387: std_logic; attribute dont_touch of I10387: signal is true;
	signal I10392: std_logic; attribute dont_touch of I10392: signal is true;
	signal I10393: std_logic; attribute dont_touch of I10393: signal is true;
	signal I10394: std_logic; attribute dont_touch of I10394: signal is true;
	signal I10399: std_logic; attribute dont_touch of I10399: signal is true;
	signal I10400: std_logic; attribute dont_touch of I10400: signal is true;
	signal I10401: std_logic; attribute dont_touch of I10401: signal is true;
	signal I10402: std_logic; attribute dont_touch of I10402: signal is true;
	signal I10403: std_logic; attribute dont_touch of I10403: signal is true;
	signal I10408: std_logic; attribute dont_touch of I10408: signal is true;
	signal I10409: std_logic; attribute dont_touch of I10409: signal is true;
	signal I10410: std_logic; attribute dont_touch of I10410: signal is true;
	signal I10415: std_logic; attribute dont_touch of I10415: signal is true;
	signal I10416: std_logic; attribute dont_touch of I10416: signal is true;
	signal I10417: std_logic; attribute dont_touch of I10417: signal is true;
	signal I10418: std_logic; attribute dont_touch of I10418: signal is true;
	signal I10423: std_logic; attribute dont_touch of I10423: signal is true;
	signal I10424: std_logic; attribute dont_touch of I10424: signal is true;
	signal I10425: std_logic; attribute dont_touch of I10425: signal is true;
	signal I10430: std_logic; attribute dont_touch of I10430: signal is true;
	signal I10431: std_logic; attribute dont_touch of I10431: signal is true;
	signal I10432: std_logic; attribute dont_touch of I10432: signal is true;
	signal I10433: std_logic; attribute dont_touch of I10433: signal is true;
	signal I10434: std_logic; attribute dont_touch of I10434: signal is true;
	signal I10439: std_logic; attribute dont_touch of I10439: signal is true;
	signal I10440: std_logic; attribute dont_touch of I10440: signal is true;
	signal I10441: std_logic; attribute dont_touch of I10441: signal is true;
	signal I10446: std_logic; attribute dont_touch of I10446: signal is true;
	signal I10447: std_logic; attribute dont_touch of I10447: signal is true;
	signal I10448: std_logic; attribute dont_touch of I10448: signal is true;
	signal I10449: std_logic; attribute dont_touch of I10449: signal is true;
	signal I10454: std_logic; attribute dont_touch of I10454: signal is true;
	signal I10455: std_logic; attribute dont_touch of I10455: signal is true;
	signal I10456: std_logic; attribute dont_touch of I10456: signal is true;
	signal I10461: std_logic; attribute dont_touch of I10461: signal is true;
	signal I10462: std_logic; attribute dont_touch of I10462: signal is true;
	signal I10463: std_logic; attribute dont_touch of I10463: signal is true;
	signal I10464: std_logic; attribute dont_touch of I10464: signal is true;
	signal I10465: std_logic; attribute dont_touch of I10465: signal is true;
	signal I10470: std_logic; attribute dont_touch of I10470: signal is true;
	signal I10471: std_logic; attribute dont_touch of I10471: signal is true;
	signal I10472: std_logic; attribute dont_touch of I10472: signal is true;
	signal I10477: std_logic; attribute dont_touch of I10477: signal is true;
	signal I10478: std_logic; attribute dont_touch of I10478: signal is true;
	signal I10479: std_logic; attribute dont_touch of I10479: signal is true;
	signal I10480: std_logic; attribute dont_touch of I10480: signal is true;
	signal I10485: std_logic; attribute dont_touch of I10485: signal is true;
	signal I10486: std_logic; attribute dont_touch of I10486: signal is true;
	signal I10487: std_logic; attribute dont_touch of I10487: signal is true;
	signal I10492: std_logic; attribute dont_touch of I10492: signal is true;
	signal I10493: std_logic; attribute dont_touch of I10493: signal is true;
	signal I10494: std_logic; attribute dont_touch of I10494: signal is true;
	signal I10495: std_logic; attribute dont_touch of I10495: signal is true;
	signal I10496: std_logic; attribute dont_touch of I10496: signal is true;
	signal I10501: std_logic; attribute dont_touch of I10501: signal is true;
	signal I10502: std_logic; attribute dont_touch of I10502: signal is true;
	signal I10503: std_logic; attribute dont_touch of I10503: signal is true;
	signal I10508: std_logic; attribute dont_touch of I10508: signal is true;
	signal I10509: std_logic; attribute dont_touch of I10509: signal is true;
	signal I10510: std_logic; attribute dont_touch of I10510: signal is true;
	signal I10511: std_logic; attribute dont_touch of I10511: signal is true;
	signal I10516: std_logic; attribute dont_touch of I10516: signal is true;
	signal I10517: std_logic; attribute dont_touch of I10517: signal is true;
	signal I10518: std_logic; attribute dont_touch of I10518: signal is true;
	signal I10523: std_logic; attribute dont_touch of I10523: signal is true;
	signal I10524: std_logic; attribute dont_touch of I10524: signal is true;
	signal I10525: std_logic; attribute dont_touch of I10525: signal is true;
	signal I10526: std_logic; attribute dont_touch of I10526: signal is true;
	signal I10527: std_logic; attribute dont_touch of I10527: signal is true;
	signal I10532: std_logic; attribute dont_touch of I10532: signal is true;
	signal I10533: std_logic; attribute dont_touch of I10533: signal is true;
	signal I10534: std_logic; attribute dont_touch of I10534: signal is true;
	signal I10539: std_logic; attribute dont_touch of I10539: signal is true;
	signal I10540: std_logic; attribute dont_touch of I10540: signal is true;
	signal I10541: std_logic; attribute dont_touch of I10541: signal is true;
	signal I10542: std_logic; attribute dont_touch of I10542: signal is true;
	signal I10547: std_logic; attribute dont_touch of I10547: signal is true;
	signal I10548: std_logic; attribute dont_touch of I10548: signal is true;
	signal I10549: std_logic; attribute dont_touch of I10549: signal is true;
	signal I10554: std_logic; attribute dont_touch of I10554: signal is true;
	signal I10555: std_logic; attribute dont_touch of I10555: signal is true;
	signal I10556: std_logic; attribute dont_touch of I10556: signal is true;
	signal I10557: std_logic; attribute dont_touch of I10557: signal is true;
	signal I10558: std_logic; attribute dont_touch of I10558: signal is true;
	signal I10563: std_logic; attribute dont_touch of I10563: signal is true;
	signal I10564: std_logic; attribute dont_touch of I10564: signal is true;
	signal I10565: std_logic; attribute dont_touch of I10565: signal is true;
	signal I10570: std_logic; attribute dont_touch of I10570: signal is true;
	signal I10571: std_logic; attribute dont_touch of I10571: signal is true;
	signal I10572: std_logic; attribute dont_touch of I10572: signal is true;
	signal I10573: std_logic; attribute dont_touch of I10573: signal is true;
	signal I10578: std_logic; attribute dont_touch of I10578: signal is true;
	signal I10579: std_logic; attribute dont_touch of I10579: signal is true;
	signal I10580: std_logic; attribute dont_touch of I10580: signal is true;
	signal I10585: std_logic; attribute dont_touch of I10585: signal is true;
	signal I10586: std_logic; attribute dont_touch of I10586: signal is true;
	signal I10587: std_logic; attribute dont_touch of I10587: signal is true;
	signal I10588: std_logic; attribute dont_touch of I10588: signal is true;
	signal I10589: std_logic; attribute dont_touch of I10589: signal is true;
	signal I10594: std_logic; attribute dont_touch of I10594: signal is true;
	signal I10595: std_logic; attribute dont_touch of I10595: signal is true;
	signal I10596: std_logic; attribute dont_touch of I10596: signal is true;
	signal I10601: std_logic; attribute dont_touch of I10601: signal is true;
	signal I10602: std_logic; attribute dont_touch of I10602: signal is true;
	signal I10603: std_logic; attribute dont_touch of I10603: signal is true;
	signal I10604: std_logic; attribute dont_touch of I10604: signal is true;
	signal I10609: std_logic; attribute dont_touch of I10609: signal is true;
	signal I10610: std_logic; attribute dont_touch of I10610: signal is true;
	signal I10611: std_logic; attribute dont_touch of I10611: signal is true;
	signal I10616: std_logic; attribute dont_touch of I10616: signal is true;
	signal I10617: std_logic; attribute dont_touch of I10617: signal is true;
	signal I10618: std_logic; attribute dont_touch of I10618: signal is true;
	signal I10619: std_logic; attribute dont_touch of I10619: signal is true;
	signal I10620: std_logic; attribute dont_touch of I10620: signal is true;
	signal I10625: std_logic; attribute dont_touch of I10625: signal is true;
	signal I10626: std_logic; attribute dont_touch of I10626: signal is true;
	signal I10627: std_logic; attribute dont_touch of I10627: signal is true;
	signal I10632: std_logic; attribute dont_touch of I10632: signal is true;
	signal I10633: std_logic; attribute dont_touch of I10633: signal is true;
	signal I10634: std_logic; attribute dont_touch of I10634: signal is true;
	signal I10635: std_logic; attribute dont_touch of I10635: signal is true;
	signal I10640: std_logic; attribute dont_touch of I10640: signal is true;
	signal I10641: std_logic; attribute dont_touch of I10641: signal is true;
	signal I10642: std_logic; attribute dont_touch of I10642: signal is true;
	signal I10647: std_logic; attribute dont_touch of I10647: signal is true;
	signal I10648: std_logic; attribute dont_touch of I10648: signal is true;
	signal I10649: std_logic; attribute dont_touch of I10649: signal is true;
	signal I10650: std_logic; attribute dont_touch of I10650: signal is true;
	signal I10651: std_logic; attribute dont_touch of I10651: signal is true;
	signal I10656: std_logic; attribute dont_touch of I10656: signal is true;
	signal I10657: std_logic; attribute dont_touch of I10657: signal is true;
	signal I10658: std_logic; attribute dont_touch of I10658: signal is true;
	signal I10663: std_logic; attribute dont_touch of I10663: signal is true;
	signal I10664: std_logic; attribute dont_touch of I10664: signal is true;
	signal I10665: std_logic; attribute dont_touch of I10665: signal is true;
	signal I10666: std_logic; attribute dont_touch of I10666: signal is true;
	signal I10671: std_logic; attribute dont_touch of I10671: signal is true;
	signal I10672: std_logic; attribute dont_touch of I10672: signal is true;
	signal I10673: std_logic; attribute dont_touch of I10673: signal is true;
	signal I10678: std_logic; attribute dont_touch of I10678: signal is true;
	signal I10679: std_logic; attribute dont_touch of I10679: signal is true;
	signal I10680: std_logic; attribute dont_touch of I10680: signal is true;
	signal I10681: std_logic; attribute dont_touch of I10681: signal is true;
	signal I10682: std_logic; attribute dont_touch of I10682: signal is true;
	signal I10687: std_logic; attribute dont_touch of I10687: signal is true;
	signal I10688: std_logic; attribute dont_touch of I10688: signal is true;
	signal I10689: std_logic; attribute dont_touch of I10689: signal is true;
	signal I10694: std_logic; attribute dont_touch of I10694: signal is true;
	signal I10695: std_logic; attribute dont_touch of I10695: signal is true;
	signal I10696: std_logic; attribute dont_touch of I10696: signal is true;
	signal I10697: std_logic; attribute dont_touch of I10697: signal is true;
	signal I10702: std_logic; attribute dont_touch of I10702: signal is true;
	signal I10703: std_logic; attribute dont_touch of I10703: signal is true;
	signal I10704: std_logic; attribute dont_touch of I10704: signal is true;
	signal I10709: std_logic; attribute dont_touch of I10709: signal is true;
	signal I10710: std_logic; attribute dont_touch of I10710: signal is true;
	signal I10711: std_logic; attribute dont_touch of I10711: signal is true;
	signal I10712: std_logic; attribute dont_touch of I10712: signal is true;
	signal I10713: std_logic; attribute dont_touch of I10713: signal is true;
	signal I10718: std_logic; attribute dont_touch of I10718: signal is true;
	signal I10719: std_logic; attribute dont_touch of I10719: signal is true;
	signal I10720: std_logic; attribute dont_touch of I10720: signal is true;
	signal I10725: std_logic; attribute dont_touch of I10725: signal is true;
	signal I10726: std_logic; attribute dont_touch of I10726: signal is true;
	signal I10727: std_logic; attribute dont_touch of I10727: signal is true;
	signal I10728: std_logic; attribute dont_touch of I10728: signal is true;
	signal I10733: std_logic; attribute dont_touch of I10733: signal is true;
	signal I10734: std_logic; attribute dont_touch of I10734: signal is true;
	signal I10735: std_logic; attribute dont_touch of I10735: signal is true;
	signal I10740: std_logic; attribute dont_touch of I10740: signal is true;
	signal I10741: std_logic; attribute dont_touch of I10741: signal is true;
	signal I10742: std_logic; attribute dont_touch of I10742: signal is true;
	signal I10743: std_logic; attribute dont_touch of I10743: signal is true;
	signal I10744: std_logic; attribute dont_touch of I10744: signal is true;
	signal I10749: std_logic; attribute dont_touch of I10749: signal is true;
	signal I10750: std_logic; attribute dont_touch of I10750: signal is true;
	signal I10751: std_logic; attribute dont_touch of I10751: signal is true;
	signal I10756: std_logic; attribute dont_touch of I10756: signal is true;
	signal I10757: std_logic; attribute dont_touch of I10757: signal is true;
	signal I10758: std_logic; attribute dont_touch of I10758: signal is true;
	signal I10759: std_logic; attribute dont_touch of I10759: signal is true;
	signal I10764: std_logic; attribute dont_touch of I10764: signal is true;
	signal I10765: std_logic; attribute dont_touch of I10765: signal is true;
	signal I10766: std_logic; attribute dont_touch of I10766: signal is true;
	signal I10771: std_logic; attribute dont_touch of I10771: signal is true;
	signal I10772: std_logic; attribute dont_touch of I10772: signal is true;
	signal I10773: std_logic; attribute dont_touch of I10773: signal is true;
	signal I10774: std_logic; attribute dont_touch of I10774: signal is true;
	signal I10775: std_logic; attribute dont_touch of I10775: signal is true;
	signal I10780: std_logic; attribute dont_touch of I10780: signal is true;
	signal I10781: std_logic; attribute dont_touch of I10781: signal is true;
	signal I10782: std_logic; attribute dont_touch of I10782: signal is true;
	signal I10787: std_logic; attribute dont_touch of I10787: signal is true;
	signal I10788: std_logic; attribute dont_touch of I10788: signal is true;
	signal I10789: std_logic; attribute dont_touch of I10789: signal is true;
	signal I10790: std_logic; attribute dont_touch of I10790: signal is true;
	signal I10795: std_logic; attribute dont_touch of I10795: signal is true;
	signal I10796: std_logic; attribute dont_touch of I10796: signal is true;
	signal I10797: std_logic; attribute dont_touch of I10797: signal is true;
	signal I10802: std_logic; attribute dont_touch of I10802: signal is true;
	signal I10803: std_logic; attribute dont_touch of I10803: signal is true;
	signal I10804: std_logic; attribute dont_touch of I10804: signal is true;
	signal I10805: std_logic; attribute dont_touch of I10805: signal is true;
	signal I10806: std_logic; attribute dont_touch of I10806: signal is true;
	signal I10811: std_logic; attribute dont_touch of I10811: signal is true;
	signal I10812: std_logic; attribute dont_touch of I10812: signal is true;
	signal I10813: std_logic; attribute dont_touch of I10813: signal is true;
	signal I10818: std_logic; attribute dont_touch of I10818: signal is true;
	signal I10819: std_logic; attribute dont_touch of I10819: signal is true;
	signal I10820: std_logic; attribute dont_touch of I10820: signal is true;
	signal I10821: std_logic; attribute dont_touch of I10821: signal is true;
	signal I10826: std_logic; attribute dont_touch of I10826: signal is true;
	signal I10827: std_logic; attribute dont_touch of I10827: signal is true;
	signal I10828: std_logic; attribute dont_touch of I10828: signal is true;
	signal I10833: std_logic; attribute dont_touch of I10833: signal is true;
	signal I10834: std_logic; attribute dont_touch of I10834: signal is true;
	signal I10835: std_logic; attribute dont_touch of I10835: signal is true;
	signal I10836: std_logic; attribute dont_touch of I10836: signal is true;
	signal I10837: std_logic; attribute dont_touch of I10837: signal is true;
	signal I10842: std_logic; attribute dont_touch of I10842: signal is true;
	signal I10843: std_logic; attribute dont_touch of I10843: signal is true;
	signal I10844: std_logic; attribute dont_touch of I10844: signal is true;
	signal I10849: std_logic; attribute dont_touch of I10849: signal is true;
	signal I10850: std_logic; attribute dont_touch of I10850: signal is true;
	signal I10851: std_logic; attribute dont_touch of I10851: signal is true;
	signal I10852: std_logic; attribute dont_touch of I10852: signal is true;
	signal I10857: std_logic; attribute dont_touch of I10857: signal is true;
	signal I10858: std_logic; attribute dont_touch of I10858: signal is true;
	signal I10859: std_logic; attribute dont_touch of I10859: signal is true;
	signal I10864: std_logic; attribute dont_touch of I10864: signal is true;
	signal I10865: std_logic; attribute dont_touch of I10865: signal is true;
	signal I10866: std_logic; attribute dont_touch of I10866: signal is true;
	signal I10867: std_logic; attribute dont_touch of I10867: signal is true;
	signal I10868: std_logic; attribute dont_touch of I10868: signal is true;
	signal I10873: std_logic; attribute dont_touch of I10873: signal is true;
	signal I10874: std_logic; attribute dont_touch of I10874: signal is true;
	signal I10875: std_logic; attribute dont_touch of I10875: signal is true;
	signal I10880: std_logic; attribute dont_touch of I10880: signal is true;
	signal I10881: std_logic; attribute dont_touch of I10881: signal is true;
	signal I10882: std_logic; attribute dont_touch of I10882: signal is true;
	signal I10883: std_logic; attribute dont_touch of I10883: signal is true;
	signal I10888: std_logic; attribute dont_touch of I10888: signal is true;
	signal I10889: std_logic; attribute dont_touch of I10889: signal is true;
	signal I10890: std_logic; attribute dont_touch of I10890: signal is true;
	signal I10895: std_logic; attribute dont_touch of I10895: signal is true;
	signal I10896: std_logic; attribute dont_touch of I10896: signal is true;
	signal I10897: std_logic; attribute dont_touch of I10897: signal is true;
	signal I10898: std_logic; attribute dont_touch of I10898: signal is true;
	signal I10899: std_logic; attribute dont_touch of I10899: signal is true;
	signal I10904: std_logic; attribute dont_touch of I10904: signal is true;
	signal I10905: std_logic; attribute dont_touch of I10905: signal is true;
	signal I10906: std_logic; attribute dont_touch of I10906: signal is true;
	signal I10911: std_logic; attribute dont_touch of I10911: signal is true;
	signal I10912: std_logic; attribute dont_touch of I10912: signal is true;
	signal I10913: std_logic; attribute dont_touch of I10913: signal is true;
	signal I10914: std_logic; attribute dont_touch of I10914: signal is true;
	signal I10919: std_logic; attribute dont_touch of I10919: signal is true;
	signal I10920: std_logic; attribute dont_touch of I10920: signal is true;
	signal I10921: std_logic; attribute dont_touch of I10921: signal is true;
	signal I10926: std_logic; attribute dont_touch of I10926: signal is true;
	signal I10927: std_logic; attribute dont_touch of I10927: signal is true;
	signal I10928: std_logic; attribute dont_touch of I10928: signal is true;
	signal I10929: std_logic; attribute dont_touch of I10929: signal is true;
	signal I10930: std_logic; attribute dont_touch of I10930: signal is true;
	signal I10935: std_logic; attribute dont_touch of I10935: signal is true;
	signal I10936: std_logic; attribute dont_touch of I10936: signal is true;
	signal I10937: std_logic; attribute dont_touch of I10937: signal is true;
	signal I10942: std_logic; attribute dont_touch of I10942: signal is true;
	signal I10943: std_logic; attribute dont_touch of I10943: signal is true;
	signal I10944: std_logic; attribute dont_touch of I10944: signal is true;
	signal I10945: std_logic; attribute dont_touch of I10945: signal is true;
	signal I10950: std_logic; attribute dont_touch of I10950: signal is true;
	signal I10951: std_logic; attribute dont_touch of I10951: signal is true;
	signal I10952: std_logic; attribute dont_touch of I10952: signal is true;
	signal I10957: std_logic; attribute dont_touch of I10957: signal is true;
	signal I10958: std_logic; attribute dont_touch of I10958: signal is true;
	signal I10959: std_logic; attribute dont_touch of I10959: signal is true;
	signal I10960: std_logic; attribute dont_touch of I10960: signal is true;
	signal I10961: std_logic; attribute dont_touch of I10961: signal is true;
	signal I10966: std_logic; attribute dont_touch of I10966: signal is true;
	signal I10967: std_logic; attribute dont_touch of I10967: signal is true;
	signal I10968: std_logic; attribute dont_touch of I10968: signal is true;
	signal I10973: std_logic; attribute dont_touch of I10973: signal is true;
	signal I10974: std_logic; attribute dont_touch of I10974: signal is true;
	signal I10975: std_logic; attribute dont_touch of I10975: signal is true;
	signal I10976: std_logic; attribute dont_touch of I10976: signal is true;
	signal I10981: std_logic; attribute dont_touch of I10981: signal is true;
	signal I10982: std_logic; attribute dont_touch of I10982: signal is true;
	signal I10983: std_logic; attribute dont_touch of I10983: signal is true;
	signal I11062: std_logic; attribute dont_touch of I11062: signal is true;
	signal I11063: std_logic; attribute dont_touch of I11063: signal is true;
	signal I11064: std_logic; attribute dont_touch of I11064: signal is true;
	signal I11075: std_logic; attribute dont_touch of I11075: signal is true;
	signal I11076: std_logic; attribute dont_touch of I11076: signal is true;
	signal I11077: std_logic; attribute dont_touch of I11077: signal is true;
	signal I11088: std_logic; attribute dont_touch of I11088: signal is true;
	signal I11089: std_logic; attribute dont_touch of I11089: signal is true;
	signal I11090: std_logic; attribute dont_touch of I11090: signal is true;
	signal I11101: std_logic; attribute dont_touch of I11101: signal is true;
	signal I11102: std_logic; attribute dont_touch of I11102: signal is true;
	signal I11103: std_logic; attribute dont_touch of I11103: signal is true;
	signal I11114: std_logic; attribute dont_touch of I11114: signal is true;
	signal I11115: std_logic; attribute dont_touch of I11115: signal is true;
	signal I11116: std_logic; attribute dont_touch of I11116: signal is true;
	signal I11127: std_logic; attribute dont_touch of I11127: signal is true;
	signal I11128: std_logic; attribute dont_touch of I11128: signal is true;
	signal I11129: std_logic; attribute dont_touch of I11129: signal is true;
	signal I11140: std_logic; attribute dont_touch of I11140: signal is true;
	signal I11141: std_logic; attribute dont_touch of I11141: signal is true;
	signal I11142: std_logic; attribute dont_touch of I11142: signal is true;
	signal I11153: std_logic; attribute dont_touch of I11153: signal is true;
	signal I11154: std_logic; attribute dont_touch of I11154: signal is true;
	signal I11155: std_logic; attribute dont_touch of I11155: signal is true;
	signal I11166: std_logic; attribute dont_touch of I11166: signal is true;
	signal I11167: std_logic; attribute dont_touch of I11167: signal is true;
	signal I11168: std_logic; attribute dont_touch of I11168: signal is true;
	signal I11179: std_logic; attribute dont_touch of I11179: signal is true;
	signal I11180: std_logic; attribute dont_touch of I11180: signal is true;
	signal I11181: std_logic; attribute dont_touch of I11181: signal is true;
	signal I11192: std_logic; attribute dont_touch of I11192: signal is true;
	signal I11193: std_logic; attribute dont_touch of I11193: signal is true;
	signal I11194: std_logic; attribute dont_touch of I11194: signal is true;
	signal I11205: std_logic; attribute dont_touch of I11205: signal is true;
	signal I11206: std_logic; attribute dont_touch of I11206: signal is true;
	signal I11207: std_logic; attribute dont_touch of I11207: signal is true;
	signal I11218: std_logic; attribute dont_touch of I11218: signal is true;
	signal I11219: std_logic; attribute dont_touch of I11219: signal is true;
	signal I11220: std_logic; attribute dont_touch of I11220: signal is true;
	signal I11231: std_logic; attribute dont_touch of I11231: signal is true;
	signal I11232: std_logic; attribute dont_touch of I11232: signal is true;
	signal I11233: std_logic; attribute dont_touch of I11233: signal is true;
	signal I11244: std_logic; attribute dont_touch of I11244: signal is true;
	signal I11245: std_logic; attribute dont_touch of I11245: signal is true;
	signal I11246: std_logic; attribute dont_touch of I11246: signal is true;
	signal I11257: std_logic; attribute dont_touch of I11257: signal is true;
	signal I11258: std_logic; attribute dont_touch of I11258: signal is true;
	signal I11259: std_logic; attribute dont_touch of I11259: signal is true;
	signal I11270: std_logic; attribute dont_touch of I11270: signal is true;
	signal I11271: std_logic; attribute dont_touch of I11271: signal is true;
	signal I11272: std_logic; attribute dont_touch of I11272: signal is true;
	signal I11283: std_logic; attribute dont_touch of I11283: signal is true;
	signal I11284: std_logic; attribute dont_touch of I11284: signal is true;
	signal I11285: std_logic; attribute dont_touch of I11285: signal is true;
	signal I11296: std_logic; attribute dont_touch of I11296: signal is true;
	signal I11297: std_logic; attribute dont_touch of I11297: signal is true;
	signal I11298: std_logic; attribute dont_touch of I11298: signal is true;
	signal I11309: std_logic; attribute dont_touch of I11309: signal is true;
	signal I11310: std_logic; attribute dont_touch of I11310: signal is true;
	signal I11311: std_logic; attribute dont_touch of I11311: signal is true;
	signal I11322: std_logic; attribute dont_touch of I11322: signal is true;
	signal I11323: std_logic; attribute dont_touch of I11323: signal is true;
	signal I11324: std_logic; attribute dont_touch of I11324: signal is true;
	signal I11335: std_logic; attribute dont_touch of I11335: signal is true;
	signal I11336: std_logic; attribute dont_touch of I11336: signal is true;
	signal I11337: std_logic; attribute dont_touch of I11337: signal is true;
	signal I11348: std_logic; attribute dont_touch of I11348: signal is true;
	signal I11349: std_logic; attribute dont_touch of I11349: signal is true;
	signal I11350: std_logic; attribute dont_touch of I11350: signal is true;
	signal I11361: std_logic; attribute dont_touch of I11361: signal is true;
	signal I11362: std_logic; attribute dont_touch of I11362: signal is true;
	signal I11363: std_logic; attribute dont_touch of I11363: signal is true;
	signal I11374: std_logic; attribute dont_touch of I11374: signal is true;
	signal I11375: std_logic; attribute dont_touch of I11375: signal is true;
	signal I11376: std_logic; attribute dont_touch of I11376: signal is true;
	signal I11387: std_logic; attribute dont_touch of I11387: signal is true;
	signal I11388: std_logic; attribute dont_touch of I11388: signal is true;
	signal I11389: std_logic; attribute dont_touch of I11389: signal is true;
	signal I11400: std_logic; attribute dont_touch of I11400: signal is true;
	signal I11401: std_logic; attribute dont_touch of I11401: signal is true;
	signal I11402: std_logic; attribute dont_touch of I11402: signal is true;
	signal I11413: std_logic; attribute dont_touch of I11413: signal is true;
	signal I11414: std_logic; attribute dont_touch of I11414: signal is true;
	signal I11415: std_logic; attribute dont_touch of I11415: signal is true;
	signal I11426: std_logic; attribute dont_touch of I11426: signal is true;
	signal I11427: std_logic; attribute dont_touch of I11427: signal is true;
	signal I11428: std_logic; attribute dont_touch of I11428: signal is true;
	signal I11439: std_logic; attribute dont_touch of I11439: signal is true;
	signal I11440: std_logic; attribute dont_touch of I11440: signal is true;
	signal I11441: std_logic; attribute dont_touch of I11441: signal is true;
	signal I11452: std_logic; attribute dont_touch of I11452: signal is true;
	signal I11453: std_logic; attribute dont_touch of I11453: signal is true;
	signal I11454: std_logic; attribute dont_touch of I11454: signal is true;
	signal I11465: std_logic; attribute dont_touch of I11465: signal is true;
	signal I11466: std_logic; attribute dont_touch of I11466: signal is true;
	signal I11467: std_logic; attribute dont_touch of I11467: signal is true;
	signal I11479: std_logic; attribute dont_touch of I11479: signal is true;
	signal I11480: std_logic; attribute dont_touch of I11480: signal is true;
	signal I11481: std_logic; attribute dont_touch of I11481: signal is true;
	signal I11482: std_logic; attribute dont_touch of I11482: signal is true;
	signal I11487: std_logic; attribute dont_touch of I11487: signal is true;
	signal I11488: std_logic; attribute dont_touch of I11488: signal is true;
	signal I11489: std_logic; attribute dont_touch of I11489: signal is true;
	signal I11494: std_logic; attribute dont_touch of I11494: signal is true;
	signal I11495: std_logic; attribute dont_touch of I11495: signal is true;
	signal I11496: std_logic; attribute dont_touch of I11496: signal is true;
	signal I11497: std_logic; attribute dont_touch of I11497: signal is true;
	signal I11502: std_logic; attribute dont_touch of I11502: signal is true;
	signal I11503: std_logic; attribute dont_touch of I11503: signal is true;
	signal I11504: std_logic; attribute dont_touch of I11504: signal is true;
	signal I11509: std_logic; attribute dont_touch of I11509: signal is true;
	signal I11510: std_logic; attribute dont_touch of I11510: signal is true;
	signal I11511: std_logic; attribute dont_touch of I11511: signal is true;
	signal I11512: std_logic; attribute dont_touch of I11512: signal is true;
	signal I11517: std_logic; attribute dont_touch of I11517: signal is true;
	signal I11518: std_logic; attribute dont_touch of I11518: signal is true;
	signal I11519: std_logic; attribute dont_touch of I11519: signal is true;
	signal I11524: std_logic; attribute dont_touch of I11524: signal is true;
	signal I11525: std_logic; attribute dont_touch of I11525: signal is true;
	signal I11526: std_logic; attribute dont_touch of I11526: signal is true;
	signal I11531: std_logic; attribute dont_touch of I11531: signal is true;
	signal I11532: std_logic; attribute dont_touch of I11532: signal is true;
	signal I11533: std_logic; attribute dont_touch of I11533: signal is true;
	signal I11538: std_logic; attribute dont_touch of I11538: signal is true;
	signal I11539: std_logic; attribute dont_touch of I11539: signal is true;
	signal I11540: std_logic; attribute dont_touch of I11540: signal is true;
	signal I11545: std_logic; attribute dont_touch of I11545: signal is true;
	signal I11546: std_logic; attribute dont_touch of I11546: signal is true;
	signal I11547: std_logic; attribute dont_touch of I11547: signal is true;
	signal I11552: std_logic; attribute dont_touch of I11552: signal is true;
	signal I11553: std_logic; attribute dont_touch of I11553: signal is true;
	signal I11554: std_logic; attribute dont_touch of I11554: signal is true;
	signal I11559: std_logic; attribute dont_touch of I11559: signal is true;
	signal I11560: std_logic; attribute dont_touch of I11560: signal is true;
	signal I11561: std_logic; attribute dont_touch of I11561: signal is true;
	signal I11566: std_logic; attribute dont_touch of I11566: signal is true;
	signal I11567: std_logic; attribute dont_touch of I11567: signal is true;
	signal I11568: std_logic; attribute dont_touch of I11568: signal is true;
	signal I11573: std_logic; attribute dont_touch of I11573: signal is true;
	signal I11574: std_logic; attribute dont_touch of I11574: signal is true;
	signal I11575: std_logic; attribute dont_touch of I11575: signal is true;
	signal I11580: std_logic; attribute dont_touch of I11580: signal is true;
	signal I11581: std_logic; attribute dont_touch of I11581: signal is true;
	signal I11582: std_logic; attribute dont_touch of I11582: signal is true;
	signal I11587: std_logic; attribute dont_touch of I11587: signal is true;
	signal I11588: std_logic; attribute dont_touch of I11588: signal is true;
	signal I11589: std_logic; attribute dont_touch of I11589: signal is true;
	signal I11594: std_logic; attribute dont_touch of I11594: signal is true;
	signal I11595: std_logic; attribute dont_touch of I11595: signal is true;
	signal I11596: std_logic; attribute dont_touch of I11596: signal is true;
	signal I11601: std_logic; attribute dont_touch of I11601: signal is true;
	signal I11602: std_logic; attribute dont_touch of I11602: signal is true;
	signal I11603: std_logic; attribute dont_touch of I11603: signal is true;
	signal I11608: std_logic; attribute dont_touch of I11608: signal is true;
	signal I11609: std_logic; attribute dont_touch of I11609: signal is true;
	signal I11610: std_logic; attribute dont_touch of I11610: signal is true;
	signal I11615: std_logic; attribute dont_touch of I11615: signal is true;
	signal I11616: std_logic; attribute dont_touch of I11616: signal is true;
	signal I11617: std_logic; attribute dont_touch of I11617: signal is true;
	signal I11622: std_logic; attribute dont_touch of I11622: signal is true;
	signal I11623: std_logic; attribute dont_touch of I11623: signal is true;
	signal I11624: std_logic; attribute dont_touch of I11624: signal is true;
	signal I11629: std_logic; attribute dont_touch of I11629: signal is true;
	signal I11630: std_logic; attribute dont_touch of I11630: signal is true;
	signal I11631: std_logic; attribute dont_touch of I11631: signal is true;
	signal I11636: std_logic; attribute dont_touch of I11636: signal is true;
	signal I11637: std_logic; attribute dont_touch of I11637: signal is true;
	signal I11638: std_logic; attribute dont_touch of I11638: signal is true;
	signal I11643: std_logic; attribute dont_touch of I11643: signal is true;
	signal I11644: std_logic; attribute dont_touch of I11644: signal is true;
	signal I11645: std_logic; attribute dont_touch of I11645: signal is true;
	signal I11650: std_logic; attribute dont_touch of I11650: signal is true;
	signal I11651: std_logic; attribute dont_touch of I11651: signal is true;
	signal I11652: std_logic; attribute dont_touch of I11652: signal is true;
	signal I11657: std_logic; attribute dont_touch of I11657: signal is true;
	signal I11658: std_logic; attribute dont_touch of I11658: signal is true;
	signal I11659: std_logic; attribute dont_touch of I11659: signal is true;
	signal I11664: std_logic; attribute dont_touch of I11664: signal is true;
	signal I11665: std_logic; attribute dont_touch of I11665: signal is true;
	signal I11666: std_logic; attribute dont_touch of I11666: signal is true;
	signal I11671: std_logic; attribute dont_touch of I11671: signal is true;
	signal I11672: std_logic; attribute dont_touch of I11672: signal is true;
	signal I11673: std_logic; attribute dont_touch of I11673: signal is true;
	signal I11678: std_logic; attribute dont_touch of I11678: signal is true;
	signal I11679: std_logic; attribute dont_touch of I11679: signal is true;
	signal I11680: std_logic; attribute dont_touch of I11680: signal is true;
	signal I11685: std_logic; attribute dont_touch of I11685: signal is true;
	signal I11686: std_logic; attribute dont_touch of I11686: signal is true;
	signal I11687: std_logic; attribute dont_touch of I11687: signal is true;
	signal I11692: std_logic; attribute dont_touch of I11692: signal is true;
	signal I11693: std_logic; attribute dont_touch of I11693: signal is true;
	signal I11694: std_logic; attribute dont_touch of I11694: signal is true;
	signal I11699: std_logic; attribute dont_touch of I11699: signal is true;
	signal I11700: std_logic; attribute dont_touch of I11700: signal is true;
	signal I11701: std_logic; attribute dont_touch of I11701: signal is true;
	signal I11706: std_logic; attribute dont_touch of I11706: signal is true;
	signal I11707: std_logic; attribute dont_touch of I11707: signal is true;
	signal I11708: std_logic; attribute dont_touch of I11708: signal is true;
	signal I11713: std_logic; attribute dont_touch of I11713: signal is true;
	signal I11714: std_logic; attribute dont_touch of I11714: signal is true;
	signal I11715: std_logic; attribute dont_touch of I11715: signal is true;
	signal I11720: std_logic; attribute dont_touch of I11720: signal is true;
	signal I11721: std_logic; attribute dont_touch of I11721: signal is true;
	signal I11722: std_logic; attribute dont_touch of I11722: signal is true;
	signal I14001: std_logic; attribute dont_touch of I14001: signal is true;
	signal I14002: std_logic; attribute dont_touch of I14002: signal is true;
	signal I14003: std_logic; attribute dont_touch of I14003: signal is true;
	signal I14004: std_logic; attribute dont_touch of I14004: signal is true;
	signal I14005: std_logic; attribute dont_touch of I14005: signal is true;
	signal I14010: std_logic; attribute dont_touch of I14010: signal is true;
	signal I14011: std_logic; attribute dont_touch of I14011: signal is true;
	signal I14012: std_logic; attribute dont_touch of I14012: signal is true;
	signal I14017: std_logic; attribute dont_touch of I14017: signal is true;
	signal I14018: std_logic; attribute dont_touch of I14018: signal is true;
	signal I14019: std_logic; attribute dont_touch of I14019: signal is true;
	signal I14020: std_logic; attribute dont_touch of I14020: signal is true;
	signal I14025: std_logic; attribute dont_touch of I14025: signal is true;
	signal I14026: std_logic; attribute dont_touch of I14026: signal is true;
	signal I14027: std_logic; attribute dont_touch of I14027: signal is true;
	signal I14032: std_logic; attribute dont_touch of I14032: signal is true;
	signal I14033: std_logic; attribute dont_touch of I14033: signal is true;
	signal I14034: std_logic; attribute dont_touch of I14034: signal is true;
	signal I14035: std_logic; attribute dont_touch of I14035: signal is true;
	signal I14036: std_logic; attribute dont_touch of I14036: signal is true;
	signal I14041: std_logic; attribute dont_touch of I14041: signal is true;
	signal I14042: std_logic; attribute dont_touch of I14042: signal is true;
	signal I14043: std_logic; attribute dont_touch of I14043: signal is true;
	signal I14048: std_logic; attribute dont_touch of I14048: signal is true;
	signal I14049: std_logic; attribute dont_touch of I14049: signal is true;
	signal I14050: std_logic; attribute dont_touch of I14050: signal is true;
	signal I14051: std_logic; attribute dont_touch of I14051: signal is true;
	signal I14056: std_logic; attribute dont_touch of I14056: signal is true;
	signal I14057: std_logic; attribute dont_touch of I14057: signal is true;
	signal I14058: std_logic; attribute dont_touch of I14058: signal is true;
	signal I14063: std_logic; attribute dont_touch of I14063: signal is true;
	signal I14064: std_logic; attribute dont_touch of I14064: signal is true;
	signal I14065: std_logic; attribute dont_touch of I14065: signal is true;
	signal I14066: std_logic; attribute dont_touch of I14066: signal is true;
	signal I14067: std_logic; attribute dont_touch of I14067: signal is true;
	signal I14072: std_logic; attribute dont_touch of I14072: signal is true;
	signal I14073: std_logic; attribute dont_touch of I14073: signal is true;
	signal I14074: std_logic; attribute dont_touch of I14074: signal is true;
	signal I14079: std_logic; attribute dont_touch of I14079: signal is true;
	signal I14080: std_logic; attribute dont_touch of I14080: signal is true;
	signal I14081: std_logic; attribute dont_touch of I14081: signal is true;
	signal I14082: std_logic; attribute dont_touch of I14082: signal is true;
	signal I14087: std_logic; attribute dont_touch of I14087: signal is true;
	signal I14088: std_logic; attribute dont_touch of I14088: signal is true;
	signal I14089: std_logic; attribute dont_touch of I14089: signal is true;
	signal I14094: std_logic; attribute dont_touch of I14094: signal is true;
	signal I14095: std_logic; attribute dont_touch of I14095: signal is true;
	signal I14096: std_logic; attribute dont_touch of I14096: signal is true;
	signal I14097: std_logic; attribute dont_touch of I14097: signal is true;
	signal I14098: std_logic; attribute dont_touch of I14098: signal is true;
	signal I14103: std_logic; attribute dont_touch of I14103: signal is true;
	signal I14104: std_logic; attribute dont_touch of I14104: signal is true;
	signal I14105: std_logic; attribute dont_touch of I14105: signal is true;
	signal I14110: std_logic; attribute dont_touch of I14110: signal is true;
	signal I14111: std_logic; attribute dont_touch of I14111: signal is true;
	signal I14112: std_logic; attribute dont_touch of I14112: signal is true;
	signal I14113: std_logic; attribute dont_touch of I14113: signal is true;
	signal I14118: std_logic; attribute dont_touch of I14118: signal is true;
	signal I14119: std_logic; attribute dont_touch of I14119: signal is true;
	signal I14120: std_logic; attribute dont_touch of I14120: signal is true;
	signal I14125: std_logic; attribute dont_touch of I14125: signal is true;
	signal I14126: std_logic; attribute dont_touch of I14126: signal is true;
	signal I14127: std_logic; attribute dont_touch of I14127: signal is true;
	signal I14128: std_logic; attribute dont_touch of I14128: signal is true;
	signal I14129: std_logic; attribute dont_touch of I14129: signal is true;
	signal I14134: std_logic; attribute dont_touch of I14134: signal is true;
	signal I14135: std_logic; attribute dont_touch of I14135: signal is true;
	signal I14136: std_logic; attribute dont_touch of I14136: signal is true;
	signal I14141: std_logic; attribute dont_touch of I14141: signal is true;
	signal I14142: std_logic; attribute dont_touch of I14142: signal is true;
	signal I14143: std_logic; attribute dont_touch of I14143: signal is true;
	signal I14144: std_logic; attribute dont_touch of I14144: signal is true;
	signal I14149: std_logic; attribute dont_touch of I14149: signal is true;
	signal I14150: std_logic; attribute dont_touch of I14150: signal is true;
	signal I14151: std_logic; attribute dont_touch of I14151: signal is true;
	signal I14156: std_logic; attribute dont_touch of I14156: signal is true;
	signal I14157: std_logic; attribute dont_touch of I14157: signal is true;
	signal I14158: std_logic; attribute dont_touch of I14158: signal is true;
	signal I14159: std_logic; attribute dont_touch of I14159: signal is true;
	signal I14160: std_logic; attribute dont_touch of I14160: signal is true;
	signal I14165: std_logic; attribute dont_touch of I14165: signal is true;
	signal I14166: std_logic; attribute dont_touch of I14166: signal is true;
	signal I14167: std_logic; attribute dont_touch of I14167: signal is true;
	signal I14172: std_logic; attribute dont_touch of I14172: signal is true;
	signal I14173: std_logic; attribute dont_touch of I14173: signal is true;
	signal I14174: std_logic; attribute dont_touch of I14174: signal is true;
	signal I14175: std_logic; attribute dont_touch of I14175: signal is true;
	signal I14180: std_logic; attribute dont_touch of I14180: signal is true;
	signal I14181: std_logic; attribute dont_touch of I14181: signal is true;
	signal I14182: std_logic; attribute dont_touch of I14182: signal is true;
	signal I14187: std_logic; attribute dont_touch of I14187: signal is true;
	signal I14188: std_logic; attribute dont_touch of I14188: signal is true;
	signal I14189: std_logic; attribute dont_touch of I14189: signal is true;
	signal I14190: std_logic; attribute dont_touch of I14190: signal is true;
	signal I14191: std_logic; attribute dont_touch of I14191: signal is true;
	signal I14196: std_logic; attribute dont_touch of I14196: signal is true;
	signal I14197: std_logic; attribute dont_touch of I14197: signal is true;
	signal I14198: std_logic; attribute dont_touch of I14198: signal is true;
	signal I14203: std_logic; attribute dont_touch of I14203: signal is true;
	signal I14204: std_logic; attribute dont_touch of I14204: signal is true;
	signal I14205: std_logic; attribute dont_touch of I14205: signal is true;
	signal I14206: std_logic; attribute dont_touch of I14206: signal is true;
	signal I14211: std_logic; attribute dont_touch of I14211: signal is true;
	signal I14212: std_logic; attribute dont_touch of I14212: signal is true;
	signal I14213: std_logic; attribute dont_touch of I14213: signal is true;
	signal I14218: std_logic; attribute dont_touch of I14218: signal is true;
	signal I14219: std_logic; attribute dont_touch of I14219: signal is true;
	signal I14220: std_logic; attribute dont_touch of I14220: signal is true;
	signal I14221: std_logic; attribute dont_touch of I14221: signal is true;
	signal I14222: std_logic; attribute dont_touch of I14222: signal is true;
	signal I14227: std_logic; attribute dont_touch of I14227: signal is true;
	signal I14228: std_logic; attribute dont_touch of I14228: signal is true;
	signal I14229: std_logic; attribute dont_touch of I14229: signal is true;
	signal I14234: std_logic; attribute dont_touch of I14234: signal is true;
	signal I14235: std_logic; attribute dont_touch of I14235: signal is true;
	signal I14236: std_logic; attribute dont_touch of I14236: signal is true;
	signal I14237: std_logic; attribute dont_touch of I14237: signal is true;
	signal I14242: std_logic; attribute dont_touch of I14242: signal is true;
	signal I14243: std_logic; attribute dont_touch of I14243: signal is true;
	signal I14244: std_logic; attribute dont_touch of I14244: signal is true;
	signal I14249: std_logic; attribute dont_touch of I14249: signal is true;
	signal I14250: std_logic; attribute dont_touch of I14250: signal is true;
	signal I14251: std_logic; attribute dont_touch of I14251: signal is true;
	signal I14252: std_logic; attribute dont_touch of I14252: signal is true;
	signal I14253: std_logic; attribute dont_touch of I14253: signal is true;
	signal I14258: std_logic; attribute dont_touch of I14258: signal is true;
	signal I14259: std_logic; attribute dont_touch of I14259: signal is true;
	signal I14260: std_logic; attribute dont_touch of I14260: signal is true;
	signal I14265: std_logic; attribute dont_touch of I14265: signal is true;
	signal I14266: std_logic; attribute dont_touch of I14266: signal is true;
	signal I14267: std_logic; attribute dont_touch of I14267: signal is true;
	signal I14268: std_logic; attribute dont_touch of I14268: signal is true;
	signal I14273: std_logic; attribute dont_touch of I14273: signal is true;
	signal I14274: std_logic; attribute dont_touch of I14274: signal is true;
	signal I14275: std_logic; attribute dont_touch of I14275: signal is true;
	signal I14280: std_logic; attribute dont_touch of I14280: signal is true;
	signal I14281: std_logic; attribute dont_touch of I14281: signal is true;
	signal I14282: std_logic; attribute dont_touch of I14282: signal is true;
	signal I14283: std_logic; attribute dont_touch of I14283: signal is true;
	signal I14284: std_logic; attribute dont_touch of I14284: signal is true;
	signal I14289: std_logic; attribute dont_touch of I14289: signal is true;
	signal I14290: std_logic; attribute dont_touch of I14290: signal is true;
	signal I14291: std_logic; attribute dont_touch of I14291: signal is true;
	signal I14296: std_logic; attribute dont_touch of I14296: signal is true;
	signal I14297: std_logic; attribute dont_touch of I14297: signal is true;
	signal I14298: std_logic; attribute dont_touch of I14298: signal is true;
	signal I14299: std_logic; attribute dont_touch of I14299: signal is true;
	signal I14304: std_logic; attribute dont_touch of I14304: signal is true;
	signal I14305: std_logic; attribute dont_touch of I14305: signal is true;
	signal I14306: std_logic; attribute dont_touch of I14306: signal is true;
	signal I14311: std_logic; attribute dont_touch of I14311: signal is true;
	signal I14312: std_logic; attribute dont_touch of I14312: signal is true;
	signal I14313: std_logic; attribute dont_touch of I14313: signal is true;
	signal I14314: std_logic; attribute dont_touch of I14314: signal is true;
	signal I14315: std_logic; attribute dont_touch of I14315: signal is true;
	signal I14320: std_logic; attribute dont_touch of I14320: signal is true;
	signal I14321: std_logic; attribute dont_touch of I14321: signal is true;
	signal I14322: std_logic; attribute dont_touch of I14322: signal is true;
	signal I14327: std_logic; attribute dont_touch of I14327: signal is true;
	signal I14328: std_logic; attribute dont_touch of I14328: signal is true;
	signal I14329: std_logic; attribute dont_touch of I14329: signal is true;
	signal I14330: std_logic; attribute dont_touch of I14330: signal is true;
	signal I14335: std_logic; attribute dont_touch of I14335: signal is true;
	signal I14336: std_logic; attribute dont_touch of I14336: signal is true;
	signal I14337: std_logic; attribute dont_touch of I14337: signal is true;
	signal I14342: std_logic; attribute dont_touch of I14342: signal is true;
	signal I14343: std_logic; attribute dont_touch of I14343: signal is true;
	signal I14344: std_logic; attribute dont_touch of I14344: signal is true;
	signal I14345: std_logic; attribute dont_touch of I14345: signal is true;
	signal I14346: std_logic; attribute dont_touch of I14346: signal is true;
	signal I14351: std_logic; attribute dont_touch of I14351: signal is true;
	signal I14352: std_logic; attribute dont_touch of I14352: signal is true;
	signal I14353: std_logic; attribute dont_touch of I14353: signal is true;
	signal I14358: std_logic; attribute dont_touch of I14358: signal is true;
	signal I14359: std_logic; attribute dont_touch of I14359: signal is true;
	signal I14360: std_logic; attribute dont_touch of I14360: signal is true;
	signal I14361: std_logic; attribute dont_touch of I14361: signal is true;
	signal I14366: std_logic; attribute dont_touch of I14366: signal is true;
	signal I14367: std_logic; attribute dont_touch of I14367: signal is true;
	signal I14368: std_logic; attribute dont_touch of I14368: signal is true;
	signal I14373: std_logic; attribute dont_touch of I14373: signal is true;
	signal I14374: std_logic; attribute dont_touch of I14374: signal is true;
	signal I14375: std_logic; attribute dont_touch of I14375: signal is true;
	signal I14376: std_logic; attribute dont_touch of I14376: signal is true;
	signal I14377: std_logic; attribute dont_touch of I14377: signal is true;
	signal I14382: std_logic; attribute dont_touch of I14382: signal is true;
	signal I14383: std_logic; attribute dont_touch of I14383: signal is true;
	signal I14384: std_logic; attribute dont_touch of I14384: signal is true;
	signal I14389: std_logic; attribute dont_touch of I14389: signal is true;
	signal I14390: std_logic; attribute dont_touch of I14390: signal is true;
	signal I14391: std_logic; attribute dont_touch of I14391: signal is true;
	signal I14392: std_logic; attribute dont_touch of I14392: signal is true;
	signal I14397: std_logic; attribute dont_touch of I14397: signal is true;
	signal I14398: std_logic; attribute dont_touch of I14398: signal is true;
	signal I14399: std_logic; attribute dont_touch of I14399: signal is true;
	signal I14404: std_logic; attribute dont_touch of I14404: signal is true;
	signal I14405: std_logic; attribute dont_touch of I14405: signal is true;
	signal I14406: std_logic; attribute dont_touch of I14406: signal is true;
	signal I14407: std_logic; attribute dont_touch of I14407: signal is true;
	signal I14408: std_logic; attribute dont_touch of I14408: signal is true;
	signal I14413: std_logic; attribute dont_touch of I14413: signal is true;
	signal I14414: std_logic; attribute dont_touch of I14414: signal is true;
	signal I14415: std_logic; attribute dont_touch of I14415: signal is true;
	signal I14420: std_logic; attribute dont_touch of I14420: signal is true;
	signal I14421: std_logic; attribute dont_touch of I14421: signal is true;
	signal I14422: std_logic; attribute dont_touch of I14422: signal is true;
	signal I14423: std_logic; attribute dont_touch of I14423: signal is true;
	signal I14428: std_logic; attribute dont_touch of I14428: signal is true;
	signal I14429: std_logic; attribute dont_touch of I14429: signal is true;
	signal I14430: std_logic; attribute dont_touch of I14430: signal is true;
	signal I14435: std_logic; attribute dont_touch of I14435: signal is true;
	signal I14436: std_logic; attribute dont_touch of I14436: signal is true;
	signal I14437: std_logic; attribute dont_touch of I14437: signal is true;
	signal I14438: std_logic; attribute dont_touch of I14438: signal is true;
	signal I14439: std_logic; attribute dont_touch of I14439: signal is true;
	signal I14444: std_logic; attribute dont_touch of I14444: signal is true;
	signal I14445: std_logic; attribute dont_touch of I14445: signal is true;
	signal I14446: std_logic; attribute dont_touch of I14446: signal is true;
	signal I14451: std_logic; attribute dont_touch of I14451: signal is true;
	signal I14452: std_logic; attribute dont_touch of I14452: signal is true;
	signal I14453: std_logic; attribute dont_touch of I14453: signal is true;
	signal I14454: std_logic; attribute dont_touch of I14454: signal is true;
	signal I14459: std_logic; attribute dont_touch of I14459: signal is true;
	signal I14460: std_logic; attribute dont_touch of I14460: signal is true;
	signal I14461: std_logic; attribute dont_touch of I14461: signal is true;
	signal I14466: std_logic; attribute dont_touch of I14466: signal is true;
	signal I14467: std_logic; attribute dont_touch of I14467: signal is true;
	signal I14468: std_logic; attribute dont_touch of I14468: signal is true;
	signal I14469: std_logic; attribute dont_touch of I14469: signal is true;
	signal I14470: std_logic; attribute dont_touch of I14470: signal is true;
	signal I14475: std_logic; attribute dont_touch of I14475: signal is true;
	signal I14476: std_logic; attribute dont_touch of I14476: signal is true;
	signal I14477: std_logic; attribute dont_touch of I14477: signal is true;
	signal I14482: std_logic; attribute dont_touch of I14482: signal is true;
	signal I14483: std_logic; attribute dont_touch of I14483: signal is true;
	signal I14484: std_logic; attribute dont_touch of I14484: signal is true;
	signal I14485: std_logic; attribute dont_touch of I14485: signal is true;
	signal I14490: std_logic; attribute dont_touch of I14490: signal is true;
	signal I14491: std_logic; attribute dont_touch of I14491: signal is true;
	signal I14492: std_logic; attribute dont_touch of I14492: signal is true;
	signal I14497: std_logic; attribute dont_touch of I14497: signal is true;
	signal I14498: std_logic; attribute dont_touch of I14498: signal is true;
	signal I14499: std_logic; attribute dont_touch of I14499: signal is true;
	signal I14500: std_logic; attribute dont_touch of I14500: signal is true;
	signal I14501: std_logic; attribute dont_touch of I14501: signal is true;
	signal I14506: std_logic; attribute dont_touch of I14506: signal is true;
	signal I14507: std_logic; attribute dont_touch of I14507: signal is true;
	signal I14508: std_logic; attribute dont_touch of I14508: signal is true;
	signal I14513: std_logic; attribute dont_touch of I14513: signal is true;
	signal I14514: std_logic; attribute dont_touch of I14514: signal is true;
	signal I14515: std_logic; attribute dont_touch of I14515: signal is true;
	signal I14516: std_logic; attribute dont_touch of I14516: signal is true;
	signal I14521: std_logic; attribute dont_touch of I14521: signal is true;
	signal I14522: std_logic; attribute dont_touch of I14522: signal is true;
	signal I14523: std_logic; attribute dont_touch of I14523: signal is true;
	signal I14528: std_logic; attribute dont_touch of I14528: signal is true;
	signal I14529: std_logic; attribute dont_touch of I14529: signal is true;
	signal I14530: std_logic; attribute dont_touch of I14530: signal is true;
	signal I14531: std_logic; attribute dont_touch of I14531: signal is true;
	signal I14532: std_logic; attribute dont_touch of I14532: signal is true;
	signal I14537: std_logic; attribute dont_touch of I14537: signal is true;
	signal I14538: std_logic; attribute dont_touch of I14538: signal is true;
	signal I14539: std_logic; attribute dont_touch of I14539: signal is true;
	signal I14544: std_logic; attribute dont_touch of I14544: signal is true;
	signal I14545: std_logic; attribute dont_touch of I14545: signal is true;
	signal I14546: std_logic; attribute dont_touch of I14546: signal is true;
	signal I14547: std_logic; attribute dont_touch of I14547: signal is true;
	signal I14552: std_logic; attribute dont_touch of I14552: signal is true;
	signal I14553: std_logic; attribute dont_touch of I14553: signal is true;
	signal I14554: std_logic; attribute dont_touch of I14554: signal is true;
	signal I14559: std_logic; attribute dont_touch of I14559: signal is true;
	signal I14560: std_logic; attribute dont_touch of I14560: signal is true;
	signal I14561: std_logic; attribute dont_touch of I14561: signal is true;
	signal I14562: std_logic; attribute dont_touch of I14562: signal is true;
	signal I14563: std_logic; attribute dont_touch of I14563: signal is true;
	signal I14568: std_logic; attribute dont_touch of I14568: signal is true;
	signal I14569: std_logic; attribute dont_touch of I14569: signal is true;
	signal I14570: std_logic; attribute dont_touch of I14570: signal is true;
	signal I14575: std_logic; attribute dont_touch of I14575: signal is true;
	signal I14576: std_logic; attribute dont_touch of I14576: signal is true;
	signal I14577: std_logic; attribute dont_touch of I14577: signal is true;
	signal I14578: std_logic; attribute dont_touch of I14578: signal is true;
	signal I14583: std_logic; attribute dont_touch of I14583: signal is true;
	signal I14584: std_logic; attribute dont_touch of I14584: signal is true;
	signal I14585: std_logic; attribute dont_touch of I14585: signal is true;
	signal I14590: std_logic; attribute dont_touch of I14590: signal is true;
	signal I14591: std_logic; attribute dont_touch of I14591: signal is true;
	signal I14592: std_logic; attribute dont_touch of I14592: signal is true;
	signal I14593: std_logic; attribute dont_touch of I14593: signal is true;
	signal I14594: std_logic; attribute dont_touch of I14594: signal is true;
	signal I14599: std_logic; attribute dont_touch of I14599: signal is true;
	signal I14600: std_logic; attribute dont_touch of I14600: signal is true;
	signal I14601: std_logic; attribute dont_touch of I14601: signal is true;
	signal I14606: std_logic; attribute dont_touch of I14606: signal is true;
	signal I14607: std_logic; attribute dont_touch of I14607: signal is true;
	signal I14608: std_logic; attribute dont_touch of I14608: signal is true;
	signal I14609: std_logic; attribute dont_touch of I14609: signal is true;
	signal I14614: std_logic; attribute dont_touch of I14614: signal is true;
	signal I14615: std_logic; attribute dont_touch of I14615: signal is true;
	signal I14616: std_logic; attribute dont_touch of I14616: signal is true;
	signal I14621: std_logic; attribute dont_touch of I14621: signal is true;
	signal I14622: std_logic; attribute dont_touch of I14622: signal is true;
	signal I14623: std_logic; attribute dont_touch of I14623: signal is true;
	signal I14624: std_logic; attribute dont_touch of I14624: signal is true;
	signal I14625: std_logic; attribute dont_touch of I14625: signal is true;
	signal I14630: std_logic; attribute dont_touch of I14630: signal is true;
	signal I14631: std_logic; attribute dont_touch of I14631: signal is true;
	signal I14632: std_logic; attribute dont_touch of I14632: signal is true;
	signal I14637: std_logic; attribute dont_touch of I14637: signal is true;
	signal I14638: std_logic; attribute dont_touch of I14638: signal is true;
	signal I14639: std_logic; attribute dont_touch of I14639: signal is true;
	signal I14640: std_logic; attribute dont_touch of I14640: signal is true;
	signal I14645: std_logic; attribute dont_touch of I14645: signal is true;
	signal I14646: std_logic; attribute dont_touch of I14646: signal is true;
	signal I14647: std_logic; attribute dont_touch of I14647: signal is true;
	signal I14652: std_logic; attribute dont_touch of I14652: signal is true;
	signal I14653: std_logic; attribute dont_touch of I14653: signal is true;
	signal I14654: std_logic; attribute dont_touch of I14654: signal is true;
	signal I14655: std_logic; attribute dont_touch of I14655: signal is true;
	signal I14656: std_logic; attribute dont_touch of I14656: signal is true;
	signal I14661: std_logic; attribute dont_touch of I14661: signal is true;
	signal I14662: std_logic; attribute dont_touch of I14662: signal is true;
	signal I14663: std_logic; attribute dont_touch of I14663: signal is true;
	signal I14668: std_logic; attribute dont_touch of I14668: signal is true;
	signal I14669: std_logic; attribute dont_touch of I14669: signal is true;
	signal I14670: std_logic; attribute dont_touch of I14670: signal is true;
	signal I14671: std_logic; attribute dont_touch of I14671: signal is true;
	signal I14676: std_logic; attribute dont_touch of I14676: signal is true;
	signal I14677: std_logic; attribute dont_touch of I14677: signal is true;
	signal I14678: std_logic; attribute dont_touch of I14678: signal is true;
	signal I14683: std_logic; attribute dont_touch of I14683: signal is true;
	signal I14684: std_logic; attribute dont_touch of I14684: signal is true;
	signal I14685: std_logic; attribute dont_touch of I14685: signal is true;
	signal I14686: std_logic; attribute dont_touch of I14686: signal is true;
	signal I14687: std_logic; attribute dont_touch of I14687: signal is true;
	signal I14692: std_logic; attribute dont_touch of I14692: signal is true;
	signal I14693: std_logic; attribute dont_touch of I14693: signal is true;
	signal I14694: std_logic; attribute dont_touch of I14694: signal is true;
	signal I14699: std_logic; attribute dont_touch of I14699: signal is true;
	signal I14700: std_logic; attribute dont_touch of I14700: signal is true;
	signal I14701: std_logic; attribute dont_touch of I14701: signal is true;
	signal I14702: std_logic; attribute dont_touch of I14702: signal is true;
	signal I14707: std_logic; attribute dont_touch of I14707: signal is true;
	signal I14708: std_logic; attribute dont_touch of I14708: signal is true;
	signal I14709: std_logic; attribute dont_touch of I14709: signal is true;
	signal I14714: std_logic; attribute dont_touch of I14714: signal is true;
	signal I14715: std_logic; attribute dont_touch of I14715: signal is true;
	signal I14716: std_logic; attribute dont_touch of I14716: signal is true;
	signal I14717: std_logic; attribute dont_touch of I14717: signal is true;
	signal I14718: std_logic; attribute dont_touch of I14718: signal is true;
	signal I14723: std_logic; attribute dont_touch of I14723: signal is true;
	signal I14724: std_logic; attribute dont_touch of I14724: signal is true;
	signal I14725: std_logic; attribute dont_touch of I14725: signal is true;
	signal I14730: std_logic; attribute dont_touch of I14730: signal is true;
	signal I14731: std_logic; attribute dont_touch of I14731: signal is true;
	signal I14732: std_logic; attribute dont_touch of I14732: signal is true;
	signal I14733: std_logic; attribute dont_touch of I14733: signal is true;
	signal I14738: std_logic; attribute dont_touch of I14738: signal is true;
	signal I14739: std_logic; attribute dont_touch of I14739: signal is true;
	signal I14740: std_logic; attribute dont_touch of I14740: signal is true;
	signal I14745: std_logic; attribute dont_touch of I14745: signal is true;
	signal I14746: std_logic; attribute dont_touch of I14746: signal is true;
	signal I14747: std_logic; attribute dont_touch of I14747: signal is true;
	signal I14748: std_logic; attribute dont_touch of I14748: signal is true;
	signal I14749: std_logic; attribute dont_touch of I14749: signal is true;
	signal I14754: std_logic; attribute dont_touch of I14754: signal is true;
	signal I14755: std_logic; attribute dont_touch of I14755: signal is true;
	signal I14756: std_logic; attribute dont_touch of I14756: signal is true;
	signal I14761: std_logic; attribute dont_touch of I14761: signal is true;
	signal I14762: std_logic; attribute dont_touch of I14762: signal is true;
	signal I14763: std_logic; attribute dont_touch of I14763: signal is true;
	signal I14764: std_logic; attribute dont_touch of I14764: signal is true;
	signal I14769: std_logic; attribute dont_touch of I14769: signal is true;
	signal I14770: std_logic; attribute dont_touch of I14770: signal is true;
	signal I14771: std_logic; attribute dont_touch of I14771: signal is true;
	signal I14776: std_logic; attribute dont_touch of I14776: signal is true;
	signal I14777: std_logic; attribute dont_touch of I14777: signal is true;
	signal I14778: std_logic; attribute dont_touch of I14778: signal is true;
	signal I14779: std_logic; attribute dont_touch of I14779: signal is true;
	signal I14780: std_logic; attribute dont_touch of I14780: signal is true;
	signal I14785: std_logic; attribute dont_touch of I14785: signal is true;
	signal I14786: std_logic; attribute dont_touch of I14786: signal is true;
	signal I14787: std_logic; attribute dont_touch of I14787: signal is true;
	signal I14792: std_logic; attribute dont_touch of I14792: signal is true;
	signal I14793: std_logic; attribute dont_touch of I14793: signal is true;
	signal I14794: std_logic; attribute dont_touch of I14794: signal is true;
	signal I14795: std_logic; attribute dont_touch of I14795: signal is true;
	signal I14800: std_logic; attribute dont_touch of I14800: signal is true;
	signal I14801: std_logic; attribute dont_touch of I14801: signal is true;
	signal I14802: std_logic; attribute dont_touch of I14802: signal is true;
	signal I14807: std_logic; attribute dont_touch of I14807: signal is true;
	signal I14808: std_logic; attribute dont_touch of I14808: signal is true;
	signal I14809: std_logic; attribute dont_touch of I14809: signal is true;
	signal I14810: std_logic; attribute dont_touch of I14810: signal is true;
	signal I14811: std_logic; attribute dont_touch of I14811: signal is true;
	signal I14816: std_logic; attribute dont_touch of I14816: signal is true;
	signal I14817: std_logic; attribute dont_touch of I14817: signal is true;
	signal I14818: std_logic; attribute dont_touch of I14818: signal is true;
	signal I14823: std_logic; attribute dont_touch of I14823: signal is true;
	signal I14824: std_logic; attribute dont_touch of I14824: signal is true;
	signal I14825: std_logic; attribute dont_touch of I14825: signal is true;
	signal I14826: std_logic; attribute dont_touch of I14826: signal is true;
	signal I14831: std_logic; attribute dont_touch of I14831: signal is true;
	signal I14832: std_logic; attribute dont_touch of I14832: signal is true;
	signal I14833: std_logic; attribute dont_touch of I14833: signal is true;
	signal I14838: std_logic; attribute dont_touch of I14838: signal is true;
	signal I14839: std_logic; attribute dont_touch of I14839: signal is true;
	signal I14840: std_logic; attribute dont_touch of I14840: signal is true;
	signal I14841: std_logic; attribute dont_touch of I14841: signal is true;
	signal I14842: std_logic; attribute dont_touch of I14842: signal is true;
	signal I14847: std_logic; attribute dont_touch of I14847: signal is true;
	signal I14848: std_logic; attribute dont_touch of I14848: signal is true;
	signal I14849: std_logic; attribute dont_touch of I14849: signal is true;
	signal I14854: std_logic; attribute dont_touch of I14854: signal is true;
	signal I14855: std_logic; attribute dont_touch of I14855: signal is true;
	signal I14856: std_logic; attribute dont_touch of I14856: signal is true;
	signal I14857: std_logic; attribute dont_touch of I14857: signal is true;
	signal I14862: std_logic; attribute dont_touch of I14862: signal is true;
	signal I14863: std_logic; attribute dont_touch of I14863: signal is true;
	signal I14864: std_logic; attribute dont_touch of I14864: signal is true;
	signal I14869: std_logic; attribute dont_touch of I14869: signal is true;
	signal I14870: std_logic; attribute dont_touch of I14870: signal is true;
	signal I14871: std_logic; attribute dont_touch of I14871: signal is true;
	signal I14872: std_logic; attribute dont_touch of I14872: signal is true;
	signal I14873: std_logic; attribute dont_touch of I14873: signal is true;
	signal I14878: std_logic; attribute dont_touch of I14878: signal is true;
	signal I14879: std_logic; attribute dont_touch of I14879: signal is true;
	signal I14880: std_logic; attribute dont_touch of I14880: signal is true;
	signal I14885: std_logic; attribute dont_touch of I14885: signal is true;
	signal I14886: std_logic; attribute dont_touch of I14886: signal is true;
	signal I14887: std_logic; attribute dont_touch of I14887: signal is true;
	signal I14888: std_logic; attribute dont_touch of I14888: signal is true;
	signal I14893: std_logic; attribute dont_touch of I14893: signal is true;
	signal I14894: std_logic; attribute dont_touch of I14894: signal is true;
	signal I14895: std_logic; attribute dont_touch of I14895: signal is true;
	signal I14900: std_logic; attribute dont_touch of I14900: signal is true;
	signal I14901: std_logic; attribute dont_touch of I14901: signal is true;
	signal I14902: std_logic; attribute dont_touch of I14902: signal is true;
	signal I14903: std_logic; attribute dont_touch of I14903: signal is true;
	signal I14904: std_logic; attribute dont_touch of I14904: signal is true;
	signal I14909: std_logic; attribute dont_touch of I14909: signal is true;
	signal I14910: std_logic; attribute dont_touch of I14910: signal is true;
	signal I14911: std_logic; attribute dont_touch of I14911: signal is true;
	signal I14916: std_logic; attribute dont_touch of I14916: signal is true;
	signal I14917: std_logic; attribute dont_touch of I14917: signal is true;
	signal I14918: std_logic; attribute dont_touch of I14918: signal is true;
	signal I14919: std_logic; attribute dont_touch of I14919: signal is true;
	signal I14924: std_logic; attribute dont_touch of I14924: signal is true;
	signal I14925: std_logic; attribute dont_touch of I14925: signal is true;
	signal I14926: std_logic; attribute dont_touch of I14926: signal is true;
	signal I14931: std_logic; attribute dont_touch of I14931: signal is true;
	signal I14932: std_logic; attribute dont_touch of I14932: signal is true;
	signal I14933: std_logic; attribute dont_touch of I14933: signal is true;
	signal I14934: std_logic; attribute dont_touch of I14934: signal is true;
	signal I14935: std_logic; attribute dont_touch of I14935: signal is true;
	signal I14940: std_logic; attribute dont_touch of I14940: signal is true;
	signal I14941: std_logic; attribute dont_touch of I14941: signal is true;
	signal I14942: std_logic; attribute dont_touch of I14942: signal is true;
	signal I14947: std_logic; attribute dont_touch of I14947: signal is true;
	signal I14948: std_logic; attribute dont_touch of I14948: signal is true;
	signal I14949: std_logic; attribute dont_touch of I14949: signal is true;
	signal I14950: std_logic; attribute dont_touch of I14950: signal is true;
	signal I14955: std_logic; attribute dont_touch of I14955: signal is true;
	signal I14956: std_logic; attribute dont_touch of I14956: signal is true;
	signal I14957: std_logic; attribute dont_touch of I14957: signal is true;
	signal I14962: std_logic; attribute dont_touch of I14962: signal is true;
	signal I14963: std_logic; attribute dont_touch of I14963: signal is true;
	signal I14964: std_logic; attribute dont_touch of I14964: signal is true;
	signal I14965: std_logic; attribute dont_touch of I14965: signal is true;
	signal I14966: std_logic; attribute dont_touch of I14966: signal is true;
	signal I14971: std_logic; attribute dont_touch of I14971: signal is true;
	signal I14972: std_logic; attribute dont_touch of I14972: signal is true;
	signal I14973: std_logic; attribute dont_touch of I14973: signal is true;
	signal I14978: std_logic; attribute dont_touch of I14978: signal is true;
	signal I14979: std_logic; attribute dont_touch of I14979: signal is true;
	signal I14980: std_logic; attribute dont_touch of I14980: signal is true;
	signal I14981: std_logic; attribute dont_touch of I14981: signal is true;
	signal I14986: std_logic; attribute dont_touch of I14986: signal is true;
	signal I14987: std_logic; attribute dont_touch of I14987: signal is true;
	signal I14988: std_logic; attribute dont_touch of I14988: signal is true;
	signal I15067: std_logic; attribute dont_touch of I15067: signal is true;
	signal I15068: std_logic; attribute dont_touch of I15068: signal is true;
	signal I15069: std_logic; attribute dont_touch of I15069: signal is true;
	signal I15080: std_logic; attribute dont_touch of I15080: signal is true;
	signal I15081: std_logic; attribute dont_touch of I15081: signal is true;
	signal I15082: std_logic; attribute dont_touch of I15082: signal is true;
	signal I15093: std_logic; attribute dont_touch of I15093: signal is true;
	signal I15094: std_logic; attribute dont_touch of I15094: signal is true;
	signal I15095: std_logic; attribute dont_touch of I15095: signal is true;
	signal I15106: std_logic; attribute dont_touch of I15106: signal is true;
	signal I15107: std_logic; attribute dont_touch of I15107: signal is true;
	signal I15108: std_logic; attribute dont_touch of I15108: signal is true;
	signal I15119: std_logic; attribute dont_touch of I15119: signal is true;
	signal I15120: std_logic; attribute dont_touch of I15120: signal is true;
	signal I15121: std_logic; attribute dont_touch of I15121: signal is true;
	signal I15132: std_logic; attribute dont_touch of I15132: signal is true;
	signal I15133: std_logic; attribute dont_touch of I15133: signal is true;
	signal I15134: std_logic; attribute dont_touch of I15134: signal is true;
	signal I15145: std_logic; attribute dont_touch of I15145: signal is true;
	signal I15146: std_logic; attribute dont_touch of I15146: signal is true;
	signal I15147: std_logic; attribute dont_touch of I15147: signal is true;
	signal I15158: std_logic; attribute dont_touch of I15158: signal is true;
	signal I15159: std_logic; attribute dont_touch of I15159: signal is true;
	signal I15160: std_logic; attribute dont_touch of I15160: signal is true;
	signal I15171: std_logic; attribute dont_touch of I15171: signal is true;
	signal I15172: std_logic; attribute dont_touch of I15172: signal is true;
	signal I15173: std_logic; attribute dont_touch of I15173: signal is true;
	signal I15184: std_logic; attribute dont_touch of I15184: signal is true;
	signal I15185: std_logic; attribute dont_touch of I15185: signal is true;
	signal I15186: std_logic; attribute dont_touch of I15186: signal is true;
	signal I15197: std_logic; attribute dont_touch of I15197: signal is true;
	signal I15198: std_logic; attribute dont_touch of I15198: signal is true;
	signal I15199: std_logic; attribute dont_touch of I15199: signal is true;
	signal I15210: std_logic; attribute dont_touch of I15210: signal is true;
	signal I15211: std_logic; attribute dont_touch of I15211: signal is true;
	signal I15212: std_logic; attribute dont_touch of I15212: signal is true;
	signal I15223: std_logic; attribute dont_touch of I15223: signal is true;
	signal I15224: std_logic; attribute dont_touch of I15224: signal is true;
	signal I15225: std_logic; attribute dont_touch of I15225: signal is true;
	signal I15236: std_logic; attribute dont_touch of I15236: signal is true;
	signal I15237: std_logic; attribute dont_touch of I15237: signal is true;
	signal I15238: std_logic; attribute dont_touch of I15238: signal is true;
	signal I15249: std_logic; attribute dont_touch of I15249: signal is true;
	signal I15250: std_logic; attribute dont_touch of I15250: signal is true;
	signal I15251: std_logic; attribute dont_touch of I15251: signal is true;
	signal I15262: std_logic; attribute dont_touch of I15262: signal is true;
	signal I15263: std_logic; attribute dont_touch of I15263: signal is true;
	signal I15264: std_logic; attribute dont_touch of I15264: signal is true;
	signal I15275: std_logic; attribute dont_touch of I15275: signal is true;
	signal I15276: std_logic; attribute dont_touch of I15276: signal is true;
	signal I15277: std_logic; attribute dont_touch of I15277: signal is true;
	signal I15288: std_logic; attribute dont_touch of I15288: signal is true;
	signal I15289: std_logic; attribute dont_touch of I15289: signal is true;
	signal I15290: std_logic; attribute dont_touch of I15290: signal is true;
	signal I15301: std_logic; attribute dont_touch of I15301: signal is true;
	signal I15302: std_logic; attribute dont_touch of I15302: signal is true;
	signal I15303: std_logic; attribute dont_touch of I15303: signal is true;
	signal I15314: std_logic; attribute dont_touch of I15314: signal is true;
	signal I15315: std_logic; attribute dont_touch of I15315: signal is true;
	signal I15316: std_logic; attribute dont_touch of I15316: signal is true;
	signal I15327: std_logic; attribute dont_touch of I15327: signal is true;
	signal I15328: std_logic; attribute dont_touch of I15328: signal is true;
	signal I15329: std_logic; attribute dont_touch of I15329: signal is true;
	signal I15340: std_logic; attribute dont_touch of I15340: signal is true;
	signal I15341: std_logic; attribute dont_touch of I15341: signal is true;
	signal I15342: std_logic; attribute dont_touch of I15342: signal is true;
	signal I15353: std_logic; attribute dont_touch of I15353: signal is true;
	signal I15354: std_logic; attribute dont_touch of I15354: signal is true;
	signal I15355: std_logic; attribute dont_touch of I15355: signal is true;
	signal I15366: std_logic; attribute dont_touch of I15366: signal is true;
	signal I15367: std_logic; attribute dont_touch of I15367: signal is true;
	signal I15368: std_logic; attribute dont_touch of I15368: signal is true;
	signal I15379: std_logic; attribute dont_touch of I15379: signal is true;
	signal I15380: std_logic; attribute dont_touch of I15380: signal is true;
	signal I15381: std_logic; attribute dont_touch of I15381: signal is true;
	signal I15392: std_logic; attribute dont_touch of I15392: signal is true;
	signal I15393: std_logic; attribute dont_touch of I15393: signal is true;
	signal I15394: std_logic; attribute dont_touch of I15394: signal is true;
	signal I15405: std_logic; attribute dont_touch of I15405: signal is true;
	signal I15406: std_logic; attribute dont_touch of I15406: signal is true;
	signal I15407: std_logic; attribute dont_touch of I15407: signal is true;
	signal I15418: std_logic; attribute dont_touch of I15418: signal is true;
	signal I15419: std_logic; attribute dont_touch of I15419: signal is true;
	signal I15420: std_logic; attribute dont_touch of I15420: signal is true;
	signal I15431: std_logic; attribute dont_touch of I15431: signal is true;
	signal I15432: std_logic; attribute dont_touch of I15432: signal is true;
	signal I15433: std_logic; attribute dont_touch of I15433: signal is true;
	signal I15444: std_logic; attribute dont_touch of I15444: signal is true;
	signal I15445: std_logic; attribute dont_touch of I15445: signal is true;
	signal I15446: std_logic; attribute dont_touch of I15446: signal is true;
	signal I15457: std_logic; attribute dont_touch of I15457: signal is true;
	signal I15458: std_logic; attribute dont_touch of I15458: signal is true;
	signal I15459: std_logic; attribute dont_touch of I15459: signal is true;
	signal I15470: std_logic; attribute dont_touch of I15470: signal is true;
	signal I15471: std_logic; attribute dont_touch of I15471: signal is true;
	signal I15472: std_logic; attribute dont_touch of I15472: signal is true;
	signal I15484: std_logic; attribute dont_touch of I15484: signal is true;
	signal I15485: std_logic; attribute dont_touch of I15485: signal is true;
	signal I15486: std_logic; attribute dont_touch of I15486: signal is true;
	signal I15487: std_logic; attribute dont_touch of I15487: signal is true;
	signal I15492: std_logic; attribute dont_touch of I15492: signal is true;
	signal I15493: std_logic; attribute dont_touch of I15493: signal is true;
	signal I15494: std_logic; attribute dont_touch of I15494: signal is true;
	signal I15499: std_logic; attribute dont_touch of I15499: signal is true;
	signal I15500: std_logic; attribute dont_touch of I15500: signal is true;
	signal I15501: std_logic; attribute dont_touch of I15501: signal is true;
	signal I15502: std_logic; attribute dont_touch of I15502: signal is true;
	signal I15507: std_logic; attribute dont_touch of I15507: signal is true;
	signal I15508: std_logic; attribute dont_touch of I15508: signal is true;
	signal I15509: std_logic; attribute dont_touch of I15509: signal is true;
	signal I15514: std_logic; attribute dont_touch of I15514: signal is true;
	signal I15515: std_logic; attribute dont_touch of I15515: signal is true;
	signal I15516: std_logic; attribute dont_touch of I15516: signal is true;
	signal I15517: std_logic; attribute dont_touch of I15517: signal is true;
	signal I15522: std_logic; attribute dont_touch of I15522: signal is true;
	signal I15523: std_logic; attribute dont_touch of I15523: signal is true;
	signal I15524: std_logic; attribute dont_touch of I15524: signal is true;
	signal I15529: std_logic; attribute dont_touch of I15529: signal is true;
	signal I15530: std_logic; attribute dont_touch of I15530: signal is true;
	signal I15531: std_logic; attribute dont_touch of I15531: signal is true;
	signal I15536: std_logic; attribute dont_touch of I15536: signal is true;
	signal I15537: std_logic; attribute dont_touch of I15537: signal is true;
	signal I15538: std_logic; attribute dont_touch of I15538: signal is true;
	signal I15543: std_logic; attribute dont_touch of I15543: signal is true;
	signal I15544: std_logic; attribute dont_touch of I15544: signal is true;
	signal I15545: std_logic; attribute dont_touch of I15545: signal is true;
	signal I15550: std_logic; attribute dont_touch of I15550: signal is true;
	signal I15551: std_logic; attribute dont_touch of I15551: signal is true;
	signal I15552: std_logic; attribute dont_touch of I15552: signal is true;
	signal I15557: std_logic; attribute dont_touch of I15557: signal is true;
	signal I15558: std_logic; attribute dont_touch of I15558: signal is true;
	signal I15559: std_logic; attribute dont_touch of I15559: signal is true;
	signal I15564: std_logic; attribute dont_touch of I15564: signal is true;
	signal I15565: std_logic; attribute dont_touch of I15565: signal is true;
	signal I15566: std_logic; attribute dont_touch of I15566: signal is true;
	signal I15571: std_logic; attribute dont_touch of I15571: signal is true;
	signal I15572: std_logic; attribute dont_touch of I15572: signal is true;
	signal I15573: std_logic; attribute dont_touch of I15573: signal is true;
	signal I15578: std_logic; attribute dont_touch of I15578: signal is true;
	signal I15579: std_logic; attribute dont_touch of I15579: signal is true;
	signal I15580: std_logic; attribute dont_touch of I15580: signal is true;
	signal I15585: std_logic; attribute dont_touch of I15585: signal is true;
	signal I15586: std_logic; attribute dont_touch of I15586: signal is true;
	signal I15587: std_logic; attribute dont_touch of I15587: signal is true;
	signal I15592: std_logic; attribute dont_touch of I15592: signal is true;
	signal I15593: std_logic; attribute dont_touch of I15593: signal is true;
	signal I15594: std_logic; attribute dont_touch of I15594: signal is true;
	signal I15599: std_logic; attribute dont_touch of I15599: signal is true;
	signal I15600: std_logic; attribute dont_touch of I15600: signal is true;
	signal I15601: std_logic; attribute dont_touch of I15601: signal is true;
	signal I15606: std_logic; attribute dont_touch of I15606: signal is true;
	signal I15607: std_logic; attribute dont_touch of I15607: signal is true;
	signal I15608: std_logic; attribute dont_touch of I15608: signal is true;
	signal I15613: std_logic; attribute dont_touch of I15613: signal is true;
	signal I15614: std_logic; attribute dont_touch of I15614: signal is true;
	signal I15615: std_logic; attribute dont_touch of I15615: signal is true;
	signal I15620: std_logic; attribute dont_touch of I15620: signal is true;
	signal I15621: std_logic; attribute dont_touch of I15621: signal is true;
	signal I15622: std_logic; attribute dont_touch of I15622: signal is true;
	signal I15627: std_logic; attribute dont_touch of I15627: signal is true;
	signal I15628: std_logic; attribute dont_touch of I15628: signal is true;
	signal I15629: std_logic; attribute dont_touch of I15629: signal is true;
	signal I15634: std_logic; attribute dont_touch of I15634: signal is true;
	signal I15635: std_logic; attribute dont_touch of I15635: signal is true;
	signal I15636: std_logic; attribute dont_touch of I15636: signal is true;
	signal I15641: std_logic; attribute dont_touch of I15641: signal is true;
	signal I15642: std_logic; attribute dont_touch of I15642: signal is true;
	signal I15643: std_logic; attribute dont_touch of I15643: signal is true;
	signal I15648: std_logic; attribute dont_touch of I15648: signal is true;
	signal I15649: std_logic; attribute dont_touch of I15649: signal is true;
	signal I15650: std_logic; attribute dont_touch of I15650: signal is true;
	signal I15655: std_logic; attribute dont_touch of I15655: signal is true;
	signal I15656: std_logic; attribute dont_touch of I15656: signal is true;
	signal I15657: std_logic; attribute dont_touch of I15657: signal is true;
	signal I15662: std_logic; attribute dont_touch of I15662: signal is true;
	signal I15663: std_logic; attribute dont_touch of I15663: signal is true;
	signal I15664: std_logic; attribute dont_touch of I15664: signal is true;
	signal I15669: std_logic; attribute dont_touch of I15669: signal is true;
	signal I15670: std_logic; attribute dont_touch of I15670: signal is true;
	signal I15671: std_logic; attribute dont_touch of I15671: signal is true;
	signal I15676: std_logic; attribute dont_touch of I15676: signal is true;
	signal I15677: std_logic; attribute dont_touch of I15677: signal is true;
	signal I15678: std_logic; attribute dont_touch of I15678: signal is true;
	signal I15683: std_logic; attribute dont_touch of I15683: signal is true;
	signal I15684: std_logic; attribute dont_touch of I15684: signal is true;
	signal I15685: std_logic; attribute dont_touch of I15685: signal is true;
	signal I15690: std_logic; attribute dont_touch of I15690: signal is true;
	signal I15691: std_logic; attribute dont_touch of I15691: signal is true;
	signal I15692: std_logic; attribute dont_touch of I15692: signal is true;
	signal I15697: std_logic; attribute dont_touch of I15697: signal is true;
	signal I15698: std_logic; attribute dont_touch of I15698: signal is true;
	signal I15699: std_logic; attribute dont_touch of I15699: signal is true;
	signal I15704: std_logic; attribute dont_touch of I15704: signal is true;
	signal I15705: std_logic; attribute dont_touch of I15705: signal is true;
	signal I15706: std_logic; attribute dont_touch of I15706: signal is true;
	signal I15711: std_logic; attribute dont_touch of I15711: signal is true;
	signal I15712: std_logic; attribute dont_touch of I15712: signal is true;
	signal I15713: std_logic; attribute dont_touch of I15713: signal is true;
	signal I15718: std_logic; attribute dont_touch of I15718: signal is true;
	signal I15719: std_logic; attribute dont_touch of I15719: signal is true;
	signal I15720: std_logic; attribute dont_touch of I15720: signal is true;
	signal I15725: std_logic; attribute dont_touch of I15725: signal is true;
	signal I15726: std_logic; attribute dont_touch of I15726: signal is true;
	signal I15727: std_logic; attribute dont_touch of I15727: signal is true;
	signal I18006: std_logic; attribute dont_touch of I18006: signal is true;
	signal I18007: std_logic; attribute dont_touch of I18007: signal is true;
	signal I18008: std_logic; attribute dont_touch of I18008: signal is true;
	signal I18009: std_logic; attribute dont_touch of I18009: signal is true;
	signal I18010: std_logic; attribute dont_touch of I18010: signal is true;
	signal I18015: std_logic; attribute dont_touch of I18015: signal is true;
	signal I18016: std_logic; attribute dont_touch of I18016: signal is true;
	signal I18017: std_logic; attribute dont_touch of I18017: signal is true;
	signal I18022: std_logic; attribute dont_touch of I18022: signal is true;
	signal I18023: std_logic; attribute dont_touch of I18023: signal is true;
	signal I18024: std_logic; attribute dont_touch of I18024: signal is true;
	signal I18025: std_logic; attribute dont_touch of I18025: signal is true;
	signal I18030: std_logic; attribute dont_touch of I18030: signal is true;
	signal I18031: std_logic; attribute dont_touch of I18031: signal is true;
	signal I18032: std_logic; attribute dont_touch of I18032: signal is true;
	signal I18037: std_logic; attribute dont_touch of I18037: signal is true;
	signal I18038: std_logic; attribute dont_touch of I18038: signal is true;
	signal I18039: std_logic; attribute dont_touch of I18039: signal is true;
	signal I18040: std_logic; attribute dont_touch of I18040: signal is true;
	signal I18041: std_logic; attribute dont_touch of I18041: signal is true;
	signal I18046: std_logic; attribute dont_touch of I18046: signal is true;
	signal I18047: std_logic; attribute dont_touch of I18047: signal is true;
	signal I18048: std_logic; attribute dont_touch of I18048: signal is true;
	signal I18053: std_logic; attribute dont_touch of I18053: signal is true;
	signal I18054: std_logic; attribute dont_touch of I18054: signal is true;
	signal I18055: std_logic; attribute dont_touch of I18055: signal is true;
	signal I18056: std_logic; attribute dont_touch of I18056: signal is true;
	signal I18061: std_logic; attribute dont_touch of I18061: signal is true;
	signal I18062: std_logic; attribute dont_touch of I18062: signal is true;
	signal I18063: std_logic; attribute dont_touch of I18063: signal is true;
	signal I18068: std_logic; attribute dont_touch of I18068: signal is true;
	signal I18069: std_logic; attribute dont_touch of I18069: signal is true;
	signal I18070: std_logic; attribute dont_touch of I18070: signal is true;
	signal I18071: std_logic; attribute dont_touch of I18071: signal is true;
	signal I18072: std_logic; attribute dont_touch of I18072: signal is true;
	signal I18077: std_logic; attribute dont_touch of I18077: signal is true;
	signal I18078: std_logic; attribute dont_touch of I18078: signal is true;
	signal I18079: std_logic; attribute dont_touch of I18079: signal is true;
	signal I18084: std_logic; attribute dont_touch of I18084: signal is true;
	signal I18085: std_logic; attribute dont_touch of I18085: signal is true;
	signal I18086: std_logic; attribute dont_touch of I18086: signal is true;
	signal I18087: std_logic; attribute dont_touch of I18087: signal is true;
	signal I18092: std_logic; attribute dont_touch of I18092: signal is true;
	signal I18093: std_logic; attribute dont_touch of I18093: signal is true;
	signal I18094: std_logic; attribute dont_touch of I18094: signal is true;
	signal I18099: std_logic; attribute dont_touch of I18099: signal is true;
	signal I18100: std_logic; attribute dont_touch of I18100: signal is true;
	signal I18101: std_logic; attribute dont_touch of I18101: signal is true;
	signal I18102: std_logic; attribute dont_touch of I18102: signal is true;
	signal I18103: std_logic; attribute dont_touch of I18103: signal is true;
	signal I18108: std_logic; attribute dont_touch of I18108: signal is true;
	signal I18109: std_logic; attribute dont_touch of I18109: signal is true;
	signal I18110: std_logic; attribute dont_touch of I18110: signal is true;
	signal I18115: std_logic; attribute dont_touch of I18115: signal is true;
	signal I18116: std_logic; attribute dont_touch of I18116: signal is true;
	signal I18117: std_logic; attribute dont_touch of I18117: signal is true;
	signal I18118: std_logic; attribute dont_touch of I18118: signal is true;
	signal I18123: std_logic; attribute dont_touch of I18123: signal is true;
	signal I18124: std_logic; attribute dont_touch of I18124: signal is true;
	signal I18125: std_logic; attribute dont_touch of I18125: signal is true;
	signal I18130: std_logic; attribute dont_touch of I18130: signal is true;
	signal I18131: std_logic; attribute dont_touch of I18131: signal is true;
	signal I18132: std_logic; attribute dont_touch of I18132: signal is true;
	signal I18133: std_logic; attribute dont_touch of I18133: signal is true;
	signal I18134: std_logic; attribute dont_touch of I18134: signal is true;
	signal I18139: std_logic; attribute dont_touch of I18139: signal is true;
	signal I18140: std_logic; attribute dont_touch of I18140: signal is true;
	signal I18141: std_logic; attribute dont_touch of I18141: signal is true;
	signal I18146: std_logic; attribute dont_touch of I18146: signal is true;
	signal I18147: std_logic; attribute dont_touch of I18147: signal is true;
	signal I18148: std_logic; attribute dont_touch of I18148: signal is true;
	signal I18149: std_logic; attribute dont_touch of I18149: signal is true;
	signal I18154: std_logic; attribute dont_touch of I18154: signal is true;
	signal I18155: std_logic; attribute dont_touch of I18155: signal is true;
	signal I18156: std_logic; attribute dont_touch of I18156: signal is true;
	signal I18161: std_logic; attribute dont_touch of I18161: signal is true;
	signal I18162: std_logic; attribute dont_touch of I18162: signal is true;
	signal I18163: std_logic; attribute dont_touch of I18163: signal is true;
	signal I18164: std_logic; attribute dont_touch of I18164: signal is true;
	signal I18165: std_logic; attribute dont_touch of I18165: signal is true;
	signal I18170: std_logic; attribute dont_touch of I18170: signal is true;
	signal I18171: std_logic; attribute dont_touch of I18171: signal is true;
	signal I18172: std_logic; attribute dont_touch of I18172: signal is true;
	signal I18177: std_logic; attribute dont_touch of I18177: signal is true;
	signal I18178: std_logic; attribute dont_touch of I18178: signal is true;
	signal I18179: std_logic; attribute dont_touch of I18179: signal is true;
	signal I18180: std_logic; attribute dont_touch of I18180: signal is true;
	signal I18185: std_logic; attribute dont_touch of I18185: signal is true;
	signal I18186: std_logic; attribute dont_touch of I18186: signal is true;
	signal I18187: std_logic; attribute dont_touch of I18187: signal is true;
	signal I18192: std_logic; attribute dont_touch of I18192: signal is true;
	signal I18193: std_logic; attribute dont_touch of I18193: signal is true;
	signal I18194: std_logic; attribute dont_touch of I18194: signal is true;
	signal I18195: std_logic; attribute dont_touch of I18195: signal is true;
	signal I18196: std_logic; attribute dont_touch of I18196: signal is true;
	signal I18201: std_logic; attribute dont_touch of I18201: signal is true;
	signal I18202: std_logic; attribute dont_touch of I18202: signal is true;
	signal I18203: std_logic; attribute dont_touch of I18203: signal is true;
	signal I18208: std_logic; attribute dont_touch of I18208: signal is true;
	signal I18209: std_logic; attribute dont_touch of I18209: signal is true;
	signal I18210: std_logic; attribute dont_touch of I18210: signal is true;
	signal I18211: std_logic; attribute dont_touch of I18211: signal is true;
	signal I18216: std_logic; attribute dont_touch of I18216: signal is true;
	signal I18217: std_logic; attribute dont_touch of I18217: signal is true;
	signal I18218: std_logic; attribute dont_touch of I18218: signal is true;
	signal I18223: std_logic; attribute dont_touch of I18223: signal is true;
	signal I18224: std_logic; attribute dont_touch of I18224: signal is true;
	signal I18225: std_logic; attribute dont_touch of I18225: signal is true;
	signal I18226: std_logic; attribute dont_touch of I18226: signal is true;
	signal I18227: std_logic; attribute dont_touch of I18227: signal is true;
	signal I18232: std_logic; attribute dont_touch of I18232: signal is true;
	signal I18233: std_logic; attribute dont_touch of I18233: signal is true;
	signal I18234: std_logic; attribute dont_touch of I18234: signal is true;
	signal I18239: std_logic; attribute dont_touch of I18239: signal is true;
	signal I18240: std_logic; attribute dont_touch of I18240: signal is true;
	signal I18241: std_logic; attribute dont_touch of I18241: signal is true;
	signal I18242: std_logic; attribute dont_touch of I18242: signal is true;
	signal I18247: std_logic; attribute dont_touch of I18247: signal is true;
	signal I18248: std_logic; attribute dont_touch of I18248: signal is true;
	signal I18249: std_logic; attribute dont_touch of I18249: signal is true;
	signal I18254: std_logic; attribute dont_touch of I18254: signal is true;
	signal I18255: std_logic; attribute dont_touch of I18255: signal is true;
	signal I18256: std_logic; attribute dont_touch of I18256: signal is true;
	signal I18257: std_logic; attribute dont_touch of I18257: signal is true;
	signal I18258: std_logic; attribute dont_touch of I18258: signal is true;
	signal I18263: std_logic; attribute dont_touch of I18263: signal is true;
	signal I18264: std_logic; attribute dont_touch of I18264: signal is true;
	signal I18265: std_logic; attribute dont_touch of I18265: signal is true;
	signal I18270: std_logic; attribute dont_touch of I18270: signal is true;
	signal I18271: std_logic; attribute dont_touch of I18271: signal is true;
	signal I18272: std_logic; attribute dont_touch of I18272: signal is true;
	signal I18273: std_logic; attribute dont_touch of I18273: signal is true;
	signal I18278: std_logic; attribute dont_touch of I18278: signal is true;
	signal I18279: std_logic; attribute dont_touch of I18279: signal is true;
	signal I18280: std_logic; attribute dont_touch of I18280: signal is true;
	signal I18285: std_logic; attribute dont_touch of I18285: signal is true;
	signal I18286: std_logic; attribute dont_touch of I18286: signal is true;
	signal I18287: std_logic; attribute dont_touch of I18287: signal is true;
	signal I18288: std_logic; attribute dont_touch of I18288: signal is true;
	signal I18289: std_logic; attribute dont_touch of I18289: signal is true;
	signal I18294: std_logic; attribute dont_touch of I18294: signal is true;
	signal I18295: std_logic; attribute dont_touch of I18295: signal is true;
	signal I18296: std_logic; attribute dont_touch of I18296: signal is true;
	signal I18301: std_logic; attribute dont_touch of I18301: signal is true;
	signal I18302: std_logic; attribute dont_touch of I18302: signal is true;
	signal I18303: std_logic; attribute dont_touch of I18303: signal is true;
	signal I18304: std_logic; attribute dont_touch of I18304: signal is true;
	signal I18309: std_logic; attribute dont_touch of I18309: signal is true;
	signal I18310: std_logic; attribute dont_touch of I18310: signal is true;
	signal I18311: std_logic; attribute dont_touch of I18311: signal is true;
	signal I18316: std_logic; attribute dont_touch of I18316: signal is true;
	signal I18317: std_logic; attribute dont_touch of I18317: signal is true;
	signal I18318: std_logic; attribute dont_touch of I18318: signal is true;
	signal I18319: std_logic; attribute dont_touch of I18319: signal is true;
	signal I18320: std_logic; attribute dont_touch of I18320: signal is true;
	signal I18325: std_logic; attribute dont_touch of I18325: signal is true;
	signal I18326: std_logic; attribute dont_touch of I18326: signal is true;
	signal I18327: std_logic; attribute dont_touch of I18327: signal is true;
	signal I18332: std_logic; attribute dont_touch of I18332: signal is true;
	signal I18333: std_logic; attribute dont_touch of I18333: signal is true;
	signal I18334: std_logic; attribute dont_touch of I18334: signal is true;
	signal I18335: std_logic; attribute dont_touch of I18335: signal is true;
	signal I18340: std_logic; attribute dont_touch of I18340: signal is true;
	signal I18341: std_logic; attribute dont_touch of I18341: signal is true;
	signal I18342: std_logic; attribute dont_touch of I18342: signal is true;
	signal I18347: std_logic; attribute dont_touch of I18347: signal is true;
	signal I18348: std_logic; attribute dont_touch of I18348: signal is true;
	signal I18349: std_logic; attribute dont_touch of I18349: signal is true;
	signal I18350: std_logic; attribute dont_touch of I18350: signal is true;
	signal I18351: std_logic; attribute dont_touch of I18351: signal is true;
	signal I18356: std_logic; attribute dont_touch of I18356: signal is true;
	signal I18357: std_logic; attribute dont_touch of I18357: signal is true;
	signal I18358: std_logic; attribute dont_touch of I18358: signal is true;
	signal I18363: std_logic; attribute dont_touch of I18363: signal is true;
	signal I18364: std_logic; attribute dont_touch of I18364: signal is true;
	signal I18365: std_logic; attribute dont_touch of I18365: signal is true;
	signal I18366: std_logic; attribute dont_touch of I18366: signal is true;
	signal I18371: std_logic; attribute dont_touch of I18371: signal is true;
	signal I18372: std_logic; attribute dont_touch of I18372: signal is true;
	signal I18373: std_logic; attribute dont_touch of I18373: signal is true;
	signal I18378: std_logic; attribute dont_touch of I18378: signal is true;
	signal I18379: std_logic; attribute dont_touch of I18379: signal is true;
	signal I18380: std_logic; attribute dont_touch of I18380: signal is true;
	signal I18381: std_logic; attribute dont_touch of I18381: signal is true;
	signal I18382: std_logic; attribute dont_touch of I18382: signal is true;
	signal I18387: std_logic; attribute dont_touch of I18387: signal is true;
	signal I18388: std_logic; attribute dont_touch of I18388: signal is true;
	signal I18389: std_logic; attribute dont_touch of I18389: signal is true;
	signal I18394: std_logic; attribute dont_touch of I18394: signal is true;
	signal I18395: std_logic; attribute dont_touch of I18395: signal is true;
	signal I18396: std_logic; attribute dont_touch of I18396: signal is true;
	signal I18397: std_logic; attribute dont_touch of I18397: signal is true;
	signal I18402: std_logic; attribute dont_touch of I18402: signal is true;
	signal I18403: std_logic; attribute dont_touch of I18403: signal is true;
	signal I18404: std_logic; attribute dont_touch of I18404: signal is true;
	signal I18409: std_logic; attribute dont_touch of I18409: signal is true;
	signal I18410: std_logic; attribute dont_touch of I18410: signal is true;
	signal I18411: std_logic; attribute dont_touch of I18411: signal is true;
	signal I18412: std_logic; attribute dont_touch of I18412: signal is true;
	signal I18413: std_logic; attribute dont_touch of I18413: signal is true;
	signal I18418: std_logic; attribute dont_touch of I18418: signal is true;
	signal I18419: std_logic; attribute dont_touch of I18419: signal is true;
	signal I18420: std_logic; attribute dont_touch of I18420: signal is true;
	signal I18425: std_logic; attribute dont_touch of I18425: signal is true;
	signal I18426: std_logic; attribute dont_touch of I18426: signal is true;
	signal I18427: std_logic; attribute dont_touch of I18427: signal is true;
	signal I18428: std_logic; attribute dont_touch of I18428: signal is true;
	signal I18433: std_logic; attribute dont_touch of I18433: signal is true;
	signal I18434: std_logic; attribute dont_touch of I18434: signal is true;
	signal I18435: std_logic; attribute dont_touch of I18435: signal is true;
	signal I18440: std_logic; attribute dont_touch of I18440: signal is true;
	signal I18441: std_logic; attribute dont_touch of I18441: signal is true;
	signal I18442: std_logic; attribute dont_touch of I18442: signal is true;
	signal I18443: std_logic; attribute dont_touch of I18443: signal is true;
	signal I18444: std_logic; attribute dont_touch of I18444: signal is true;
	signal I18449: std_logic; attribute dont_touch of I18449: signal is true;
	signal I18450: std_logic; attribute dont_touch of I18450: signal is true;
	signal I18451: std_logic; attribute dont_touch of I18451: signal is true;
	signal I18456: std_logic; attribute dont_touch of I18456: signal is true;
	signal I18457: std_logic; attribute dont_touch of I18457: signal is true;
	signal I18458: std_logic; attribute dont_touch of I18458: signal is true;
	signal I18459: std_logic; attribute dont_touch of I18459: signal is true;
	signal I18464: std_logic; attribute dont_touch of I18464: signal is true;
	signal I18465: std_logic; attribute dont_touch of I18465: signal is true;
	signal I18466: std_logic; attribute dont_touch of I18466: signal is true;
	signal I18471: std_logic; attribute dont_touch of I18471: signal is true;
	signal I18472: std_logic; attribute dont_touch of I18472: signal is true;
	signal I18473: std_logic; attribute dont_touch of I18473: signal is true;
	signal I18474: std_logic; attribute dont_touch of I18474: signal is true;
	signal I18475: std_logic; attribute dont_touch of I18475: signal is true;
	signal I18480: std_logic; attribute dont_touch of I18480: signal is true;
	signal I18481: std_logic; attribute dont_touch of I18481: signal is true;
	signal I18482: std_logic; attribute dont_touch of I18482: signal is true;
	signal I18487: std_logic; attribute dont_touch of I18487: signal is true;
	signal I18488: std_logic; attribute dont_touch of I18488: signal is true;
	signal I18489: std_logic; attribute dont_touch of I18489: signal is true;
	signal I18490: std_logic; attribute dont_touch of I18490: signal is true;
	signal I18495: std_logic; attribute dont_touch of I18495: signal is true;
	signal I18496: std_logic; attribute dont_touch of I18496: signal is true;
	signal I18497: std_logic; attribute dont_touch of I18497: signal is true;
	signal I18502: std_logic; attribute dont_touch of I18502: signal is true;
	signal I18503: std_logic; attribute dont_touch of I18503: signal is true;
	signal I18504: std_logic; attribute dont_touch of I18504: signal is true;
	signal I18505: std_logic; attribute dont_touch of I18505: signal is true;
	signal I18506: std_logic; attribute dont_touch of I18506: signal is true;
	signal I18511: std_logic; attribute dont_touch of I18511: signal is true;
	signal I18512: std_logic; attribute dont_touch of I18512: signal is true;
	signal I18513: std_logic; attribute dont_touch of I18513: signal is true;
	signal I18518: std_logic; attribute dont_touch of I18518: signal is true;
	signal I18519: std_logic; attribute dont_touch of I18519: signal is true;
	signal I18520: std_logic; attribute dont_touch of I18520: signal is true;
	signal I18521: std_logic; attribute dont_touch of I18521: signal is true;
	signal I18526: std_logic; attribute dont_touch of I18526: signal is true;
	signal I18527: std_logic; attribute dont_touch of I18527: signal is true;
	signal I18528: std_logic; attribute dont_touch of I18528: signal is true;
	signal I18533: std_logic; attribute dont_touch of I18533: signal is true;
	signal I18534: std_logic; attribute dont_touch of I18534: signal is true;
	signal I18535: std_logic; attribute dont_touch of I18535: signal is true;
	signal I18536: std_logic; attribute dont_touch of I18536: signal is true;
	signal I18537: std_logic; attribute dont_touch of I18537: signal is true;
	signal I18542: std_logic; attribute dont_touch of I18542: signal is true;
	signal I18543: std_logic; attribute dont_touch of I18543: signal is true;
	signal I18544: std_logic; attribute dont_touch of I18544: signal is true;
	signal I18549: std_logic; attribute dont_touch of I18549: signal is true;
	signal I18550: std_logic; attribute dont_touch of I18550: signal is true;
	signal I18551: std_logic; attribute dont_touch of I18551: signal is true;
	signal I18552: std_logic; attribute dont_touch of I18552: signal is true;
	signal I18557: std_logic; attribute dont_touch of I18557: signal is true;
	signal I18558: std_logic; attribute dont_touch of I18558: signal is true;
	signal I18559: std_logic; attribute dont_touch of I18559: signal is true;
	signal I18564: std_logic; attribute dont_touch of I18564: signal is true;
	signal I18565: std_logic; attribute dont_touch of I18565: signal is true;
	signal I18566: std_logic; attribute dont_touch of I18566: signal is true;
	signal I18567: std_logic; attribute dont_touch of I18567: signal is true;
	signal I18568: std_logic; attribute dont_touch of I18568: signal is true;
	signal I18573: std_logic; attribute dont_touch of I18573: signal is true;
	signal I18574: std_logic; attribute dont_touch of I18574: signal is true;
	signal I18575: std_logic; attribute dont_touch of I18575: signal is true;
	signal I18580: std_logic; attribute dont_touch of I18580: signal is true;
	signal I18581: std_logic; attribute dont_touch of I18581: signal is true;
	signal I18582: std_logic; attribute dont_touch of I18582: signal is true;
	signal I18583: std_logic; attribute dont_touch of I18583: signal is true;
	signal I18588: std_logic; attribute dont_touch of I18588: signal is true;
	signal I18589: std_logic; attribute dont_touch of I18589: signal is true;
	signal I18590: std_logic; attribute dont_touch of I18590: signal is true;
	signal I18595: std_logic; attribute dont_touch of I18595: signal is true;
	signal I18596: std_logic; attribute dont_touch of I18596: signal is true;
	signal I18597: std_logic; attribute dont_touch of I18597: signal is true;
	signal I18598: std_logic; attribute dont_touch of I18598: signal is true;
	signal I18599: std_logic; attribute dont_touch of I18599: signal is true;
	signal I18604: std_logic; attribute dont_touch of I18604: signal is true;
	signal I18605: std_logic; attribute dont_touch of I18605: signal is true;
	signal I18606: std_logic; attribute dont_touch of I18606: signal is true;
	signal I18611: std_logic; attribute dont_touch of I18611: signal is true;
	signal I18612: std_logic; attribute dont_touch of I18612: signal is true;
	signal I18613: std_logic; attribute dont_touch of I18613: signal is true;
	signal I18614: std_logic; attribute dont_touch of I18614: signal is true;
	signal I18619: std_logic; attribute dont_touch of I18619: signal is true;
	signal I18620: std_logic; attribute dont_touch of I18620: signal is true;
	signal I18621: std_logic; attribute dont_touch of I18621: signal is true;
	signal I18626: std_logic; attribute dont_touch of I18626: signal is true;
	signal I18627: std_logic; attribute dont_touch of I18627: signal is true;
	signal I18628: std_logic; attribute dont_touch of I18628: signal is true;
	signal I18629: std_logic; attribute dont_touch of I18629: signal is true;
	signal I18630: std_logic; attribute dont_touch of I18630: signal is true;
	signal I18635: std_logic; attribute dont_touch of I18635: signal is true;
	signal I18636: std_logic; attribute dont_touch of I18636: signal is true;
	signal I18637: std_logic; attribute dont_touch of I18637: signal is true;
	signal I18642: std_logic; attribute dont_touch of I18642: signal is true;
	signal I18643: std_logic; attribute dont_touch of I18643: signal is true;
	signal I18644: std_logic; attribute dont_touch of I18644: signal is true;
	signal I18645: std_logic; attribute dont_touch of I18645: signal is true;
	signal I18650: std_logic; attribute dont_touch of I18650: signal is true;
	signal I18651: std_logic; attribute dont_touch of I18651: signal is true;
	signal I18652: std_logic; attribute dont_touch of I18652: signal is true;
	signal I18657: std_logic; attribute dont_touch of I18657: signal is true;
	signal I18658: std_logic; attribute dont_touch of I18658: signal is true;
	signal I18659: std_logic; attribute dont_touch of I18659: signal is true;
	signal I18660: std_logic; attribute dont_touch of I18660: signal is true;
	signal I18661: std_logic; attribute dont_touch of I18661: signal is true;
	signal I18666: std_logic; attribute dont_touch of I18666: signal is true;
	signal I18667: std_logic; attribute dont_touch of I18667: signal is true;
	signal I18668: std_logic; attribute dont_touch of I18668: signal is true;
	signal I18673: std_logic; attribute dont_touch of I18673: signal is true;
	signal I18674: std_logic; attribute dont_touch of I18674: signal is true;
	signal I18675: std_logic; attribute dont_touch of I18675: signal is true;
	signal I18676: std_logic; attribute dont_touch of I18676: signal is true;
	signal I18681: std_logic; attribute dont_touch of I18681: signal is true;
	signal I18682: std_logic; attribute dont_touch of I18682: signal is true;
	signal I18683: std_logic; attribute dont_touch of I18683: signal is true;
	signal I18688: std_logic; attribute dont_touch of I18688: signal is true;
	signal I18689: std_logic; attribute dont_touch of I18689: signal is true;
	signal I18690: std_logic; attribute dont_touch of I18690: signal is true;
	signal I18691: std_logic; attribute dont_touch of I18691: signal is true;
	signal I18692: std_logic; attribute dont_touch of I18692: signal is true;
	signal I18697: std_logic; attribute dont_touch of I18697: signal is true;
	signal I18698: std_logic; attribute dont_touch of I18698: signal is true;
	signal I18699: std_logic; attribute dont_touch of I18699: signal is true;
	signal I18704: std_logic; attribute dont_touch of I18704: signal is true;
	signal I18705: std_logic; attribute dont_touch of I18705: signal is true;
	signal I18706: std_logic; attribute dont_touch of I18706: signal is true;
	signal I18707: std_logic; attribute dont_touch of I18707: signal is true;
	signal I18712: std_logic; attribute dont_touch of I18712: signal is true;
	signal I18713: std_logic; attribute dont_touch of I18713: signal is true;
	signal I18714: std_logic; attribute dont_touch of I18714: signal is true;
	signal I18719: std_logic; attribute dont_touch of I18719: signal is true;
	signal I18720: std_logic; attribute dont_touch of I18720: signal is true;
	signal I18721: std_logic; attribute dont_touch of I18721: signal is true;
	signal I18722: std_logic; attribute dont_touch of I18722: signal is true;
	signal I18723: std_logic; attribute dont_touch of I18723: signal is true;
	signal I18728: std_logic; attribute dont_touch of I18728: signal is true;
	signal I18729: std_logic; attribute dont_touch of I18729: signal is true;
	signal I18730: std_logic; attribute dont_touch of I18730: signal is true;
	signal I18735: std_logic; attribute dont_touch of I18735: signal is true;
	signal I18736: std_logic; attribute dont_touch of I18736: signal is true;
	signal I18737: std_logic; attribute dont_touch of I18737: signal is true;
	signal I18738: std_logic; attribute dont_touch of I18738: signal is true;
	signal I18743: std_logic; attribute dont_touch of I18743: signal is true;
	signal I18744: std_logic; attribute dont_touch of I18744: signal is true;
	signal I18745: std_logic; attribute dont_touch of I18745: signal is true;
	signal I18750: std_logic; attribute dont_touch of I18750: signal is true;
	signal I18751: std_logic; attribute dont_touch of I18751: signal is true;
	signal I18752: std_logic; attribute dont_touch of I18752: signal is true;
	signal I18753: std_logic; attribute dont_touch of I18753: signal is true;
	signal I18754: std_logic; attribute dont_touch of I18754: signal is true;
	signal I18759: std_logic; attribute dont_touch of I18759: signal is true;
	signal I18760: std_logic; attribute dont_touch of I18760: signal is true;
	signal I18761: std_logic; attribute dont_touch of I18761: signal is true;
	signal I18766: std_logic; attribute dont_touch of I18766: signal is true;
	signal I18767: std_logic; attribute dont_touch of I18767: signal is true;
	signal I18768: std_logic; attribute dont_touch of I18768: signal is true;
	signal I18769: std_logic; attribute dont_touch of I18769: signal is true;
	signal I18774: std_logic; attribute dont_touch of I18774: signal is true;
	signal I18775: std_logic; attribute dont_touch of I18775: signal is true;
	signal I18776: std_logic; attribute dont_touch of I18776: signal is true;
	signal I18781: std_logic; attribute dont_touch of I18781: signal is true;
	signal I18782: std_logic; attribute dont_touch of I18782: signal is true;
	signal I18783: std_logic; attribute dont_touch of I18783: signal is true;
	signal I18784: std_logic; attribute dont_touch of I18784: signal is true;
	signal I18785: std_logic; attribute dont_touch of I18785: signal is true;
	signal I18790: std_logic; attribute dont_touch of I18790: signal is true;
	signal I18791: std_logic; attribute dont_touch of I18791: signal is true;
	signal I18792: std_logic; attribute dont_touch of I18792: signal is true;
	signal I18797: std_logic; attribute dont_touch of I18797: signal is true;
	signal I18798: std_logic; attribute dont_touch of I18798: signal is true;
	signal I18799: std_logic; attribute dont_touch of I18799: signal is true;
	signal I18800: std_logic; attribute dont_touch of I18800: signal is true;
	signal I18805: std_logic; attribute dont_touch of I18805: signal is true;
	signal I18806: std_logic; attribute dont_touch of I18806: signal is true;
	signal I18807: std_logic; attribute dont_touch of I18807: signal is true;
	signal I18812: std_logic; attribute dont_touch of I18812: signal is true;
	signal I18813: std_logic; attribute dont_touch of I18813: signal is true;
	signal I18814: std_logic; attribute dont_touch of I18814: signal is true;
	signal I18815: std_logic; attribute dont_touch of I18815: signal is true;
	signal I18816: std_logic; attribute dont_touch of I18816: signal is true;
	signal I18821: std_logic; attribute dont_touch of I18821: signal is true;
	signal I18822: std_logic; attribute dont_touch of I18822: signal is true;
	signal I18823: std_logic; attribute dont_touch of I18823: signal is true;
	signal I18828: std_logic; attribute dont_touch of I18828: signal is true;
	signal I18829: std_logic; attribute dont_touch of I18829: signal is true;
	signal I18830: std_logic; attribute dont_touch of I18830: signal is true;
	signal I18831: std_logic; attribute dont_touch of I18831: signal is true;
	signal I18836: std_logic; attribute dont_touch of I18836: signal is true;
	signal I18837: std_logic; attribute dont_touch of I18837: signal is true;
	signal I18838: std_logic; attribute dont_touch of I18838: signal is true;
	signal I18843: std_logic; attribute dont_touch of I18843: signal is true;
	signal I18844: std_logic; attribute dont_touch of I18844: signal is true;
	signal I18845: std_logic; attribute dont_touch of I18845: signal is true;
	signal I18846: std_logic; attribute dont_touch of I18846: signal is true;
	signal I18847: std_logic; attribute dont_touch of I18847: signal is true;
	signal I18852: std_logic; attribute dont_touch of I18852: signal is true;
	signal I18853: std_logic; attribute dont_touch of I18853: signal is true;
	signal I18854: std_logic; attribute dont_touch of I18854: signal is true;
	signal I18859: std_logic; attribute dont_touch of I18859: signal is true;
	signal I18860: std_logic; attribute dont_touch of I18860: signal is true;
	signal I18861: std_logic; attribute dont_touch of I18861: signal is true;
	signal I18862: std_logic; attribute dont_touch of I18862: signal is true;
	signal I18867: std_logic; attribute dont_touch of I18867: signal is true;
	signal I18868: std_logic; attribute dont_touch of I18868: signal is true;
	signal I18869: std_logic; attribute dont_touch of I18869: signal is true;
	signal I18874: std_logic; attribute dont_touch of I18874: signal is true;
	signal I18875: std_logic; attribute dont_touch of I18875: signal is true;
	signal I18876: std_logic; attribute dont_touch of I18876: signal is true;
	signal I18877: std_logic; attribute dont_touch of I18877: signal is true;
	signal I18878: std_logic; attribute dont_touch of I18878: signal is true;
	signal I18883: std_logic; attribute dont_touch of I18883: signal is true;
	signal I18884: std_logic; attribute dont_touch of I18884: signal is true;
	signal I18885: std_logic; attribute dont_touch of I18885: signal is true;
	signal I18890: std_logic; attribute dont_touch of I18890: signal is true;
	signal I18891: std_logic; attribute dont_touch of I18891: signal is true;
	signal I18892: std_logic; attribute dont_touch of I18892: signal is true;
	signal I18893: std_logic; attribute dont_touch of I18893: signal is true;
	signal I18898: std_logic; attribute dont_touch of I18898: signal is true;
	signal I18899: std_logic; attribute dont_touch of I18899: signal is true;
	signal I18900: std_logic; attribute dont_touch of I18900: signal is true;
	signal I18905: std_logic; attribute dont_touch of I18905: signal is true;
	signal I18906: std_logic; attribute dont_touch of I18906: signal is true;
	signal I18907: std_logic; attribute dont_touch of I18907: signal is true;
	signal I18908: std_logic; attribute dont_touch of I18908: signal is true;
	signal I18909: std_logic; attribute dont_touch of I18909: signal is true;
	signal I18914: std_logic; attribute dont_touch of I18914: signal is true;
	signal I18915: std_logic; attribute dont_touch of I18915: signal is true;
	signal I18916: std_logic; attribute dont_touch of I18916: signal is true;
	signal I18921: std_logic; attribute dont_touch of I18921: signal is true;
	signal I18922: std_logic; attribute dont_touch of I18922: signal is true;
	signal I18923: std_logic; attribute dont_touch of I18923: signal is true;
	signal I18924: std_logic; attribute dont_touch of I18924: signal is true;
	signal I18929: std_logic; attribute dont_touch of I18929: signal is true;
	signal I18930: std_logic; attribute dont_touch of I18930: signal is true;
	signal I18931: std_logic; attribute dont_touch of I18931: signal is true;
	signal I18936: std_logic; attribute dont_touch of I18936: signal is true;
	signal I18937: std_logic; attribute dont_touch of I18937: signal is true;
	signal I18938: std_logic; attribute dont_touch of I18938: signal is true;
	signal I18939: std_logic; attribute dont_touch of I18939: signal is true;
	signal I18940: std_logic; attribute dont_touch of I18940: signal is true;
	signal I18945: std_logic; attribute dont_touch of I18945: signal is true;
	signal I18946: std_logic; attribute dont_touch of I18946: signal is true;
	signal I18947: std_logic; attribute dont_touch of I18947: signal is true;
	signal I18952: std_logic; attribute dont_touch of I18952: signal is true;
	signal I18953: std_logic; attribute dont_touch of I18953: signal is true;
	signal I18954: std_logic; attribute dont_touch of I18954: signal is true;
	signal I18955: std_logic; attribute dont_touch of I18955: signal is true;
	signal I18960: std_logic; attribute dont_touch of I18960: signal is true;
	signal I18961: std_logic; attribute dont_touch of I18961: signal is true;
	signal I18962: std_logic; attribute dont_touch of I18962: signal is true;
	signal I18967: std_logic; attribute dont_touch of I18967: signal is true;
	signal I18968: std_logic; attribute dont_touch of I18968: signal is true;
	signal I18969: std_logic; attribute dont_touch of I18969: signal is true;
	signal I18970: std_logic; attribute dont_touch of I18970: signal is true;
	signal I18971: std_logic; attribute dont_touch of I18971: signal is true;
	signal I18976: std_logic; attribute dont_touch of I18976: signal is true;
	signal I18977: std_logic; attribute dont_touch of I18977: signal is true;
	signal I18978: std_logic; attribute dont_touch of I18978: signal is true;
	signal I18983: std_logic; attribute dont_touch of I18983: signal is true;
	signal I18984: std_logic; attribute dont_touch of I18984: signal is true;
	signal I18985: std_logic; attribute dont_touch of I18985: signal is true;
	signal I18986: std_logic; attribute dont_touch of I18986: signal is true;
	signal I18991: std_logic; attribute dont_touch of I18991: signal is true;
	signal I18992: std_logic; attribute dont_touch of I18992: signal is true;
	signal I18993: std_logic; attribute dont_touch of I18993: signal is true;
	signal I19072: std_logic; attribute dont_touch of I19072: signal is true;
	signal I19073: std_logic; attribute dont_touch of I19073: signal is true;
	signal I19074: std_logic; attribute dont_touch of I19074: signal is true;
	signal I19085: std_logic; attribute dont_touch of I19085: signal is true;
	signal I19086: std_logic; attribute dont_touch of I19086: signal is true;
	signal I19087: std_logic; attribute dont_touch of I19087: signal is true;
	signal I19098: std_logic; attribute dont_touch of I19098: signal is true;
	signal I19099: std_logic; attribute dont_touch of I19099: signal is true;
	signal I19100: std_logic; attribute dont_touch of I19100: signal is true;
	signal I19111: std_logic; attribute dont_touch of I19111: signal is true;
	signal I19112: std_logic; attribute dont_touch of I19112: signal is true;
	signal I19113: std_logic; attribute dont_touch of I19113: signal is true;
	signal I19124: std_logic; attribute dont_touch of I19124: signal is true;
	signal I19125: std_logic; attribute dont_touch of I19125: signal is true;
	signal I19126: std_logic; attribute dont_touch of I19126: signal is true;
	signal I19137: std_logic; attribute dont_touch of I19137: signal is true;
	signal I19138: std_logic; attribute dont_touch of I19138: signal is true;
	signal I19139: std_logic; attribute dont_touch of I19139: signal is true;
	signal I19150: std_logic; attribute dont_touch of I19150: signal is true;
	signal I19151: std_logic; attribute dont_touch of I19151: signal is true;
	signal I19152: std_logic; attribute dont_touch of I19152: signal is true;
	signal I19163: std_logic; attribute dont_touch of I19163: signal is true;
	signal I19164: std_logic; attribute dont_touch of I19164: signal is true;
	signal I19165: std_logic; attribute dont_touch of I19165: signal is true;
	signal I19176: std_logic; attribute dont_touch of I19176: signal is true;
	signal I19177: std_logic; attribute dont_touch of I19177: signal is true;
	signal I19178: std_logic; attribute dont_touch of I19178: signal is true;
	signal I19189: std_logic; attribute dont_touch of I19189: signal is true;
	signal I19190: std_logic; attribute dont_touch of I19190: signal is true;
	signal I19191: std_logic; attribute dont_touch of I19191: signal is true;
	signal I19202: std_logic; attribute dont_touch of I19202: signal is true;
	signal I19203: std_logic; attribute dont_touch of I19203: signal is true;
	signal I19204: std_logic; attribute dont_touch of I19204: signal is true;
	signal I19215: std_logic; attribute dont_touch of I19215: signal is true;
	signal I19216: std_logic; attribute dont_touch of I19216: signal is true;
	signal I19217: std_logic; attribute dont_touch of I19217: signal is true;
	signal I19228: std_logic; attribute dont_touch of I19228: signal is true;
	signal I19229: std_logic; attribute dont_touch of I19229: signal is true;
	signal I19230: std_logic; attribute dont_touch of I19230: signal is true;
	signal I19241: std_logic; attribute dont_touch of I19241: signal is true;
	signal I19242: std_logic; attribute dont_touch of I19242: signal is true;
	signal I19243: std_logic; attribute dont_touch of I19243: signal is true;
	signal I19254: std_logic; attribute dont_touch of I19254: signal is true;
	signal I19255: std_logic; attribute dont_touch of I19255: signal is true;
	signal I19256: std_logic; attribute dont_touch of I19256: signal is true;
	signal I19267: std_logic; attribute dont_touch of I19267: signal is true;
	signal I19268: std_logic; attribute dont_touch of I19268: signal is true;
	signal I19269: std_logic; attribute dont_touch of I19269: signal is true;
	signal I19280: std_logic; attribute dont_touch of I19280: signal is true;
	signal I19281: std_logic; attribute dont_touch of I19281: signal is true;
	signal I19282: std_logic; attribute dont_touch of I19282: signal is true;
	signal I19293: std_logic; attribute dont_touch of I19293: signal is true;
	signal I19294: std_logic; attribute dont_touch of I19294: signal is true;
	signal I19295: std_logic; attribute dont_touch of I19295: signal is true;
	signal I19306: std_logic; attribute dont_touch of I19306: signal is true;
	signal I19307: std_logic; attribute dont_touch of I19307: signal is true;
	signal I19308: std_logic; attribute dont_touch of I19308: signal is true;
	signal I19319: std_logic; attribute dont_touch of I19319: signal is true;
	signal I19320: std_logic; attribute dont_touch of I19320: signal is true;
	signal I19321: std_logic; attribute dont_touch of I19321: signal is true;
	signal I19332: std_logic; attribute dont_touch of I19332: signal is true;
	signal I19333: std_logic; attribute dont_touch of I19333: signal is true;
	signal I19334: std_logic; attribute dont_touch of I19334: signal is true;
	signal I19345: std_logic; attribute dont_touch of I19345: signal is true;
	signal I19346: std_logic; attribute dont_touch of I19346: signal is true;
	signal I19347: std_logic; attribute dont_touch of I19347: signal is true;
	signal I19358: std_logic; attribute dont_touch of I19358: signal is true;
	signal I19359: std_logic; attribute dont_touch of I19359: signal is true;
	signal I19360: std_logic; attribute dont_touch of I19360: signal is true;
	signal I19371: std_logic; attribute dont_touch of I19371: signal is true;
	signal I19372: std_logic; attribute dont_touch of I19372: signal is true;
	signal I19373: std_logic; attribute dont_touch of I19373: signal is true;
	signal I19384: std_logic; attribute dont_touch of I19384: signal is true;
	signal I19385: std_logic; attribute dont_touch of I19385: signal is true;
	signal I19386: std_logic; attribute dont_touch of I19386: signal is true;
	signal I19397: std_logic; attribute dont_touch of I19397: signal is true;
	signal I19398: std_logic; attribute dont_touch of I19398: signal is true;
	signal I19399: std_logic; attribute dont_touch of I19399: signal is true;
	signal I19410: std_logic; attribute dont_touch of I19410: signal is true;
	signal I19411: std_logic; attribute dont_touch of I19411: signal is true;
	signal I19412: std_logic; attribute dont_touch of I19412: signal is true;
	signal I19423: std_logic; attribute dont_touch of I19423: signal is true;
	signal I19424: std_logic; attribute dont_touch of I19424: signal is true;
	signal I19425: std_logic; attribute dont_touch of I19425: signal is true;
	signal I19436: std_logic; attribute dont_touch of I19436: signal is true;
	signal I19437: std_logic; attribute dont_touch of I19437: signal is true;
	signal I19438: std_logic; attribute dont_touch of I19438: signal is true;
	signal I19449: std_logic; attribute dont_touch of I19449: signal is true;
	signal I19450: std_logic; attribute dont_touch of I19450: signal is true;
	signal I19451: std_logic; attribute dont_touch of I19451: signal is true;
	signal I19462: std_logic; attribute dont_touch of I19462: signal is true;
	signal I19463: std_logic; attribute dont_touch of I19463: signal is true;
	signal I19464: std_logic; attribute dont_touch of I19464: signal is true;
	signal I19475: std_logic; attribute dont_touch of I19475: signal is true;
	signal I19476: std_logic; attribute dont_touch of I19476: signal is true;
	signal I19477: std_logic; attribute dont_touch of I19477: signal is true;
	signal I19489: std_logic; attribute dont_touch of I19489: signal is true;
	signal I19490: std_logic; attribute dont_touch of I19490: signal is true;
	signal I19491: std_logic; attribute dont_touch of I19491: signal is true;
	signal I19492: std_logic; attribute dont_touch of I19492: signal is true;
	signal I19497: std_logic; attribute dont_touch of I19497: signal is true;
	signal I19498: std_logic; attribute dont_touch of I19498: signal is true;
	signal I19499: std_logic; attribute dont_touch of I19499: signal is true;
	signal I19504: std_logic; attribute dont_touch of I19504: signal is true;
	signal I19505: std_logic; attribute dont_touch of I19505: signal is true;
	signal I19506: std_logic; attribute dont_touch of I19506: signal is true;
	signal I19507: std_logic; attribute dont_touch of I19507: signal is true;
	signal I19512: std_logic; attribute dont_touch of I19512: signal is true;
	signal I19513: std_logic; attribute dont_touch of I19513: signal is true;
	signal I19514: std_logic; attribute dont_touch of I19514: signal is true;
	signal I19519: std_logic; attribute dont_touch of I19519: signal is true;
	signal I19520: std_logic; attribute dont_touch of I19520: signal is true;
	signal I19521: std_logic; attribute dont_touch of I19521: signal is true;
	signal I19522: std_logic; attribute dont_touch of I19522: signal is true;
	signal I19527: std_logic; attribute dont_touch of I19527: signal is true;
	signal I19528: std_logic; attribute dont_touch of I19528: signal is true;
	signal I19529: std_logic; attribute dont_touch of I19529: signal is true;
	signal I19534: std_logic; attribute dont_touch of I19534: signal is true;
	signal I19535: std_logic; attribute dont_touch of I19535: signal is true;
	signal I19536: std_logic; attribute dont_touch of I19536: signal is true;
	signal I19541: std_logic; attribute dont_touch of I19541: signal is true;
	signal I19542: std_logic; attribute dont_touch of I19542: signal is true;
	signal I19543: std_logic; attribute dont_touch of I19543: signal is true;
	signal I19548: std_logic; attribute dont_touch of I19548: signal is true;
	signal I19549: std_logic; attribute dont_touch of I19549: signal is true;
	signal I19550: std_logic; attribute dont_touch of I19550: signal is true;
	signal I19555: std_logic; attribute dont_touch of I19555: signal is true;
	signal I19556: std_logic; attribute dont_touch of I19556: signal is true;
	signal I19557: std_logic; attribute dont_touch of I19557: signal is true;
	signal I19562: std_logic; attribute dont_touch of I19562: signal is true;
	signal I19563: std_logic; attribute dont_touch of I19563: signal is true;
	signal I19564: std_logic; attribute dont_touch of I19564: signal is true;
	signal I19569: std_logic; attribute dont_touch of I19569: signal is true;
	signal I19570: std_logic; attribute dont_touch of I19570: signal is true;
	signal I19571: std_logic; attribute dont_touch of I19571: signal is true;
	signal I19576: std_logic; attribute dont_touch of I19576: signal is true;
	signal I19577: std_logic; attribute dont_touch of I19577: signal is true;
	signal I19578: std_logic; attribute dont_touch of I19578: signal is true;
	signal I19583: std_logic; attribute dont_touch of I19583: signal is true;
	signal I19584: std_logic; attribute dont_touch of I19584: signal is true;
	signal I19585: std_logic; attribute dont_touch of I19585: signal is true;
	signal I19590: std_logic; attribute dont_touch of I19590: signal is true;
	signal I19591: std_logic; attribute dont_touch of I19591: signal is true;
	signal I19592: std_logic; attribute dont_touch of I19592: signal is true;
	signal I19597: std_logic; attribute dont_touch of I19597: signal is true;
	signal I19598: std_logic; attribute dont_touch of I19598: signal is true;
	signal I19599: std_logic; attribute dont_touch of I19599: signal is true;
	signal I19604: std_logic; attribute dont_touch of I19604: signal is true;
	signal I19605: std_logic; attribute dont_touch of I19605: signal is true;
	signal I19606: std_logic; attribute dont_touch of I19606: signal is true;
	signal I19611: std_logic; attribute dont_touch of I19611: signal is true;
	signal I19612: std_logic; attribute dont_touch of I19612: signal is true;
	signal I19613: std_logic; attribute dont_touch of I19613: signal is true;
	signal I19618: std_logic; attribute dont_touch of I19618: signal is true;
	signal I19619: std_logic; attribute dont_touch of I19619: signal is true;
	signal I19620: std_logic; attribute dont_touch of I19620: signal is true;
	signal I19625: std_logic; attribute dont_touch of I19625: signal is true;
	signal I19626: std_logic; attribute dont_touch of I19626: signal is true;
	signal I19627: std_logic; attribute dont_touch of I19627: signal is true;
	signal I19632: std_logic; attribute dont_touch of I19632: signal is true;
	signal I19633: std_logic; attribute dont_touch of I19633: signal is true;
	signal I19634: std_logic; attribute dont_touch of I19634: signal is true;
	signal I19639: std_logic; attribute dont_touch of I19639: signal is true;
	signal I19640: std_logic; attribute dont_touch of I19640: signal is true;
	signal I19641: std_logic; attribute dont_touch of I19641: signal is true;
	signal I19646: std_logic; attribute dont_touch of I19646: signal is true;
	signal I19647: std_logic; attribute dont_touch of I19647: signal is true;
	signal I19648: std_logic; attribute dont_touch of I19648: signal is true;
	signal I19653: std_logic; attribute dont_touch of I19653: signal is true;
	signal I19654: std_logic; attribute dont_touch of I19654: signal is true;
	signal I19655: std_logic; attribute dont_touch of I19655: signal is true;
	signal I19660: std_logic; attribute dont_touch of I19660: signal is true;
	signal I19661: std_logic; attribute dont_touch of I19661: signal is true;
	signal I19662: std_logic; attribute dont_touch of I19662: signal is true;
	signal I19667: std_logic; attribute dont_touch of I19667: signal is true;
	signal I19668: std_logic; attribute dont_touch of I19668: signal is true;
	signal I19669: std_logic; attribute dont_touch of I19669: signal is true;
	signal I19674: std_logic; attribute dont_touch of I19674: signal is true;
	signal I19675: std_logic; attribute dont_touch of I19675: signal is true;
	signal I19676: std_logic; attribute dont_touch of I19676: signal is true;
	signal I19681: std_logic; attribute dont_touch of I19681: signal is true;
	signal I19682: std_logic; attribute dont_touch of I19682: signal is true;
	signal I19683: std_logic; attribute dont_touch of I19683: signal is true;
	signal I19688: std_logic; attribute dont_touch of I19688: signal is true;
	signal I19689: std_logic; attribute dont_touch of I19689: signal is true;
	signal I19690: std_logic; attribute dont_touch of I19690: signal is true;
	signal I19695: std_logic; attribute dont_touch of I19695: signal is true;
	signal I19696: std_logic; attribute dont_touch of I19696: signal is true;
	signal I19697: std_logic; attribute dont_touch of I19697: signal is true;
	signal I19702: std_logic; attribute dont_touch of I19702: signal is true;
	signal I19703: std_logic; attribute dont_touch of I19703: signal is true;
	signal I19704: std_logic; attribute dont_touch of I19704: signal is true;
	signal I19709: std_logic; attribute dont_touch of I19709: signal is true;
	signal I19710: std_logic; attribute dont_touch of I19710: signal is true;
	signal I19711: std_logic; attribute dont_touch of I19711: signal is true;
	signal I19716: std_logic; attribute dont_touch of I19716: signal is true;
	signal I19717: std_logic; attribute dont_touch of I19717: signal is true;
	signal I19718: std_logic; attribute dont_touch of I19718: signal is true;
	signal I19723: std_logic; attribute dont_touch of I19723: signal is true;
	signal I19724: std_logic; attribute dont_touch of I19724: signal is true;
	signal I19725: std_logic; attribute dont_touch of I19725: signal is true;
	signal I19730: std_logic; attribute dont_touch of I19730: signal is true;
	signal I19731: std_logic; attribute dont_touch of I19731: signal is true;
	signal I19732: std_logic; attribute dont_touch of I19732: signal is true;
	signal I22011: std_logic; attribute dont_touch of I22011: signal is true;
	signal I22012: std_logic; attribute dont_touch of I22012: signal is true;
	signal I22013: std_logic; attribute dont_touch of I22013: signal is true;
	signal I22014: std_logic; attribute dont_touch of I22014: signal is true;
	signal I22015: std_logic; attribute dont_touch of I22015: signal is true;
	signal I22020: std_logic; attribute dont_touch of I22020: signal is true;
	signal I22021: std_logic; attribute dont_touch of I22021: signal is true;
	signal I22022: std_logic; attribute dont_touch of I22022: signal is true;
	signal I22027: std_logic; attribute dont_touch of I22027: signal is true;
	signal I22028: std_logic; attribute dont_touch of I22028: signal is true;
	signal I22029: std_logic; attribute dont_touch of I22029: signal is true;
	signal I22030: std_logic; attribute dont_touch of I22030: signal is true;
	signal I22035: std_logic; attribute dont_touch of I22035: signal is true;
	signal I22036: std_logic; attribute dont_touch of I22036: signal is true;
	signal I22037: std_logic; attribute dont_touch of I22037: signal is true;
	signal I22042: std_logic; attribute dont_touch of I22042: signal is true;
	signal I22043: std_logic; attribute dont_touch of I22043: signal is true;
	signal I22044: std_logic; attribute dont_touch of I22044: signal is true;
	signal I22045: std_logic; attribute dont_touch of I22045: signal is true;
	signal I22046: std_logic; attribute dont_touch of I22046: signal is true;
	signal I22051: std_logic; attribute dont_touch of I22051: signal is true;
	signal I22052: std_logic; attribute dont_touch of I22052: signal is true;
	signal I22053: std_logic; attribute dont_touch of I22053: signal is true;
	signal I22058: std_logic; attribute dont_touch of I22058: signal is true;
	signal I22059: std_logic; attribute dont_touch of I22059: signal is true;
	signal I22060: std_logic; attribute dont_touch of I22060: signal is true;
	signal I22061: std_logic; attribute dont_touch of I22061: signal is true;
	signal I22066: std_logic; attribute dont_touch of I22066: signal is true;
	signal I22067: std_logic; attribute dont_touch of I22067: signal is true;
	signal I22068: std_logic; attribute dont_touch of I22068: signal is true;
	signal I22073: std_logic; attribute dont_touch of I22073: signal is true;
	signal I22074: std_logic; attribute dont_touch of I22074: signal is true;
	signal I22075: std_logic; attribute dont_touch of I22075: signal is true;
	signal I22076: std_logic; attribute dont_touch of I22076: signal is true;
	signal I22077: std_logic; attribute dont_touch of I22077: signal is true;
	signal I22082: std_logic; attribute dont_touch of I22082: signal is true;
	signal I22083: std_logic; attribute dont_touch of I22083: signal is true;
	signal I22084: std_logic; attribute dont_touch of I22084: signal is true;
	signal I22089: std_logic; attribute dont_touch of I22089: signal is true;
	signal I22090: std_logic; attribute dont_touch of I22090: signal is true;
	signal I22091: std_logic; attribute dont_touch of I22091: signal is true;
	signal I22092: std_logic; attribute dont_touch of I22092: signal is true;
	signal I22097: std_logic; attribute dont_touch of I22097: signal is true;
	signal I22098: std_logic; attribute dont_touch of I22098: signal is true;
	signal I22099: std_logic; attribute dont_touch of I22099: signal is true;
	signal I22104: std_logic; attribute dont_touch of I22104: signal is true;
	signal I22105: std_logic; attribute dont_touch of I22105: signal is true;
	signal I22106: std_logic; attribute dont_touch of I22106: signal is true;
	signal I22107: std_logic; attribute dont_touch of I22107: signal is true;
	signal I22108: std_logic; attribute dont_touch of I22108: signal is true;
	signal I22113: std_logic; attribute dont_touch of I22113: signal is true;
	signal I22114: std_logic; attribute dont_touch of I22114: signal is true;
	signal I22115: std_logic; attribute dont_touch of I22115: signal is true;
	signal I22120: std_logic; attribute dont_touch of I22120: signal is true;
	signal I22121: std_logic; attribute dont_touch of I22121: signal is true;
	signal I22122: std_logic; attribute dont_touch of I22122: signal is true;
	signal I22123: std_logic; attribute dont_touch of I22123: signal is true;
	signal I22128: std_logic; attribute dont_touch of I22128: signal is true;
	signal I22129: std_logic; attribute dont_touch of I22129: signal is true;
	signal I22130: std_logic; attribute dont_touch of I22130: signal is true;
	signal I22135: std_logic; attribute dont_touch of I22135: signal is true;
	signal I22136: std_logic; attribute dont_touch of I22136: signal is true;
	signal I22137: std_logic; attribute dont_touch of I22137: signal is true;
	signal I22138: std_logic; attribute dont_touch of I22138: signal is true;
	signal I22139: std_logic; attribute dont_touch of I22139: signal is true;
	signal I22144: std_logic; attribute dont_touch of I22144: signal is true;
	signal I22145: std_logic; attribute dont_touch of I22145: signal is true;
	signal I22146: std_logic; attribute dont_touch of I22146: signal is true;
	signal I22151: std_logic; attribute dont_touch of I22151: signal is true;
	signal I22152: std_logic; attribute dont_touch of I22152: signal is true;
	signal I22153: std_logic; attribute dont_touch of I22153: signal is true;
	signal I22154: std_logic; attribute dont_touch of I22154: signal is true;
	signal I22159: std_logic; attribute dont_touch of I22159: signal is true;
	signal I22160: std_logic; attribute dont_touch of I22160: signal is true;
	signal I22161: std_logic; attribute dont_touch of I22161: signal is true;
	signal I22166: std_logic; attribute dont_touch of I22166: signal is true;
	signal I22167: std_logic; attribute dont_touch of I22167: signal is true;
	signal I22168: std_logic; attribute dont_touch of I22168: signal is true;
	signal I22169: std_logic; attribute dont_touch of I22169: signal is true;
	signal I22170: std_logic; attribute dont_touch of I22170: signal is true;
	signal I22175: std_logic; attribute dont_touch of I22175: signal is true;
	signal I22176: std_logic; attribute dont_touch of I22176: signal is true;
	signal I22177: std_logic; attribute dont_touch of I22177: signal is true;
	signal I22182: std_logic; attribute dont_touch of I22182: signal is true;
	signal I22183: std_logic; attribute dont_touch of I22183: signal is true;
	signal I22184: std_logic; attribute dont_touch of I22184: signal is true;
	signal I22185: std_logic; attribute dont_touch of I22185: signal is true;
	signal I22190: std_logic; attribute dont_touch of I22190: signal is true;
	signal I22191: std_logic; attribute dont_touch of I22191: signal is true;
	signal I22192: std_logic; attribute dont_touch of I22192: signal is true;
	signal I22197: std_logic; attribute dont_touch of I22197: signal is true;
	signal I22198: std_logic; attribute dont_touch of I22198: signal is true;
	signal I22199: std_logic; attribute dont_touch of I22199: signal is true;
	signal I22200: std_logic; attribute dont_touch of I22200: signal is true;
	signal I22201: std_logic; attribute dont_touch of I22201: signal is true;
	signal I22206: std_logic; attribute dont_touch of I22206: signal is true;
	signal I22207: std_logic; attribute dont_touch of I22207: signal is true;
	signal I22208: std_logic; attribute dont_touch of I22208: signal is true;
	signal I22213: std_logic; attribute dont_touch of I22213: signal is true;
	signal I22214: std_logic; attribute dont_touch of I22214: signal is true;
	signal I22215: std_logic; attribute dont_touch of I22215: signal is true;
	signal I22216: std_logic; attribute dont_touch of I22216: signal is true;
	signal I22221: std_logic; attribute dont_touch of I22221: signal is true;
	signal I22222: std_logic; attribute dont_touch of I22222: signal is true;
	signal I22223: std_logic; attribute dont_touch of I22223: signal is true;
	signal I22228: std_logic; attribute dont_touch of I22228: signal is true;
	signal I22229: std_logic; attribute dont_touch of I22229: signal is true;
	signal I22230: std_logic; attribute dont_touch of I22230: signal is true;
	signal I22231: std_logic; attribute dont_touch of I22231: signal is true;
	signal I22232: std_logic; attribute dont_touch of I22232: signal is true;
	signal I22237: std_logic; attribute dont_touch of I22237: signal is true;
	signal I22238: std_logic; attribute dont_touch of I22238: signal is true;
	signal I22239: std_logic; attribute dont_touch of I22239: signal is true;
	signal I22244: std_logic; attribute dont_touch of I22244: signal is true;
	signal I22245: std_logic; attribute dont_touch of I22245: signal is true;
	signal I22246: std_logic; attribute dont_touch of I22246: signal is true;
	signal I22247: std_logic; attribute dont_touch of I22247: signal is true;
	signal I22252: std_logic; attribute dont_touch of I22252: signal is true;
	signal I22253: std_logic; attribute dont_touch of I22253: signal is true;
	signal I22254: std_logic; attribute dont_touch of I22254: signal is true;
	signal I22259: std_logic; attribute dont_touch of I22259: signal is true;
	signal I22260: std_logic; attribute dont_touch of I22260: signal is true;
	signal I22261: std_logic; attribute dont_touch of I22261: signal is true;
	signal I22262: std_logic; attribute dont_touch of I22262: signal is true;
	signal I22263: std_logic; attribute dont_touch of I22263: signal is true;
	signal I22268: std_logic; attribute dont_touch of I22268: signal is true;
	signal I22269: std_logic; attribute dont_touch of I22269: signal is true;
	signal I22270: std_logic; attribute dont_touch of I22270: signal is true;
	signal I22275: std_logic; attribute dont_touch of I22275: signal is true;
	signal I22276: std_logic; attribute dont_touch of I22276: signal is true;
	signal I22277: std_logic; attribute dont_touch of I22277: signal is true;
	signal I22278: std_logic; attribute dont_touch of I22278: signal is true;
	signal I22283: std_logic; attribute dont_touch of I22283: signal is true;
	signal I22284: std_logic; attribute dont_touch of I22284: signal is true;
	signal I22285: std_logic; attribute dont_touch of I22285: signal is true;
	signal I22290: std_logic; attribute dont_touch of I22290: signal is true;
	signal I22291: std_logic; attribute dont_touch of I22291: signal is true;
	signal I22292: std_logic; attribute dont_touch of I22292: signal is true;
	signal I22293: std_logic; attribute dont_touch of I22293: signal is true;
	signal I22294: std_logic; attribute dont_touch of I22294: signal is true;
	signal I22299: std_logic; attribute dont_touch of I22299: signal is true;
	signal I22300: std_logic; attribute dont_touch of I22300: signal is true;
	signal I22301: std_logic; attribute dont_touch of I22301: signal is true;
	signal I22306: std_logic; attribute dont_touch of I22306: signal is true;
	signal I22307: std_logic; attribute dont_touch of I22307: signal is true;
	signal I22308: std_logic; attribute dont_touch of I22308: signal is true;
	signal I22309: std_logic; attribute dont_touch of I22309: signal is true;
	signal I22314: std_logic; attribute dont_touch of I22314: signal is true;
	signal I22315: std_logic; attribute dont_touch of I22315: signal is true;
	signal I22316: std_logic; attribute dont_touch of I22316: signal is true;
	signal I22321: std_logic; attribute dont_touch of I22321: signal is true;
	signal I22322: std_logic; attribute dont_touch of I22322: signal is true;
	signal I22323: std_logic; attribute dont_touch of I22323: signal is true;
	signal I22324: std_logic; attribute dont_touch of I22324: signal is true;
	signal I22325: std_logic; attribute dont_touch of I22325: signal is true;
	signal I22330: std_logic; attribute dont_touch of I22330: signal is true;
	signal I22331: std_logic; attribute dont_touch of I22331: signal is true;
	signal I22332: std_logic; attribute dont_touch of I22332: signal is true;
	signal I22337: std_logic; attribute dont_touch of I22337: signal is true;
	signal I22338: std_logic; attribute dont_touch of I22338: signal is true;
	signal I22339: std_logic; attribute dont_touch of I22339: signal is true;
	signal I22340: std_logic; attribute dont_touch of I22340: signal is true;
	signal I22345: std_logic; attribute dont_touch of I22345: signal is true;
	signal I22346: std_logic; attribute dont_touch of I22346: signal is true;
	signal I22347: std_logic; attribute dont_touch of I22347: signal is true;
	signal I22352: std_logic; attribute dont_touch of I22352: signal is true;
	signal I22353: std_logic; attribute dont_touch of I22353: signal is true;
	signal I22354: std_logic; attribute dont_touch of I22354: signal is true;
	signal I22355: std_logic; attribute dont_touch of I22355: signal is true;
	signal I22356: std_logic; attribute dont_touch of I22356: signal is true;
	signal I22361: std_logic; attribute dont_touch of I22361: signal is true;
	signal I22362: std_logic; attribute dont_touch of I22362: signal is true;
	signal I22363: std_logic; attribute dont_touch of I22363: signal is true;
	signal I22368: std_logic; attribute dont_touch of I22368: signal is true;
	signal I22369: std_logic; attribute dont_touch of I22369: signal is true;
	signal I22370: std_logic; attribute dont_touch of I22370: signal is true;
	signal I22371: std_logic; attribute dont_touch of I22371: signal is true;
	signal I22376: std_logic; attribute dont_touch of I22376: signal is true;
	signal I22377: std_logic; attribute dont_touch of I22377: signal is true;
	signal I22378: std_logic; attribute dont_touch of I22378: signal is true;
	signal I22383: std_logic; attribute dont_touch of I22383: signal is true;
	signal I22384: std_logic; attribute dont_touch of I22384: signal is true;
	signal I22385: std_logic; attribute dont_touch of I22385: signal is true;
	signal I22386: std_logic; attribute dont_touch of I22386: signal is true;
	signal I22387: std_logic; attribute dont_touch of I22387: signal is true;
	signal I22392: std_logic; attribute dont_touch of I22392: signal is true;
	signal I22393: std_logic; attribute dont_touch of I22393: signal is true;
	signal I22394: std_logic; attribute dont_touch of I22394: signal is true;
	signal I22399: std_logic; attribute dont_touch of I22399: signal is true;
	signal I22400: std_logic; attribute dont_touch of I22400: signal is true;
	signal I22401: std_logic; attribute dont_touch of I22401: signal is true;
	signal I22402: std_logic; attribute dont_touch of I22402: signal is true;
	signal I22407: std_logic; attribute dont_touch of I22407: signal is true;
	signal I22408: std_logic; attribute dont_touch of I22408: signal is true;
	signal I22409: std_logic; attribute dont_touch of I22409: signal is true;
	signal I22414: std_logic; attribute dont_touch of I22414: signal is true;
	signal I22415: std_logic; attribute dont_touch of I22415: signal is true;
	signal I22416: std_logic; attribute dont_touch of I22416: signal is true;
	signal I22417: std_logic; attribute dont_touch of I22417: signal is true;
	signal I22418: std_logic; attribute dont_touch of I22418: signal is true;
	signal I22423: std_logic; attribute dont_touch of I22423: signal is true;
	signal I22424: std_logic; attribute dont_touch of I22424: signal is true;
	signal I22425: std_logic; attribute dont_touch of I22425: signal is true;
	signal I22430: std_logic; attribute dont_touch of I22430: signal is true;
	signal I22431: std_logic; attribute dont_touch of I22431: signal is true;
	signal I22432: std_logic; attribute dont_touch of I22432: signal is true;
	signal I22433: std_logic; attribute dont_touch of I22433: signal is true;
	signal I22438: std_logic; attribute dont_touch of I22438: signal is true;
	signal I22439: std_logic; attribute dont_touch of I22439: signal is true;
	signal I22440: std_logic; attribute dont_touch of I22440: signal is true;
	signal I22445: std_logic; attribute dont_touch of I22445: signal is true;
	signal I22446: std_logic; attribute dont_touch of I22446: signal is true;
	signal I22447: std_logic; attribute dont_touch of I22447: signal is true;
	signal I22448: std_logic; attribute dont_touch of I22448: signal is true;
	signal I22449: std_logic; attribute dont_touch of I22449: signal is true;
	signal I22454: std_logic; attribute dont_touch of I22454: signal is true;
	signal I22455: std_logic; attribute dont_touch of I22455: signal is true;
	signal I22456: std_logic; attribute dont_touch of I22456: signal is true;
	signal I22461: std_logic; attribute dont_touch of I22461: signal is true;
	signal I22462: std_logic; attribute dont_touch of I22462: signal is true;
	signal I22463: std_logic; attribute dont_touch of I22463: signal is true;
	signal I22464: std_logic; attribute dont_touch of I22464: signal is true;
	signal I22469: std_logic; attribute dont_touch of I22469: signal is true;
	signal I22470: std_logic; attribute dont_touch of I22470: signal is true;
	signal I22471: std_logic; attribute dont_touch of I22471: signal is true;
	signal I22476: std_logic; attribute dont_touch of I22476: signal is true;
	signal I22477: std_logic; attribute dont_touch of I22477: signal is true;
	signal I22478: std_logic; attribute dont_touch of I22478: signal is true;
	signal I22479: std_logic; attribute dont_touch of I22479: signal is true;
	signal I22480: std_logic; attribute dont_touch of I22480: signal is true;
	signal I22485: std_logic; attribute dont_touch of I22485: signal is true;
	signal I22486: std_logic; attribute dont_touch of I22486: signal is true;
	signal I22487: std_logic; attribute dont_touch of I22487: signal is true;
	signal I22492: std_logic; attribute dont_touch of I22492: signal is true;
	signal I22493: std_logic; attribute dont_touch of I22493: signal is true;
	signal I22494: std_logic; attribute dont_touch of I22494: signal is true;
	signal I22495: std_logic; attribute dont_touch of I22495: signal is true;
	signal I22500: std_logic; attribute dont_touch of I22500: signal is true;
	signal I22501: std_logic; attribute dont_touch of I22501: signal is true;
	signal I22502: std_logic; attribute dont_touch of I22502: signal is true;
	signal I22507: std_logic; attribute dont_touch of I22507: signal is true;
	signal I22508: std_logic; attribute dont_touch of I22508: signal is true;
	signal I22509: std_logic; attribute dont_touch of I22509: signal is true;
	signal I22510: std_logic; attribute dont_touch of I22510: signal is true;
	signal I22511: std_logic; attribute dont_touch of I22511: signal is true;
	signal I22516: std_logic; attribute dont_touch of I22516: signal is true;
	signal I22517: std_logic; attribute dont_touch of I22517: signal is true;
	signal I22518: std_logic; attribute dont_touch of I22518: signal is true;
	signal I22523: std_logic; attribute dont_touch of I22523: signal is true;
	signal I22524: std_logic; attribute dont_touch of I22524: signal is true;
	signal I22525: std_logic; attribute dont_touch of I22525: signal is true;
	signal I22526: std_logic; attribute dont_touch of I22526: signal is true;
	signal I22531: std_logic; attribute dont_touch of I22531: signal is true;
	signal I22532: std_logic; attribute dont_touch of I22532: signal is true;
	signal I22533: std_logic; attribute dont_touch of I22533: signal is true;
	signal I22538: std_logic; attribute dont_touch of I22538: signal is true;
	signal I22539: std_logic; attribute dont_touch of I22539: signal is true;
	signal I22540: std_logic; attribute dont_touch of I22540: signal is true;
	signal I22541: std_logic; attribute dont_touch of I22541: signal is true;
	signal I22542: std_logic; attribute dont_touch of I22542: signal is true;
	signal I22547: std_logic; attribute dont_touch of I22547: signal is true;
	signal I22548: std_logic; attribute dont_touch of I22548: signal is true;
	signal I22549: std_logic; attribute dont_touch of I22549: signal is true;
	signal I22554: std_logic; attribute dont_touch of I22554: signal is true;
	signal I22555: std_logic; attribute dont_touch of I22555: signal is true;
	signal I22556: std_logic; attribute dont_touch of I22556: signal is true;
	signal I22557: std_logic; attribute dont_touch of I22557: signal is true;
	signal I22562: std_logic; attribute dont_touch of I22562: signal is true;
	signal I22563: std_logic; attribute dont_touch of I22563: signal is true;
	signal I22564: std_logic; attribute dont_touch of I22564: signal is true;
	signal I22569: std_logic; attribute dont_touch of I22569: signal is true;
	signal I22570: std_logic; attribute dont_touch of I22570: signal is true;
	signal I22571: std_logic; attribute dont_touch of I22571: signal is true;
	signal I22572: std_logic; attribute dont_touch of I22572: signal is true;
	signal I22573: std_logic; attribute dont_touch of I22573: signal is true;
	signal I22578: std_logic; attribute dont_touch of I22578: signal is true;
	signal I22579: std_logic; attribute dont_touch of I22579: signal is true;
	signal I22580: std_logic; attribute dont_touch of I22580: signal is true;
	signal I22585: std_logic; attribute dont_touch of I22585: signal is true;
	signal I22586: std_logic; attribute dont_touch of I22586: signal is true;
	signal I22587: std_logic; attribute dont_touch of I22587: signal is true;
	signal I22588: std_logic; attribute dont_touch of I22588: signal is true;
	signal I22593: std_logic; attribute dont_touch of I22593: signal is true;
	signal I22594: std_logic; attribute dont_touch of I22594: signal is true;
	signal I22595: std_logic; attribute dont_touch of I22595: signal is true;
	signal I22600: std_logic; attribute dont_touch of I22600: signal is true;
	signal I22601: std_logic; attribute dont_touch of I22601: signal is true;
	signal I22602: std_logic; attribute dont_touch of I22602: signal is true;
	signal I22603: std_logic; attribute dont_touch of I22603: signal is true;
	signal I22604: std_logic; attribute dont_touch of I22604: signal is true;
	signal I22609: std_logic; attribute dont_touch of I22609: signal is true;
	signal I22610: std_logic; attribute dont_touch of I22610: signal is true;
	signal I22611: std_logic; attribute dont_touch of I22611: signal is true;
	signal I22616: std_logic; attribute dont_touch of I22616: signal is true;
	signal I22617: std_logic; attribute dont_touch of I22617: signal is true;
	signal I22618: std_logic; attribute dont_touch of I22618: signal is true;
	signal I22619: std_logic; attribute dont_touch of I22619: signal is true;
	signal I22624: std_logic; attribute dont_touch of I22624: signal is true;
	signal I22625: std_logic; attribute dont_touch of I22625: signal is true;
	signal I22626: std_logic; attribute dont_touch of I22626: signal is true;
	signal I22631: std_logic; attribute dont_touch of I22631: signal is true;
	signal I22632: std_logic; attribute dont_touch of I22632: signal is true;
	signal I22633: std_logic; attribute dont_touch of I22633: signal is true;
	signal I22634: std_logic; attribute dont_touch of I22634: signal is true;
	signal I22635: std_logic; attribute dont_touch of I22635: signal is true;
	signal I22640: std_logic; attribute dont_touch of I22640: signal is true;
	signal I22641: std_logic; attribute dont_touch of I22641: signal is true;
	signal I22642: std_logic; attribute dont_touch of I22642: signal is true;
	signal I22647: std_logic; attribute dont_touch of I22647: signal is true;
	signal I22648: std_logic; attribute dont_touch of I22648: signal is true;
	signal I22649: std_logic; attribute dont_touch of I22649: signal is true;
	signal I22650: std_logic; attribute dont_touch of I22650: signal is true;
	signal I22655: std_logic; attribute dont_touch of I22655: signal is true;
	signal I22656: std_logic; attribute dont_touch of I22656: signal is true;
	signal I22657: std_logic; attribute dont_touch of I22657: signal is true;
	signal I22662: std_logic; attribute dont_touch of I22662: signal is true;
	signal I22663: std_logic; attribute dont_touch of I22663: signal is true;
	signal I22664: std_logic; attribute dont_touch of I22664: signal is true;
	signal I22665: std_logic; attribute dont_touch of I22665: signal is true;
	signal I22666: std_logic; attribute dont_touch of I22666: signal is true;
	signal I22671: std_logic; attribute dont_touch of I22671: signal is true;
	signal I22672: std_logic; attribute dont_touch of I22672: signal is true;
	signal I22673: std_logic; attribute dont_touch of I22673: signal is true;
	signal I22678: std_logic; attribute dont_touch of I22678: signal is true;
	signal I22679: std_logic; attribute dont_touch of I22679: signal is true;
	signal I22680: std_logic; attribute dont_touch of I22680: signal is true;
	signal I22681: std_logic; attribute dont_touch of I22681: signal is true;
	signal I22686: std_logic; attribute dont_touch of I22686: signal is true;
	signal I22687: std_logic; attribute dont_touch of I22687: signal is true;
	signal I22688: std_logic; attribute dont_touch of I22688: signal is true;
	signal I22693: std_logic; attribute dont_touch of I22693: signal is true;
	signal I22694: std_logic; attribute dont_touch of I22694: signal is true;
	signal I22695: std_logic; attribute dont_touch of I22695: signal is true;
	signal I22696: std_logic; attribute dont_touch of I22696: signal is true;
	signal I22697: std_logic; attribute dont_touch of I22697: signal is true;
	signal I22702: std_logic; attribute dont_touch of I22702: signal is true;
	signal I22703: std_logic; attribute dont_touch of I22703: signal is true;
	signal I22704: std_logic; attribute dont_touch of I22704: signal is true;
	signal I22709: std_logic; attribute dont_touch of I22709: signal is true;
	signal I22710: std_logic; attribute dont_touch of I22710: signal is true;
	signal I22711: std_logic; attribute dont_touch of I22711: signal is true;
	signal I22712: std_logic; attribute dont_touch of I22712: signal is true;
	signal I22717: std_logic; attribute dont_touch of I22717: signal is true;
	signal I22718: std_logic; attribute dont_touch of I22718: signal is true;
	signal I22719: std_logic; attribute dont_touch of I22719: signal is true;
	signal I22724: std_logic; attribute dont_touch of I22724: signal is true;
	signal I22725: std_logic; attribute dont_touch of I22725: signal is true;
	signal I22726: std_logic; attribute dont_touch of I22726: signal is true;
	signal I22727: std_logic; attribute dont_touch of I22727: signal is true;
	signal I22728: std_logic; attribute dont_touch of I22728: signal is true;
	signal I22733: std_logic; attribute dont_touch of I22733: signal is true;
	signal I22734: std_logic; attribute dont_touch of I22734: signal is true;
	signal I22735: std_logic; attribute dont_touch of I22735: signal is true;
	signal I22740: std_logic; attribute dont_touch of I22740: signal is true;
	signal I22741: std_logic; attribute dont_touch of I22741: signal is true;
	signal I22742: std_logic; attribute dont_touch of I22742: signal is true;
	signal I22743: std_logic; attribute dont_touch of I22743: signal is true;
	signal I22748: std_logic; attribute dont_touch of I22748: signal is true;
	signal I22749: std_logic; attribute dont_touch of I22749: signal is true;
	signal I22750: std_logic; attribute dont_touch of I22750: signal is true;
	signal I22755: std_logic; attribute dont_touch of I22755: signal is true;
	signal I22756: std_logic; attribute dont_touch of I22756: signal is true;
	signal I22757: std_logic; attribute dont_touch of I22757: signal is true;
	signal I22758: std_logic; attribute dont_touch of I22758: signal is true;
	signal I22759: std_logic; attribute dont_touch of I22759: signal is true;
	signal I22764: std_logic; attribute dont_touch of I22764: signal is true;
	signal I22765: std_logic; attribute dont_touch of I22765: signal is true;
	signal I22766: std_logic; attribute dont_touch of I22766: signal is true;
	signal I22771: std_logic; attribute dont_touch of I22771: signal is true;
	signal I22772: std_logic; attribute dont_touch of I22772: signal is true;
	signal I22773: std_logic; attribute dont_touch of I22773: signal is true;
	signal I22774: std_logic; attribute dont_touch of I22774: signal is true;
	signal I22779: std_logic; attribute dont_touch of I22779: signal is true;
	signal I22780: std_logic; attribute dont_touch of I22780: signal is true;
	signal I22781: std_logic; attribute dont_touch of I22781: signal is true;
	signal I22786: std_logic; attribute dont_touch of I22786: signal is true;
	signal I22787: std_logic; attribute dont_touch of I22787: signal is true;
	signal I22788: std_logic; attribute dont_touch of I22788: signal is true;
	signal I22789: std_logic; attribute dont_touch of I22789: signal is true;
	signal I22790: std_logic; attribute dont_touch of I22790: signal is true;
	signal I22795: std_logic; attribute dont_touch of I22795: signal is true;
	signal I22796: std_logic; attribute dont_touch of I22796: signal is true;
	signal I22797: std_logic; attribute dont_touch of I22797: signal is true;
	signal I22802: std_logic; attribute dont_touch of I22802: signal is true;
	signal I22803: std_logic; attribute dont_touch of I22803: signal is true;
	signal I22804: std_logic; attribute dont_touch of I22804: signal is true;
	signal I22805: std_logic; attribute dont_touch of I22805: signal is true;
	signal I22810: std_logic; attribute dont_touch of I22810: signal is true;
	signal I22811: std_logic; attribute dont_touch of I22811: signal is true;
	signal I22812: std_logic; attribute dont_touch of I22812: signal is true;
	signal I22817: std_logic; attribute dont_touch of I22817: signal is true;
	signal I22818: std_logic; attribute dont_touch of I22818: signal is true;
	signal I22819: std_logic; attribute dont_touch of I22819: signal is true;
	signal I22820: std_logic; attribute dont_touch of I22820: signal is true;
	signal I22821: std_logic; attribute dont_touch of I22821: signal is true;
	signal I22826: std_logic; attribute dont_touch of I22826: signal is true;
	signal I22827: std_logic; attribute dont_touch of I22827: signal is true;
	signal I22828: std_logic; attribute dont_touch of I22828: signal is true;
	signal I22833: std_logic; attribute dont_touch of I22833: signal is true;
	signal I22834: std_logic; attribute dont_touch of I22834: signal is true;
	signal I22835: std_logic; attribute dont_touch of I22835: signal is true;
	signal I22836: std_logic; attribute dont_touch of I22836: signal is true;
	signal I22841: std_logic; attribute dont_touch of I22841: signal is true;
	signal I22842: std_logic; attribute dont_touch of I22842: signal is true;
	signal I22843: std_logic; attribute dont_touch of I22843: signal is true;
	signal I22848: std_logic; attribute dont_touch of I22848: signal is true;
	signal I22849: std_logic; attribute dont_touch of I22849: signal is true;
	signal I22850: std_logic; attribute dont_touch of I22850: signal is true;
	signal I22851: std_logic; attribute dont_touch of I22851: signal is true;
	signal I22852: std_logic; attribute dont_touch of I22852: signal is true;
	signal I22857: std_logic; attribute dont_touch of I22857: signal is true;
	signal I22858: std_logic; attribute dont_touch of I22858: signal is true;
	signal I22859: std_logic; attribute dont_touch of I22859: signal is true;
	signal I22864: std_logic; attribute dont_touch of I22864: signal is true;
	signal I22865: std_logic; attribute dont_touch of I22865: signal is true;
	signal I22866: std_logic; attribute dont_touch of I22866: signal is true;
	signal I22867: std_logic; attribute dont_touch of I22867: signal is true;
	signal I22872: std_logic; attribute dont_touch of I22872: signal is true;
	signal I22873: std_logic; attribute dont_touch of I22873: signal is true;
	signal I22874: std_logic; attribute dont_touch of I22874: signal is true;
	signal I22879: std_logic; attribute dont_touch of I22879: signal is true;
	signal I22880: std_logic; attribute dont_touch of I22880: signal is true;
	signal I22881: std_logic; attribute dont_touch of I22881: signal is true;
	signal I22882: std_logic; attribute dont_touch of I22882: signal is true;
	signal I22883: std_logic; attribute dont_touch of I22883: signal is true;
	signal I22888: std_logic; attribute dont_touch of I22888: signal is true;
	signal I22889: std_logic; attribute dont_touch of I22889: signal is true;
	signal I22890: std_logic; attribute dont_touch of I22890: signal is true;
	signal I22895: std_logic; attribute dont_touch of I22895: signal is true;
	signal I22896: std_logic; attribute dont_touch of I22896: signal is true;
	signal I22897: std_logic; attribute dont_touch of I22897: signal is true;
	signal I22898: std_logic; attribute dont_touch of I22898: signal is true;
	signal I22903: std_logic; attribute dont_touch of I22903: signal is true;
	signal I22904: std_logic; attribute dont_touch of I22904: signal is true;
	signal I22905: std_logic; attribute dont_touch of I22905: signal is true;
	signal I22910: std_logic; attribute dont_touch of I22910: signal is true;
	signal I22911: std_logic; attribute dont_touch of I22911: signal is true;
	signal I22912: std_logic; attribute dont_touch of I22912: signal is true;
	signal I22913: std_logic; attribute dont_touch of I22913: signal is true;
	signal I22914: std_logic; attribute dont_touch of I22914: signal is true;
	signal I22919: std_logic; attribute dont_touch of I22919: signal is true;
	signal I22920: std_logic; attribute dont_touch of I22920: signal is true;
	signal I22921: std_logic; attribute dont_touch of I22921: signal is true;
	signal I22926: std_logic; attribute dont_touch of I22926: signal is true;
	signal I22927: std_logic; attribute dont_touch of I22927: signal is true;
	signal I22928: std_logic; attribute dont_touch of I22928: signal is true;
	signal I22929: std_logic; attribute dont_touch of I22929: signal is true;
	signal I22934: std_logic; attribute dont_touch of I22934: signal is true;
	signal I22935: std_logic; attribute dont_touch of I22935: signal is true;
	signal I22936: std_logic; attribute dont_touch of I22936: signal is true;
	signal I22941: std_logic; attribute dont_touch of I22941: signal is true;
	signal I22942: std_logic; attribute dont_touch of I22942: signal is true;
	signal I22943: std_logic; attribute dont_touch of I22943: signal is true;
	signal I22944: std_logic; attribute dont_touch of I22944: signal is true;
	signal I22945: std_logic; attribute dont_touch of I22945: signal is true;
	signal I22950: std_logic; attribute dont_touch of I22950: signal is true;
	signal I22951: std_logic; attribute dont_touch of I22951: signal is true;
	signal I22952: std_logic; attribute dont_touch of I22952: signal is true;
	signal I22957: std_logic; attribute dont_touch of I22957: signal is true;
	signal I22958: std_logic; attribute dont_touch of I22958: signal is true;
	signal I22959: std_logic; attribute dont_touch of I22959: signal is true;
	signal I22960: std_logic; attribute dont_touch of I22960: signal is true;
	signal I22965: std_logic; attribute dont_touch of I22965: signal is true;
	signal I22966: std_logic; attribute dont_touch of I22966: signal is true;
	signal I22967: std_logic; attribute dont_touch of I22967: signal is true;
	signal I22972: std_logic; attribute dont_touch of I22972: signal is true;
	signal I22973: std_logic; attribute dont_touch of I22973: signal is true;
	signal I22974: std_logic; attribute dont_touch of I22974: signal is true;
	signal I22975: std_logic; attribute dont_touch of I22975: signal is true;
	signal I22976: std_logic; attribute dont_touch of I22976: signal is true;
	signal I22981: std_logic; attribute dont_touch of I22981: signal is true;
	signal I22982: std_logic; attribute dont_touch of I22982: signal is true;
	signal I22983: std_logic; attribute dont_touch of I22983: signal is true;
	signal I22988: std_logic; attribute dont_touch of I22988: signal is true;
	signal I22989: std_logic; attribute dont_touch of I22989: signal is true;
	signal I22990: std_logic; attribute dont_touch of I22990: signal is true;
	signal I22991: std_logic; attribute dont_touch of I22991: signal is true;
	signal I22996: std_logic; attribute dont_touch of I22996: signal is true;
	signal I22997: std_logic; attribute dont_touch of I22997: signal is true;
	signal I22998: std_logic; attribute dont_touch of I22998: signal is true;
	signal I23077: std_logic; attribute dont_touch of I23077: signal is true;
	signal I23078: std_logic; attribute dont_touch of I23078: signal is true;
	signal I23079: std_logic; attribute dont_touch of I23079: signal is true;
	signal I23090: std_logic; attribute dont_touch of I23090: signal is true;
	signal I23091: std_logic; attribute dont_touch of I23091: signal is true;
	signal I23092: std_logic; attribute dont_touch of I23092: signal is true;
	signal I23103: std_logic; attribute dont_touch of I23103: signal is true;
	signal I23104: std_logic; attribute dont_touch of I23104: signal is true;
	signal I23105: std_logic; attribute dont_touch of I23105: signal is true;
	signal I23116: std_logic; attribute dont_touch of I23116: signal is true;
	signal I23117: std_logic; attribute dont_touch of I23117: signal is true;
	signal I23118: std_logic; attribute dont_touch of I23118: signal is true;
	signal I23129: std_logic; attribute dont_touch of I23129: signal is true;
	signal I23130: std_logic; attribute dont_touch of I23130: signal is true;
	signal I23131: std_logic; attribute dont_touch of I23131: signal is true;
	signal I23142: std_logic; attribute dont_touch of I23142: signal is true;
	signal I23143: std_logic; attribute dont_touch of I23143: signal is true;
	signal I23144: std_logic; attribute dont_touch of I23144: signal is true;
	signal I23155: std_logic; attribute dont_touch of I23155: signal is true;
	signal I23156: std_logic; attribute dont_touch of I23156: signal is true;
	signal I23157: std_logic; attribute dont_touch of I23157: signal is true;
	signal I23168: std_logic; attribute dont_touch of I23168: signal is true;
	signal I23169: std_logic; attribute dont_touch of I23169: signal is true;
	signal I23170: std_logic; attribute dont_touch of I23170: signal is true;
	signal I23181: std_logic; attribute dont_touch of I23181: signal is true;
	signal I23182: std_logic; attribute dont_touch of I23182: signal is true;
	signal I23183: std_logic; attribute dont_touch of I23183: signal is true;
	signal I23194: std_logic; attribute dont_touch of I23194: signal is true;
	signal I23195: std_logic; attribute dont_touch of I23195: signal is true;
	signal I23196: std_logic; attribute dont_touch of I23196: signal is true;
	signal I23207: std_logic; attribute dont_touch of I23207: signal is true;
	signal I23208: std_logic; attribute dont_touch of I23208: signal is true;
	signal I23209: std_logic; attribute dont_touch of I23209: signal is true;
	signal I23220: std_logic; attribute dont_touch of I23220: signal is true;
	signal I23221: std_logic; attribute dont_touch of I23221: signal is true;
	signal I23222: std_logic; attribute dont_touch of I23222: signal is true;
	signal I23233: std_logic; attribute dont_touch of I23233: signal is true;
	signal I23234: std_logic; attribute dont_touch of I23234: signal is true;
	signal I23235: std_logic; attribute dont_touch of I23235: signal is true;
	signal I23246: std_logic; attribute dont_touch of I23246: signal is true;
	signal I23247: std_logic; attribute dont_touch of I23247: signal is true;
	signal I23248: std_logic; attribute dont_touch of I23248: signal is true;
	signal I23259: std_logic; attribute dont_touch of I23259: signal is true;
	signal I23260: std_logic; attribute dont_touch of I23260: signal is true;
	signal I23261: std_logic; attribute dont_touch of I23261: signal is true;
	signal I23272: std_logic; attribute dont_touch of I23272: signal is true;
	signal I23273: std_logic; attribute dont_touch of I23273: signal is true;
	signal I23274: std_logic; attribute dont_touch of I23274: signal is true;
	signal I23285: std_logic; attribute dont_touch of I23285: signal is true;
	signal I23286: std_logic; attribute dont_touch of I23286: signal is true;
	signal I23287: std_logic; attribute dont_touch of I23287: signal is true;
	signal I23298: std_logic; attribute dont_touch of I23298: signal is true;
	signal I23299: std_logic; attribute dont_touch of I23299: signal is true;
	signal I23300: std_logic; attribute dont_touch of I23300: signal is true;
	signal I23311: std_logic; attribute dont_touch of I23311: signal is true;
	signal I23312: std_logic; attribute dont_touch of I23312: signal is true;
	signal I23313: std_logic; attribute dont_touch of I23313: signal is true;
	signal I23324: std_logic; attribute dont_touch of I23324: signal is true;
	signal I23325: std_logic; attribute dont_touch of I23325: signal is true;
	signal I23326: std_logic; attribute dont_touch of I23326: signal is true;
	signal I23337: std_logic; attribute dont_touch of I23337: signal is true;
	signal I23338: std_logic; attribute dont_touch of I23338: signal is true;
	signal I23339: std_logic; attribute dont_touch of I23339: signal is true;
	signal I23350: std_logic; attribute dont_touch of I23350: signal is true;
	signal I23351: std_logic; attribute dont_touch of I23351: signal is true;
	signal I23352: std_logic; attribute dont_touch of I23352: signal is true;
	signal I23363: std_logic; attribute dont_touch of I23363: signal is true;
	signal I23364: std_logic; attribute dont_touch of I23364: signal is true;
	signal I23365: std_logic; attribute dont_touch of I23365: signal is true;
	signal I23376: std_logic; attribute dont_touch of I23376: signal is true;
	signal I23377: std_logic; attribute dont_touch of I23377: signal is true;
	signal I23378: std_logic; attribute dont_touch of I23378: signal is true;
	signal I23389: std_logic; attribute dont_touch of I23389: signal is true;
	signal I23390: std_logic; attribute dont_touch of I23390: signal is true;
	signal I23391: std_logic; attribute dont_touch of I23391: signal is true;
	signal I23402: std_logic; attribute dont_touch of I23402: signal is true;
	signal I23403: std_logic; attribute dont_touch of I23403: signal is true;
	signal I23404: std_logic; attribute dont_touch of I23404: signal is true;
	signal I23415: std_logic; attribute dont_touch of I23415: signal is true;
	signal I23416: std_logic; attribute dont_touch of I23416: signal is true;
	signal I23417: std_logic; attribute dont_touch of I23417: signal is true;
	signal I23428: std_logic; attribute dont_touch of I23428: signal is true;
	signal I23429: std_logic; attribute dont_touch of I23429: signal is true;
	signal I23430: std_logic; attribute dont_touch of I23430: signal is true;
	signal I23441: std_logic; attribute dont_touch of I23441: signal is true;
	signal I23442: std_logic; attribute dont_touch of I23442: signal is true;
	signal I23443: std_logic; attribute dont_touch of I23443: signal is true;
	signal I23454: std_logic; attribute dont_touch of I23454: signal is true;
	signal I23455: std_logic; attribute dont_touch of I23455: signal is true;
	signal I23456: std_logic; attribute dont_touch of I23456: signal is true;
	signal I23467: std_logic; attribute dont_touch of I23467: signal is true;
	signal I23468: std_logic; attribute dont_touch of I23468: signal is true;
	signal I23469: std_logic; attribute dont_touch of I23469: signal is true;
	signal I23480: std_logic; attribute dont_touch of I23480: signal is true;
	signal I23481: std_logic; attribute dont_touch of I23481: signal is true;
	signal I23482: std_logic; attribute dont_touch of I23482: signal is true;
	signal I23494: std_logic; attribute dont_touch of I23494: signal is true;
	signal I23495: std_logic; attribute dont_touch of I23495: signal is true;
	signal I23496: std_logic; attribute dont_touch of I23496: signal is true;
	signal I23497: std_logic; attribute dont_touch of I23497: signal is true;
	signal I23502: std_logic; attribute dont_touch of I23502: signal is true;
	signal I23503: std_logic; attribute dont_touch of I23503: signal is true;
	signal I23504: std_logic; attribute dont_touch of I23504: signal is true;
	signal I23509: std_logic; attribute dont_touch of I23509: signal is true;
	signal I23510: std_logic; attribute dont_touch of I23510: signal is true;
	signal I23511: std_logic; attribute dont_touch of I23511: signal is true;
	signal I23512: std_logic; attribute dont_touch of I23512: signal is true;
	signal I23517: std_logic; attribute dont_touch of I23517: signal is true;
	signal I23518: std_logic; attribute dont_touch of I23518: signal is true;
	signal I23519: std_logic; attribute dont_touch of I23519: signal is true;
	signal I23524: std_logic; attribute dont_touch of I23524: signal is true;
	signal I23525: std_logic; attribute dont_touch of I23525: signal is true;
	signal I23526: std_logic; attribute dont_touch of I23526: signal is true;
	signal I23527: std_logic; attribute dont_touch of I23527: signal is true;
	signal I23532: std_logic; attribute dont_touch of I23532: signal is true;
	signal I23533: std_logic; attribute dont_touch of I23533: signal is true;
	signal I23534: std_logic; attribute dont_touch of I23534: signal is true;
	signal I23539: std_logic; attribute dont_touch of I23539: signal is true;
	signal I23540: std_logic; attribute dont_touch of I23540: signal is true;
	signal I23541: std_logic; attribute dont_touch of I23541: signal is true;
	signal I23546: std_logic; attribute dont_touch of I23546: signal is true;
	signal I23547: std_logic; attribute dont_touch of I23547: signal is true;
	signal I23548: std_logic; attribute dont_touch of I23548: signal is true;
	signal I23553: std_logic; attribute dont_touch of I23553: signal is true;
	signal I23554: std_logic; attribute dont_touch of I23554: signal is true;
	signal I23555: std_logic; attribute dont_touch of I23555: signal is true;
	signal I23560: std_logic; attribute dont_touch of I23560: signal is true;
	signal I23561: std_logic; attribute dont_touch of I23561: signal is true;
	signal I23562: std_logic; attribute dont_touch of I23562: signal is true;
	signal I23567: std_logic; attribute dont_touch of I23567: signal is true;
	signal I23568: std_logic; attribute dont_touch of I23568: signal is true;
	signal I23569: std_logic; attribute dont_touch of I23569: signal is true;
	signal I23574: std_logic; attribute dont_touch of I23574: signal is true;
	signal I23575: std_logic; attribute dont_touch of I23575: signal is true;
	signal I23576: std_logic; attribute dont_touch of I23576: signal is true;
	signal I23581: std_logic; attribute dont_touch of I23581: signal is true;
	signal I23582: std_logic; attribute dont_touch of I23582: signal is true;
	signal I23583: std_logic; attribute dont_touch of I23583: signal is true;
	signal I23588: std_logic; attribute dont_touch of I23588: signal is true;
	signal I23589: std_logic; attribute dont_touch of I23589: signal is true;
	signal I23590: std_logic; attribute dont_touch of I23590: signal is true;
	signal I23595: std_logic; attribute dont_touch of I23595: signal is true;
	signal I23596: std_logic; attribute dont_touch of I23596: signal is true;
	signal I23597: std_logic; attribute dont_touch of I23597: signal is true;
	signal I23602: std_logic; attribute dont_touch of I23602: signal is true;
	signal I23603: std_logic; attribute dont_touch of I23603: signal is true;
	signal I23604: std_logic; attribute dont_touch of I23604: signal is true;
	signal I23609: std_logic; attribute dont_touch of I23609: signal is true;
	signal I23610: std_logic; attribute dont_touch of I23610: signal is true;
	signal I23611: std_logic; attribute dont_touch of I23611: signal is true;
	signal I23616: std_logic; attribute dont_touch of I23616: signal is true;
	signal I23617: std_logic; attribute dont_touch of I23617: signal is true;
	signal I23618: std_logic; attribute dont_touch of I23618: signal is true;
	signal I23623: std_logic; attribute dont_touch of I23623: signal is true;
	signal I23624: std_logic; attribute dont_touch of I23624: signal is true;
	signal I23625: std_logic; attribute dont_touch of I23625: signal is true;
	signal I23630: std_logic; attribute dont_touch of I23630: signal is true;
	signal I23631: std_logic; attribute dont_touch of I23631: signal is true;
	signal I23632: std_logic; attribute dont_touch of I23632: signal is true;
	signal I23637: std_logic; attribute dont_touch of I23637: signal is true;
	signal I23638: std_logic; attribute dont_touch of I23638: signal is true;
	signal I23639: std_logic; attribute dont_touch of I23639: signal is true;
	signal I23644: std_logic; attribute dont_touch of I23644: signal is true;
	signal I23645: std_logic; attribute dont_touch of I23645: signal is true;
	signal I23646: std_logic; attribute dont_touch of I23646: signal is true;
	signal I23651: std_logic; attribute dont_touch of I23651: signal is true;
	signal I23652: std_logic; attribute dont_touch of I23652: signal is true;
	signal I23653: std_logic; attribute dont_touch of I23653: signal is true;
	signal I23658: std_logic; attribute dont_touch of I23658: signal is true;
	signal I23659: std_logic; attribute dont_touch of I23659: signal is true;
	signal I23660: std_logic; attribute dont_touch of I23660: signal is true;
	signal I23665: std_logic; attribute dont_touch of I23665: signal is true;
	signal I23666: std_logic; attribute dont_touch of I23666: signal is true;
	signal I23667: std_logic; attribute dont_touch of I23667: signal is true;
	signal I23672: std_logic; attribute dont_touch of I23672: signal is true;
	signal I23673: std_logic; attribute dont_touch of I23673: signal is true;
	signal I23674: std_logic; attribute dont_touch of I23674: signal is true;
	signal I23679: std_logic; attribute dont_touch of I23679: signal is true;
	signal I23680: std_logic; attribute dont_touch of I23680: signal is true;
	signal I23681: std_logic; attribute dont_touch of I23681: signal is true;
	signal I23686: std_logic; attribute dont_touch of I23686: signal is true;
	signal I23687: std_logic; attribute dont_touch of I23687: signal is true;
	signal I23688: std_logic; attribute dont_touch of I23688: signal is true;
	signal I23693: std_logic; attribute dont_touch of I23693: signal is true;
	signal I23694: std_logic; attribute dont_touch of I23694: signal is true;
	signal I23695: std_logic; attribute dont_touch of I23695: signal is true;
	signal I23700: std_logic; attribute dont_touch of I23700: signal is true;
	signal I23701: std_logic; attribute dont_touch of I23701: signal is true;
	signal I23702: std_logic; attribute dont_touch of I23702: signal is true;
	signal I23707: std_logic; attribute dont_touch of I23707: signal is true;
	signal I23708: std_logic; attribute dont_touch of I23708: signal is true;
	signal I23709: std_logic; attribute dont_touch of I23709: signal is true;
	signal I23714: std_logic; attribute dont_touch of I23714: signal is true;
	signal I23715: std_logic; attribute dont_touch of I23715: signal is true;
	signal I23716: std_logic; attribute dont_touch of I23716: signal is true;
	signal I23721: std_logic; attribute dont_touch of I23721: signal is true;
	signal I23722: std_logic; attribute dont_touch of I23722: signal is true;
	signal I23723: std_logic; attribute dont_touch of I23723: signal is true;
	signal I23728: std_logic; attribute dont_touch of I23728: signal is true;
	signal I23729: std_logic; attribute dont_touch of I23729: signal is true;
	signal I23730: std_logic; attribute dont_touch of I23730: signal is true;
	signal I23735: std_logic; attribute dont_touch of I23735: signal is true;
	signal I23736: std_logic; attribute dont_touch of I23736: signal is true;
	signal I23737: std_logic; attribute dont_touch of I23737: signal is true;
	signal I26016: std_logic; attribute dont_touch of I26016: signal is true;
	signal I26017: std_logic; attribute dont_touch of I26017: signal is true;
	signal I26018: std_logic; attribute dont_touch of I26018: signal is true;
	signal I26019: std_logic; attribute dont_touch of I26019: signal is true;
	signal I26020: std_logic; attribute dont_touch of I26020: signal is true;
	signal I26025: std_logic; attribute dont_touch of I26025: signal is true;
	signal I26026: std_logic; attribute dont_touch of I26026: signal is true;
	signal I26027: std_logic; attribute dont_touch of I26027: signal is true;
	signal I26032: std_logic; attribute dont_touch of I26032: signal is true;
	signal I26033: std_logic; attribute dont_touch of I26033: signal is true;
	signal I26034: std_logic; attribute dont_touch of I26034: signal is true;
	signal I26035: std_logic; attribute dont_touch of I26035: signal is true;
	signal I26040: std_logic; attribute dont_touch of I26040: signal is true;
	signal I26041: std_logic; attribute dont_touch of I26041: signal is true;
	signal I26042: std_logic; attribute dont_touch of I26042: signal is true;
	signal I26047: std_logic; attribute dont_touch of I26047: signal is true;
	signal I26048: std_logic; attribute dont_touch of I26048: signal is true;
	signal I26049: std_logic; attribute dont_touch of I26049: signal is true;
	signal I26050: std_logic; attribute dont_touch of I26050: signal is true;
	signal I26051: std_logic; attribute dont_touch of I26051: signal is true;
	signal I26056: std_logic; attribute dont_touch of I26056: signal is true;
	signal I26057: std_logic; attribute dont_touch of I26057: signal is true;
	signal I26058: std_logic; attribute dont_touch of I26058: signal is true;
	signal I26063: std_logic; attribute dont_touch of I26063: signal is true;
	signal I26064: std_logic; attribute dont_touch of I26064: signal is true;
	signal I26065: std_logic; attribute dont_touch of I26065: signal is true;
	signal I26066: std_logic; attribute dont_touch of I26066: signal is true;
	signal I26071: std_logic; attribute dont_touch of I26071: signal is true;
	signal I26072: std_logic; attribute dont_touch of I26072: signal is true;
	signal I26073: std_logic; attribute dont_touch of I26073: signal is true;
	signal I26078: std_logic; attribute dont_touch of I26078: signal is true;
	signal I26079: std_logic; attribute dont_touch of I26079: signal is true;
	signal I26080: std_logic; attribute dont_touch of I26080: signal is true;
	signal I26081: std_logic; attribute dont_touch of I26081: signal is true;
	signal I26082: std_logic; attribute dont_touch of I26082: signal is true;
	signal I26087: std_logic; attribute dont_touch of I26087: signal is true;
	signal I26088: std_logic; attribute dont_touch of I26088: signal is true;
	signal I26089: std_logic; attribute dont_touch of I26089: signal is true;
	signal I26094: std_logic; attribute dont_touch of I26094: signal is true;
	signal I26095: std_logic; attribute dont_touch of I26095: signal is true;
	signal I26096: std_logic; attribute dont_touch of I26096: signal is true;
	signal I26097: std_logic; attribute dont_touch of I26097: signal is true;
	signal I26102: std_logic; attribute dont_touch of I26102: signal is true;
	signal I26103: std_logic; attribute dont_touch of I26103: signal is true;
	signal I26104: std_logic; attribute dont_touch of I26104: signal is true;
	signal I26109: std_logic; attribute dont_touch of I26109: signal is true;
	signal I26110: std_logic; attribute dont_touch of I26110: signal is true;
	signal I26111: std_logic; attribute dont_touch of I26111: signal is true;
	signal I26112: std_logic; attribute dont_touch of I26112: signal is true;
	signal I26113: std_logic; attribute dont_touch of I26113: signal is true;
	signal I26118: std_logic; attribute dont_touch of I26118: signal is true;
	signal I26119: std_logic; attribute dont_touch of I26119: signal is true;
	signal I26120: std_logic; attribute dont_touch of I26120: signal is true;
	signal I26125: std_logic; attribute dont_touch of I26125: signal is true;
	signal I26126: std_logic; attribute dont_touch of I26126: signal is true;
	signal I26127: std_logic; attribute dont_touch of I26127: signal is true;
	signal I26128: std_logic; attribute dont_touch of I26128: signal is true;
	signal I26133: std_logic; attribute dont_touch of I26133: signal is true;
	signal I26134: std_logic; attribute dont_touch of I26134: signal is true;
	signal I26135: std_logic; attribute dont_touch of I26135: signal is true;
	signal I26140: std_logic; attribute dont_touch of I26140: signal is true;
	signal I26141: std_logic; attribute dont_touch of I26141: signal is true;
	signal I26142: std_logic; attribute dont_touch of I26142: signal is true;
	signal I26143: std_logic; attribute dont_touch of I26143: signal is true;
	signal I26144: std_logic; attribute dont_touch of I26144: signal is true;
	signal I26149: std_logic; attribute dont_touch of I26149: signal is true;
	signal I26150: std_logic; attribute dont_touch of I26150: signal is true;
	signal I26151: std_logic; attribute dont_touch of I26151: signal is true;
	signal I26156: std_logic; attribute dont_touch of I26156: signal is true;
	signal I26157: std_logic; attribute dont_touch of I26157: signal is true;
	signal I26158: std_logic; attribute dont_touch of I26158: signal is true;
	signal I26159: std_logic; attribute dont_touch of I26159: signal is true;
	signal I26164: std_logic; attribute dont_touch of I26164: signal is true;
	signal I26165: std_logic; attribute dont_touch of I26165: signal is true;
	signal I26166: std_logic; attribute dont_touch of I26166: signal is true;
	signal I26171: std_logic; attribute dont_touch of I26171: signal is true;
	signal I26172: std_logic; attribute dont_touch of I26172: signal is true;
	signal I26173: std_logic; attribute dont_touch of I26173: signal is true;
	signal I26174: std_logic; attribute dont_touch of I26174: signal is true;
	signal I26175: std_logic; attribute dont_touch of I26175: signal is true;
	signal I26180: std_logic; attribute dont_touch of I26180: signal is true;
	signal I26181: std_logic; attribute dont_touch of I26181: signal is true;
	signal I26182: std_logic; attribute dont_touch of I26182: signal is true;
	signal I26187: std_logic; attribute dont_touch of I26187: signal is true;
	signal I26188: std_logic; attribute dont_touch of I26188: signal is true;
	signal I26189: std_logic; attribute dont_touch of I26189: signal is true;
	signal I26190: std_logic; attribute dont_touch of I26190: signal is true;
	signal I26195: std_logic; attribute dont_touch of I26195: signal is true;
	signal I26196: std_logic; attribute dont_touch of I26196: signal is true;
	signal I26197: std_logic; attribute dont_touch of I26197: signal is true;
	signal I26202: std_logic; attribute dont_touch of I26202: signal is true;
	signal I26203: std_logic; attribute dont_touch of I26203: signal is true;
	signal I26204: std_logic; attribute dont_touch of I26204: signal is true;
	signal I26205: std_logic; attribute dont_touch of I26205: signal is true;
	signal I26206: std_logic; attribute dont_touch of I26206: signal is true;
	signal I26211: std_logic; attribute dont_touch of I26211: signal is true;
	signal I26212: std_logic; attribute dont_touch of I26212: signal is true;
	signal I26213: std_logic; attribute dont_touch of I26213: signal is true;
	signal I26218: std_logic; attribute dont_touch of I26218: signal is true;
	signal I26219: std_logic; attribute dont_touch of I26219: signal is true;
	signal I26220: std_logic; attribute dont_touch of I26220: signal is true;
	signal I26221: std_logic; attribute dont_touch of I26221: signal is true;
	signal I26226: std_logic; attribute dont_touch of I26226: signal is true;
	signal I26227: std_logic; attribute dont_touch of I26227: signal is true;
	signal I26228: std_logic; attribute dont_touch of I26228: signal is true;
	signal I26233: std_logic; attribute dont_touch of I26233: signal is true;
	signal I26234: std_logic; attribute dont_touch of I26234: signal is true;
	signal I26235: std_logic; attribute dont_touch of I26235: signal is true;
	signal I26236: std_logic; attribute dont_touch of I26236: signal is true;
	signal I26237: std_logic; attribute dont_touch of I26237: signal is true;
	signal I26242: std_logic; attribute dont_touch of I26242: signal is true;
	signal I26243: std_logic; attribute dont_touch of I26243: signal is true;
	signal I26244: std_logic; attribute dont_touch of I26244: signal is true;
	signal I26249: std_logic; attribute dont_touch of I26249: signal is true;
	signal I26250: std_logic; attribute dont_touch of I26250: signal is true;
	signal I26251: std_logic; attribute dont_touch of I26251: signal is true;
	signal I26252: std_logic; attribute dont_touch of I26252: signal is true;
	signal I26257: std_logic; attribute dont_touch of I26257: signal is true;
	signal I26258: std_logic; attribute dont_touch of I26258: signal is true;
	signal I26259: std_logic; attribute dont_touch of I26259: signal is true;
	signal I26264: std_logic; attribute dont_touch of I26264: signal is true;
	signal I26265: std_logic; attribute dont_touch of I26265: signal is true;
	signal I26266: std_logic; attribute dont_touch of I26266: signal is true;
	signal I26267: std_logic; attribute dont_touch of I26267: signal is true;
	signal I26268: std_logic; attribute dont_touch of I26268: signal is true;
	signal I26273: std_logic; attribute dont_touch of I26273: signal is true;
	signal I26274: std_logic; attribute dont_touch of I26274: signal is true;
	signal I26275: std_logic; attribute dont_touch of I26275: signal is true;
	signal I26280: std_logic; attribute dont_touch of I26280: signal is true;
	signal I26281: std_logic; attribute dont_touch of I26281: signal is true;
	signal I26282: std_logic; attribute dont_touch of I26282: signal is true;
	signal I26283: std_logic; attribute dont_touch of I26283: signal is true;
	signal I26288: std_logic; attribute dont_touch of I26288: signal is true;
	signal I26289: std_logic; attribute dont_touch of I26289: signal is true;
	signal I26290: std_logic; attribute dont_touch of I26290: signal is true;
	signal I26295: std_logic; attribute dont_touch of I26295: signal is true;
	signal I26296: std_logic; attribute dont_touch of I26296: signal is true;
	signal I26297: std_logic; attribute dont_touch of I26297: signal is true;
	signal I26298: std_logic; attribute dont_touch of I26298: signal is true;
	signal I26299: std_logic; attribute dont_touch of I26299: signal is true;
	signal I26304: std_logic; attribute dont_touch of I26304: signal is true;
	signal I26305: std_logic; attribute dont_touch of I26305: signal is true;
	signal I26306: std_logic; attribute dont_touch of I26306: signal is true;
	signal I26311: std_logic; attribute dont_touch of I26311: signal is true;
	signal I26312: std_logic; attribute dont_touch of I26312: signal is true;
	signal I26313: std_logic; attribute dont_touch of I26313: signal is true;
	signal I26314: std_logic; attribute dont_touch of I26314: signal is true;
	signal I26319: std_logic; attribute dont_touch of I26319: signal is true;
	signal I26320: std_logic; attribute dont_touch of I26320: signal is true;
	signal I26321: std_logic; attribute dont_touch of I26321: signal is true;
	signal I26326: std_logic; attribute dont_touch of I26326: signal is true;
	signal I26327: std_logic; attribute dont_touch of I26327: signal is true;
	signal I26328: std_logic; attribute dont_touch of I26328: signal is true;
	signal I26329: std_logic; attribute dont_touch of I26329: signal is true;
	signal I26330: std_logic; attribute dont_touch of I26330: signal is true;
	signal I26335: std_logic; attribute dont_touch of I26335: signal is true;
	signal I26336: std_logic; attribute dont_touch of I26336: signal is true;
	signal I26337: std_logic; attribute dont_touch of I26337: signal is true;
	signal I26342: std_logic; attribute dont_touch of I26342: signal is true;
	signal I26343: std_logic; attribute dont_touch of I26343: signal is true;
	signal I26344: std_logic; attribute dont_touch of I26344: signal is true;
	signal I26345: std_logic; attribute dont_touch of I26345: signal is true;
	signal I26350: std_logic; attribute dont_touch of I26350: signal is true;
	signal I26351: std_logic; attribute dont_touch of I26351: signal is true;
	signal I26352: std_logic; attribute dont_touch of I26352: signal is true;
	signal I26357: std_logic; attribute dont_touch of I26357: signal is true;
	signal I26358: std_logic; attribute dont_touch of I26358: signal is true;
	signal I26359: std_logic; attribute dont_touch of I26359: signal is true;
	signal I26360: std_logic; attribute dont_touch of I26360: signal is true;
	signal I26361: std_logic; attribute dont_touch of I26361: signal is true;
	signal I26366: std_logic; attribute dont_touch of I26366: signal is true;
	signal I26367: std_logic; attribute dont_touch of I26367: signal is true;
	signal I26368: std_logic; attribute dont_touch of I26368: signal is true;
	signal I26373: std_logic; attribute dont_touch of I26373: signal is true;
	signal I26374: std_logic; attribute dont_touch of I26374: signal is true;
	signal I26375: std_logic; attribute dont_touch of I26375: signal is true;
	signal I26376: std_logic; attribute dont_touch of I26376: signal is true;
	signal I26381: std_logic; attribute dont_touch of I26381: signal is true;
	signal I26382: std_logic; attribute dont_touch of I26382: signal is true;
	signal I26383: std_logic; attribute dont_touch of I26383: signal is true;
	signal I26388: std_logic; attribute dont_touch of I26388: signal is true;
	signal I26389: std_logic; attribute dont_touch of I26389: signal is true;
	signal I26390: std_logic; attribute dont_touch of I26390: signal is true;
	signal I26391: std_logic; attribute dont_touch of I26391: signal is true;
	signal I26392: std_logic; attribute dont_touch of I26392: signal is true;
	signal I26397: std_logic; attribute dont_touch of I26397: signal is true;
	signal I26398: std_logic; attribute dont_touch of I26398: signal is true;
	signal I26399: std_logic; attribute dont_touch of I26399: signal is true;
	signal I26404: std_logic; attribute dont_touch of I26404: signal is true;
	signal I26405: std_logic; attribute dont_touch of I26405: signal is true;
	signal I26406: std_logic; attribute dont_touch of I26406: signal is true;
	signal I26407: std_logic; attribute dont_touch of I26407: signal is true;
	signal I26412: std_logic; attribute dont_touch of I26412: signal is true;
	signal I26413: std_logic; attribute dont_touch of I26413: signal is true;
	signal I26414: std_logic; attribute dont_touch of I26414: signal is true;
	signal I26419: std_logic; attribute dont_touch of I26419: signal is true;
	signal I26420: std_logic; attribute dont_touch of I26420: signal is true;
	signal I26421: std_logic; attribute dont_touch of I26421: signal is true;
	signal I26422: std_logic; attribute dont_touch of I26422: signal is true;
	signal I26423: std_logic; attribute dont_touch of I26423: signal is true;
	signal I26428: std_logic; attribute dont_touch of I26428: signal is true;
	signal I26429: std_logic; attribute dont_touch of I26429: signal is true;
	signal I26430: std_logic; attribute dont_touch of I26430: signal is true;
	signal I26435: std_logic; attribute dont_touch of I26435: signal is true;
	signal I26436: std_logic; attribute dont_touch of I26436: signal is true;
	signal I26437: std_logic; attribute dont_touch of I26437: signal is true;
	signal I26438: std_logic; attribute dont_touch of I26438: signal is true;
	signal I26443: std_logic; attribute dont_touch of I26443: signal is true;
	signal I26444: std_logic; attribute dont_touch of I26444: signal is true;
	signal I26445: std_logic; attribute dont_touch of I26445: signal is true;
	signal I26450: std_logic; attribute dont_touch of I26450: signal is true;
	signal I26451: std_logic; attribute dont_touch of I26451: signal is true;
	signal I26452: std_logic; attribute dont_touch of I26452: signal is true;
	signal I26453: std_logic; attribute dont_touch of I26453: signal is true;
	signal I26454: std_logic; attribute dont_touch of I26454: signal is true;
	signal I26459: std_logic; attribute dont_touch of I26459: signal is true;
	signal I26460: std_logic; attribute dont_touch of I26460: signal is true;
	signal I26461: std_logic; attribute dont_touch of I26461: signal is true;
	signal I26466: std_logic; attribute dont_touch of I26466: signal is true;
	signal I26467: std_logic; attribute dont_touch of I26467: signal is true;
	signal I26468: std_logic; attribute dont_touch of I26468: signal is true;
	signal I26469: std_logic; attribute dont_touch of I26469: signal is true;
	signal I26474: std_logic; attribute dont_touch of I26474: signal is true;
	signal I26475: std_logic; attribute dont_touch of I26475: signal is true;
	signal I26476: std_logic; attribute dont_touch of I26476: signal is true;
	signal I26481: std_logic; attribute dont_touch of I26481: signal is true;
	signal I26482: std_logic; attribute dont_touch of I26482: signal is true;
	signal I26483: std_logic; attribute dont_touch of I26483: signal is true;
	signal I26484: std_logic; attribute dont_touch of I26484: signal is true;
	signal I26485: std_logic; attribute dont_touch of I26485: signal is true;
	signal I26490: std_logic; attribute dont_touch of I26490: signal is true;
	signal I26491: std_logic; attribute dont_touch of I26491: signal is true;
	signal I26492: std_logic; attribute dont_touch of I26492: signal is true;
	signal I26497: std_logic; attribute dont_touch of I26497: signal is true;
	signal I26498: std_logic; attribute dont_touch of I26498: signal is true;
	signal I26499: std_logic; attribute dont_touch of I26499: signal is true;
	signal I26500: std_logic; attribute dont_touch of I26500: signal is true;
	signal I26505: std_logic; attribute dont_touch of I26505: signal is true;
	signal I26506: std_logic; attribute dont_touch of I26506: signal is true;
	signal I26507: std_logic; attribute dont_touch of I26507: signal is true;
	signal I26512: std_logic; attribute dont_touch of I26512: signal is true;
	signal I26513: std_logic; attribute dont_touch of I26513: signal is true;
	signal I26514: std_logic; attribute dont_touch of I26514: signal is true;
	signal I26515: std_logic; attribute dont_touch of I26515: signal is true;
	signal I26516: std_logic; attribute dont_touch of I26516: signal is true;
	signal I26521: std_logic; attribute dont_touch of I26521: signal is true;
	signal I26522: std_logic; attribute dont_touch of I26522: signal is true;
	signal I26523: std_logic; attribute dont_touch of I26523: signal is true;
	signal I26528: std_logic; attribute dont_touch of I26528: signal is true;
	signal I26529: std_logic; attribute dont_touch of I26529: signal is true;
	signal I26530: std_logic; attribute dont_touch of I26530: signal is true;
	signal I26531: std_logic; attribute dont_touch of I26531: signal is true;
	signal I26536: std_logic; attribute dont_touch of I26536: signal is true;
	signal I26537: std_logic; attribute dont_touch of I26537: signal is true;
	signal I26538: std_logic; attribute dont_touch of I26538: signal is true;
	signal I26543: std_logic; attribute dont_touch of I26543: signal is true;
	signal I26544: std_logic; attribute dont_touch of I26544: signal is true;
	signal I26545: std_logic; attribute dont_touch of I26545: signal is true;
	signal I26546: std_logic; attribute dont_touch of I26546: signal is true;
	signal I26547: std_logic; attribute dont_touch of I26547: signal is true;
	signal I26552: std_logic; attribute dont_touch of I26552: signal is true;
	signal I26553: std_logic; attribute dont_touch of I26553: signal is true;
	signal I26554: std_logic; attribute dont_touch of I26554: signal is true;
	signal I26559: std_logic; attribute dont_touch of I26559: signal is true;
	signal I26560: std_logic; attribute dont_touch of I26560: signal is true;
	signal I26561: std_logic; attribute dont_touch of I26561: signal is true;
	signal I26562: std_logic; attribute dont_touch of I26562: signal is true;
	signal I26567: std_logic; attribute dont_touch of I26567: signal is true;
	signal I26568: std_logic; attribute dont_touch of I26568: signal is true;
	signal I26569: std_logic; attribute dont_touch of I26569: signal is true;
	signal I26574: std_logic; attribute dont_touch of I26574: signal is true;
	signal I26575: std_logic; attribute dont_touch of I26575: signal is true;
	signal I26576: std_logic; attribute dont_touch of I26576: signal is true;
	signal I26577: std_logic; attribute dont_touch of I26577: signal is true;
	signal I26578: std_logic; attribute dont_touch of I26578: signal is true;
	signal I26583: std_logic; attribute dont_touch of I26583: signal is true;
	signal I26584: std_logic; attribute dont_touch of I26584: signal is true;
	signal I26585: std_logic; attribute dont_touch of I26585: signal is true;
	signal I26590: std_logic; attribute dont_touch of I26590: signal is true;
	signal I26591: std_logic; attribute dont_touch of I26591: signal is true;
	signal I26592: std_logic; attribute dont_touch of I26592: signal is true;
	signal I26593: std_logic; attribute dont_touch of I26593: signal is true;
	signal I26598: std_logic; attribute dont_touch of I26598: signal is true;
	signal I26599: std_logic; attribute dont_touch of I26599: signal is true;
	signal I26600: std_logic; attribute dont_touch of I26600: signal is true;
	signal I26605: std_logic; attribute dont_touch of I26605: signal is true;
	signal I26606: std_logic; attribute dont_touch of I26606: signal is true;
	signal I26607: std_logic; attribute dont_touch of I26607: signal is true;
	signal I26608: std_logic; attribute dont_touch of I26608: signal is true;
	signal I26609: std_logic; attribute dont_touch of I26609: signal is true;
	signal I26614: std_logic; attribute dont_touch of I26614: signal is true;
	signal I26615: std_logic; attribute dont_touch of I26615: signal is true;
	signal I26616: std_logic; attribute dont_touch of I26616: signal is true;
	signal I26621: std_logic; attribute dont_touch of I26621: signal is true;
	signal I26622: std_logic; attribute dont_touch of I26622: signal is true;
	signal I26623: std_logic; attribute dont_touch of I26623: signal is true;
	signal I26624: std_logic; attribute dont_touch of I26624: signal is true;
	signal I26629: std_logic; attribute dont_touch of I26629: signal is true;
	signal I26630: std_logic; attribute dont_touch of I26630: signal is true;
	signal I26631: std_logic; attribute dont_touch of I26631: signal is true;
	signal I26636: std_logic; attribute dont_touch of I26636: signal is true;
	signal I26637: std_logic; attribute dont_touch of I26637: signal is true;
	signal I26638: std_logic; attribute dont_touch of I26638: signal is true;
	signal I26639: std_logic; attribute dont_touch of I26639: signal is true;
	signal I26640: std_logic; attribute dont_touch of I26640: signal is true;
	signal I26645: std_logic; attribute dont_touch of I26645: signal is true;
	signal I26646: std_logic; attribute dont_touch of I26646: signal is true;
	signal I26647: std_logic; attribute dont_touch of I26647: signal is true;
	signal I26652: std_logic; attribute dont_touch of I26652: signal is true;
	signal I26653: std_logic; attribute dont_touch of I26653: signal is true;
	signal I26654: std_logic; attribute dont_touch of I26654: signal is true;
	signal I26655: std_logic; attribute dont_touch of I26655: signal is true;
	signal I26660: std_logic; attribute dont_touch of I26660: signal is true;
	signal I26661: std_logic; attribute dont_touch of I26661: signal is true;
	signal I26662: std_logic; attribute dont_touch of I26662: signal is true;
	signal I26667: std_logic; attribute dont_touch of I26667: signal is true;
	signal I26668: std_logic; attribute dont_touch of I26668: signal is true;
	signal I26669: std_logic; attribute dont_touch of I26669: signal is true;
	signal I26670: std_logic; attribute dont_touch of I26670: signal is true;
	signal I26671: std_logic; attribute dont_touch of I26671: signal is true;
	signal I26676: std_logic; attribute dont_touch of I26676: signal is true;
	signal I26677: std_logic; attribute dont_touch of I26677: signal is true;
	signal I26678: std_logic; attribute dont_touch of I26678: signal is true;
	signal I26683: std_logic; attribute dont_touch of I26683: signal is true;
	signal I26684: std_logic; attribute dont_touch of I26684: signal is true;
	signal I26685: std_logic; attribute dont_touch of I26685: signal is true;
	signal I26686: std_logic; attribute dont_touch of I26686: signal is true;
	signal I26691: std_logic; attribute dont_touch of I26691: signal is true;
	signal I26692: std_logic; attribute dont_touch of I26692: signal is true;
	signal I26693: std_logic; attribute dont_touch of I26693: signal is true;
	signal I26698: std_logic; attribute dont_touch of I26698: signal is true;
	signal I26699: std_logic; attribute dont_touch of I26699: signal is true;
	signal I26700: std_logic; attribute dont_touch of I26700: signal is true;
	signal I26701: std_logic; attribute dont_touch of I26701: signal is true;
	signal I26702: std_logic; attribute dont_touch of I26702: signal is true;
	signal I26707: std_logic; attribute dont_touch of I26707: signal is true;
	signal I26708: std_logic; attribute dont_touch of I26708: signal is true;
	signal I26709: std_logic; attribute dont_touch of I26709: signal is true;
	signal I26714: std_logic; attribute dont_touch of I26714: signal is true;
	signal I26715: std_logic; attribute dont_touch of I26715: signal is true;
	signal I26716: std_logic; attribute dont_touch of I26716: signal is true;
	signal I26717: std_logic; attribute dont_touch of I26717: signal is true;
	signal I26722: std_logic; attribute dont_touch of I26722: signal is true;
	signal I26723: std_logic; attribute dont_touch of I26723: signal is true;
	signal I26724: std_logic; attribute dont_touch of I26724: signal is true;
	signal I26729: std_logic; attribute dont_touch of I26729: signal is true;
	signal I26730: std_logic; attribute dont_touch of I26730: signal is true;
	signal I26731: std_logic; attribute dont_touch of I26731: signal is true;
	signal I26732: std_logic; attribute dont_touch of I26732: signal is true;
	signal I26733: std_logic; attribute dont_touch of I26733: signal is true;
	signal I26738: std_logic; attribute dont_touch of I26738: signal is true;
	signal I26739: std_logic; attribute dont_touch of I26739: signal is true;
	signal I26740: std_logic; attribute dont_touch of I26740: signal is true;
	signal I26745: std_logic; attribute dont_touch of I26745: signal is true;
	signal I26746: std_logic; attribute dont_touch of I26746: signal is true;
	signal I26747: std_logic; attribute dont_touch of I26747: signal is true;
	signal I26748: std_logic; attribute dont_touch of I26748: signal is true;
	signal I26753: std_logic; attribute dont_touch of I26753: signal is true;
	signal I26754: std_logic; attribute dont_touch of I26754: signal is true;
	signal I26755: std_logic; attribute dont_touch of I26755: signal is true;
	signal I26760: std_logic; attribute dont_touch of I26760: signal is true;
	signal I26761: std_logic; attribute dont_touch of I26761: signal is true;
	signal I26762: std_logic; attribute dont_touch of I26762: signal is true;
	signal I26763: std_logic; attribute dont_touch of I26763: signal is true;
	signal I26764: std_logic; attribute dont_touch of I26764: signal is true;
	signal I26769: std_logic; attribute dont_touch of I26769: signal is true;
	signal I26770: std_logic; attribute dont_touch of I26770: signal is true;
	signal I26771: std_logic; attribute dont_touch of I26771: signal is true;
	signal I26776: std_logic; attribute dont_touch of I26776: signal is true;
	signal I26777: std_logic; attribute dont_touch of I26777: signal is true;
	signal I26778: std_logic; attribute dont_touch of I26778: signal is true;
	signal I26779: std_logic; attribute dont_touch of I26779: signal is true;
	signal I26784: std_logic; attribute dont_touch of I26784: signal is true;
	signal I26785: std_logic; attribute dont_touch of I26785: signal is true;
	signal I26786: std_logic; attribute dont_touch of I26786: signal is true;
	signal I26791: std_logic; attribute dont_touch of I26791: signal is true;
	signal I26792: std_logic; attribute dont_touch of I26792: signal is true;
	signal I26793: std_logic; attribute dont_touch of I26793: signal is true;
	signal I26794: std_logic; attribute dont_touch of I26794: signal is true;
	signal I26795: std_logic; attribute dont_touch of I26795: signal is true;
	signal I26800: std_logic; attribute dont_touch of I26800: signal is true;
	signal I26801: std_logic; attribute dont_touch of I26801: signal is true;
	signal I26802: std_logic; attribute dont_touch of I26802: signal is true;
	signal I26807: std_logic; attribute dont_touch of I26807: signal is true;
	signal I26808: std_logic; attribute dont_touch of I26808: signal is true;
	signal I26809: std_logic; attribute dont_touch of I26809: signal is true;
	signal I26810: std_logic; attribute dont_touch of I26810: signal is true;
	signal I26815: std_logic; attribute dont_touch of I26815: signal is true;
	signal I26816: std_logic; attribute dont_touch of I26816: signal is true;
	signal I26817: std_logic; attribute dont_touch of I26817: signal is true;
	signal I26822: std_logic; attribute dont_touch of I26822: signal is true;
	signal I26823: std_logic; attribute dont_touch of I26823: signal is true;
	signal I26824: std_logic; attribute dont_touch of I26824: signal is true;
	signal I26825: std_logic; attribute dont_touch of I26825: signal is true;
	signal I26826: std_logic; attribute dont_touch of I26826: signal is true;
	signal I26831: std_logic; attribute dont_touch of I26831: signal is true;
	signal I26832: std_logic; attribute dont_touch of I26832: signal is true;
	signal I26833: std_logic; attribute dont_touch of I26833: signal is true;
	signal I26838: std_logic; attribute dont_touch of I26838: signal is true;
	signal I26839: std_logic; attribute dont_touch of I26839: signal is true;
	signal I26840: std_logic; attribute dont_touch of I26840: signal is true;
	signal I26841: std_logic; attribute dont_touch of I26841: signal is true;
	signal I26846: std_logic; attribute dont_touch of I26846: signal is true;
	signal I26847: std_logic; attribute dont_touch of I26847: signal is true;
	signal I26848: std_logic; attribute dont_touch of I26848: signal is true;
	signal I26853: std_logic; attribute dont_touch of I26853: signal is true;
	signal I26854: std_logic; attribute dont_touch of I26854: signal is true;
	signal I26855: std_logic; attribute dont_touch of I26855: signal is true;
	signal I26856: std_logic; attribute dont_touch of I26856: signal is true;
	signal I26857: std_logic; attribute dont_touch of I26857: signal is true;
	signal I26862: std_logic; attribute dont_touch of I26862: signal is true;
	signal I26863: std_logic; attribute dont_touch of I26863: signal is true;
	signal I26864: std_logic; attribute dont_touch of I26864: signal is true;
	signal I26869: std_logic; attribute dont_touch of I26869: signal is true;
	signal I26870: std_logic; attribute dont_touch of I26870: signal is true;
	signal I26871: std_logic; attribute dont_touch of I26871: signal is true;
	signal I26872: std_logic; attribute dont_touch of I26872: signal is true;
	signal I26877: std_logic; attribute dont_touch of I26877: signal is true;
	signal I26878: std_logic; attribute dont_touch of I26878: signal is true;
	signal I26879: std_logic; attribute dont_touch of I26879: signal is true;
	signal I26884: std_logic; attribute dont_touch of I26884: signal is true;
	signal I26885: std_logic; attribute dont_touch of I26885: signal is true;
	signal I26886: std_logic; attribute dont_touch of I26886: signal is true;
	signal I26887: std_logic; attribute dont_touch of I26887: signal is true;
	signal I26888: std_logic; attribute dont_touch of I26888: signal is true;
	signal I26893: std_logic; attribute dont_touch of I26893: signal is true;
	signal I26894: std_logic; attribute dont_touch of I26894: signal is true;
	signal I26895: std_logic; attribute dont_touch of I26895: signal is true;
	signal I26900: std_logic; attribute dont_touch of I26900: signal is true;
	signal I26901: std_logic; attribute dont_touch of I26901: signal is true;
	signal I26902: std_logic; attribute dont_touch of I26902: signal is true;
	signal I26903: std_logic; attribute dont_touch of I26903: signal is true;
	signal I26908: std_logic; attribute dont_touch of I26908: signal is true;
	signal I26909: std_logic; attribute dont_touch of I26909: signal is true;
	signal I26910: std_logic; attribute dont_touch of I26910: signal is true;
	signal I26915: std_logic; attribute dont_touch of I26915: signal is true;
	signal I26916: std_logic; attribute dont_touch of I26916: signal is true;
	signal I26917: std_logic; attribute dont_touch of I26917: signal is true;
	signal I26918: std_logic; attribute dont_touch of I26918: signal is true;
	signal I26919: std_logic; attribute dont_touch of I26919: signal is true;
	signal I26924: std_logic; attribute dont_touch of I26924: signal is true;
	signal I26925: std_logic; attribute dont_touch of I26925: signal is true;
	signal I26926: std_logic; attribute dont_touch of I26926: signal is true;
	signal I26931: std_logic; attribute dont_touch of I26931: signal is true;
	signal I26932: std_logic; attribute dont_touch of I26932: signal is true;
	signal I26933: std_logic; attribute dont_touch of I26933: signal is true;
	signal I26934: std_logic; attribute dont_touch of I26934: signal is true;
	signal I26939: std_logic; attribute dont_touch of I26939: signal is true;
	signal I26940: std_logic; attribute dont_touch of I26940: signal is true;
	signal I26941: std_logic; attribute dont_touch of I26941: signal is true;
	signal I26946: std_logic; attribute dont_touch of I26946: signal is true;
	signal I26947: std_logic; attribute dont_touch of I26947: signal is true;
	signal I26948: std_logic; attribute dont_touch of I26948: signal is true;
	signal I26949: std_logic; attribute dont_touch of I26949: signal is true;
	signal I26950: std_logic; attribute dont_touch of I26950: signal is true;
	signal I26955: std_logic; attribute dont_touch of I26955: signal is true;
	signal I26956: std_logic; attribute dont_touch of I26956: signal is true;
	signal I26957: std_logic; attribute dont_touch of I26957: signal is true;
	signal I26962: std_logic; attribute dont_touch of I26962: signal is true;
	signal I26963: std_logic; attribute dont_touch of I26963: signal is true;
	signal I26964: std_logic; attribute dont_touch of I26964: signal is true;
	signal I26965: std_logic; attribute dont_touch of I26965: signal is true;
	signal I26970: std_logic; attribute dont_touch of I26970: signal is true;
	signal I26971: std_logic; attribute dont_touch of I26971: signal is true;
	signal I26972: std_logic; attribute dont_touch of I26972: signal is true;
	signal I26977: std_logic; attribute dont_touch of I26977: signal is true;
	signal I26978: std_logic; attribute dont_touch of I26978: signal is true;
	signal I26979: std_logic; attribute dont_touch of I26979: signal is true;
	signal I26980: std_logic; attribute dont_touch of I26980: signal is true;
	signal I26981: std_logic; attribute dont_touch of I26981: signal is true;
	signal I26986: std_logic; attribute dont_touch of I26986: signal is true;
	signal I26987: std_logic; attribute dont_touch of I26987: signal is true;
	signal I26988: std_logic; attribute dont_touch of I26988: signal is true;
	signal I26993: std_logic; attribute dont_touch of I26993: signal is true;
	signal I26994: std_logic; attribute dont_touch of I26994: signal is true;
	signal I26995: std_logic; attribute dont_touch of I26995: signal is true;
	signal I26996: std_logic; attribute dont_touch of I26996: signal is true;
	signal I27001: std_logic; attribute dont_touch of I27001: signal is true;
	signal I27002: std_logic; attribute dont_touch of I27002: signal is true;
	signal I27003: std_logic; attribute dont_touch of I27003: signal is true;
	signal I27082: std_logic; attribute dont_touch of I27082: signal is true;
	signal I27083: std_logic; attribute dont_touch of I27083: signal is true;
	signal I27084: std_logic; attribute dont_touch of I27084: signal is true;
	signal I27095: std_logic; attribute dont_touch of I27095: signal is true;
	signal I27096: std_logic; attribute dont_touch of I27096: signal is true;
	signal I27097: std_logic; attribute dont_touch of I27097: signal is true;
	signal I27108: std_logic; attribute dont_touch of I27108: signal is true;
	signal I27109: std_logic; attribute dont_touch of I27109: signal is true;
	signal I27110: std_logic; attribute dont_touch of I27110: signal is true;
	signal I27121: std_logic; attribute dont_touch of I27121: signal is true;
	signal I27122: std_logic; attribute dont_touch of I27122: signal is true;
	signal I27123: std_logic; attribute dont_touch of I27123: signal is true;
	signal I27134: std_logic; attribute dont_touch of I27134: signal is true;
	signal I27135: std_logic; attribute dont_touch of I27135: signal is true;
	signal I27136: std_logic; attribute dont_touch of I27136: signal is true;
	signal I27147: std_logic; attribute dont_touch of I27147: signal is true;
	signal I27148: std_logic; attribute dont_touch of I27148: signal is true;
	signal I27149: std_logic; attribute dont_touch of I27149: signal is true;
	signal I27160: std_logic; attribute dont_touch of I27160: signal is true;
	signal I27161: std_logic; attribute dont_touch of I27161: signal is true;
	signal I27162: std_logic; attribute dont_touch of I27162: signal is true;
	signal I27173: std_logic; attribute dont_touch of I27173: signal is true;
	signal I27174: std_logic; attribute dont_touch of I27174: signal is true;
	signal I27175: std_logic; attribute dont_touch of I27175: signal is true;
	signal I27186: std_logic; attribute dont_touch of I27186: signal is true;
	signal I27187: std_logic; attribute dont_touch of I27187: signal is true;
	signal I27188: std_logic; attribute dont_touch of I27188: signal is true;
	signal I27199: std_logic; attribute dont_touch of I27199: signal is true;
	signal I27200: std_logic; attribute dont_touch of I27200: signal is true;
	signal I27201: std_logic; attribute dont_touch of I27201: signal is true;
	signal I27212: std_logic; attribute dont_touch of I27212: signal is true;
	signal I27213: std_logic; attribute dont_touch of I27213: signal is true;
	signal I27214: std_logic; attribute dont_touch of I27214: signal is true;
	signal I27225: std_logic; attribute dont_touch of I27225: signal is true;
	signal I27226: std_logic; attribute dont_touch of I27226: signal is true;
	signal I27227: std_logic; attribute dont_touch of I27227: signal is true;
	signal I27238: std_logic; attribute dont_touch of I27238: signal is true;
	signal I27239: std_logic; attribute dont_touch of I27239: signal is true;
	signal I27240: std_logic; attribute dont_touch of I27240: signal is true;
	signal I27251: std_logic; attribute dont_touch of I27251: signal is true;
	signal I27252: std_logic; attribute dont_touch of I27252: signal is true;
	signal I27253: std_logic; attribute dont_touch of I27253: signal is true;
	signal I27264: std_logic; attribute dont_touch of I27264: signal is true;
	signal I27265: std_logic; attribute dont_touch of I27265: signal is true;
	signal I27266: std_logic; attribute dont_touch of I27266: signal is true;
	signal I27277: std_logic; attribute dont_touch of I27277: signal is true;
	signal I27278: std_logic; attribute dont_touch of I27278: signal is true;
	signal I27279: std_logic; attribute dont_touch of I27279: signal is true;
	signal I27290: std_logic; attribute dont_touch of I27290: signal is true;
	signal I27291: std_logic; attribute dont_touch of I27291: signal is true;
	signal I27292: std_logic; attribute dont_touch of I27292: signal is true;
	signal I27303: std_logic; attribute dont_touch of I27303: signal is true;
	signal I27304: std_logic; attribute dont_touch of I27304: signal is true;
	signal I27305: std_logic; attribute dont_touch of I27305: signal is true;
	signal I27316: std_logic; attribute dont_touch of I27316: signal is true;
	signal I27317: std_logic; attribute dont_touch of I27317: signal is true;
	signal I27318: std_logic; attribute dont_touch of I27318: signal is true;
	signal I27329: std_logic; attribute dont_touch of I27329: signal is true;
	signal I27330: std_logic; attribute dont_touch of I27330: signal is true;
	signal I27331: std_logic; attribute dont_touch of I27331: signal is true;
	signal I27342: std_logic; attribute dont_touch of I27342: signal is true;
	signal I27343: std_logic; attribute dont_touch of I27343: signal is true;
	signal I27344: std_logic; attribute dont_touch of I27344: signal is true;
	signal I27355: std_logic; attribute dont_touch of I27355: signal is true;
	signal I27356: std_logic; attribute dont_touch of I27356: signal is true;
	signal I27357: std_logic; attribute dont_touch of I27357: signal is true;
	signal I27368: std_logic; attribute dont_touch of I27368: signal is true;
	signal I27369: std_logic; attribute dont_touch of I27369: signal is true;
	signal I27370: std_logic; attribute dont_touch of I27370: signal is true;
	signal I27381: std_logic; attribute dont_touch of I27381: signal is true;
	signal I27382: std_logic; attribute dont_touch of I27382: signal is true;
	signal I27383: std_logic; attribute dont_touch of I27383: signal is true;
	signal I27394: std_logic; attribute dont_touch of I27394: signal is true;
	signal I27395: std_logic; attribute dont_touch of I27395: signal is true;
	signal I27396: std_logic; attribute dont_touch of I27396: signal is true;
	signal I27407: std_logic; attribute dont_touch of I27407: signal is true;
	signal I27408: std_logic; attribute dont_touch of I27408: signal is true;
	signal I27409: std_logic; attribute dont_touch of I27409: signal is true;
	signal I27420: std_logic; attribute dont_touch of I27420: signal is true;
	signal I27421: std_logic; attribute dont_touch of I27421: signal is true;
	signal I27422: std_logic; attribute dont_touch of I27422: signal is true;
	signal I27433: std_logic; attribute dont_touch of I27433: signal is true;
	signal I27434: std_logic; attribute dont_touch of I27434: signal is true;
	signal I27435: std_logic; attribute dont_touch of I27435: signal is true;
	signal I27446: std_logic; attribute dont_touch of I27446: signal is true;
	signal I27447: std_logic; attribute dont_touch of I27447: signal is true;
	signal I27448: std_logic; attribute dont_touch of I27448: signal is true;
	signal I27459: std_logic; attribute dont_touch of I27459: signal is true;
	signal I27460: std_logic; attribute dont_touch of I27460: signal is true;
	signal I27461: std_logic; attribute dont_touch of I27461: signal is true;
	signal I27472: std_logic; attribute dont_touch of I27472: signal is true;
	signal I27473: std_logic; attribute dont_touch of I27473: signal is true;
	signal I27474: std_logic; attribute dont_touch of I27474: signal is true;
	signal I27485: std_logic; attribute dont_touch of I27485: signal is true;
	signal I27486: std_logic; attribute dont_touch of I27486: signal is true;
	signal I27487: std_logic; attribute dont_touch of I27487: signal is true;
	signal I27499: std_logic; attribute dont_touch of I27499: signal is true;
	signal I27500: std_logic; attribute dont_touch of I27500: signal is true;
	signal I27501: std_logic; attribute dont_touch of I27501: signal is true;
	signal I27502: std_logic; attribute dont_touch of I27502: signal is true;
	signal I27507: std_logic; attribute dont_touch of I27507: signal is true;
	signal I27508: std_logic; attribute dont_touch of I27508: signal is true;
	signal I27509: std_logic; attribute dont_touch of I27509: signal is true;
	signal I27514: std_logic; attribute dont_touch of I27514: signal is true;
	signal I27515: std_logic; attribute dont_touch of I27515: signal is true;
	signal I27516: std_logic; attribute dont_touch of I27516: signal is true;
	signal I27517: std_logic; attribute dont_touch of I27517: signal is true;
	signal I27522: std_logic; attribute dont_touch of I27522: signal is true;
	signal I27523: std_logic; attribute dont_touch of I27523: signal is true;
	signal I27524: std_logic; attribute dont_touch of I27524: signal is true;
	signal I27529: std_logic; attribute dont_touch of I27529: signal is true;
	signal I27530: std_logic; attribute dont_touch of I27530: signal is true;
	signal I27531: std_logic; attribute dont_touch of I27531: signal is true;
	signal I27532: std_logic; attribute dont_touch of I27532: signal is true;
	signal I27537: std_logic; attribute dont_touch of I27537: signal is true;
	signal I27538: std_logic; attribute dont_touch of I27538: signal is true;
	signal I27539: std_logic; attribute dont_touch of I27539: signal is true;
	signal I27544: std_logic; attribute dont_touch of I27544: signal is true;
	signal I27545: std_logic; attribute dont_touch of I27545: signal is true;
	signal I27546: std_logic; attribute dont_touch of I27546: signal is true;
	signal I27551: std_logic; attribute dont_touch of I27551: signal is true;
	signal I27552: std_logic; attribute dont_touch of I27552: signal is true;
	signal I27553: std_logic; attribute dont_touch of I27553: signal is true;
	signal I27558: std_logic; attribute dont_touch of I27558: signal is true;
	signal I27559: std_logic; attribute dont_touch of I27559: signal is true;
	signal I27560: std_logic; attribute dont_touch of I27560: signal is true;
	signal I27565: std_logic; attribute dont_touch of I27565: signal is true;
	signal I27566: std_logic; attribute dont_touch of I27566: signal is true;
	signal I27567: std_logic; attribute dont_touch of I27567: signal is true;
	signal I27572: std_logic; attribute dont_touch of I27572: signal is true;
	signal I27573: std_logic; attribute dont_touch of I27573: signal is true;
	signal I27574: std_logic; attribute dont_touch of I27574: signal is true;
	signal I27579: std_logic; attribute dont_touch of I27579: signal is true;
	signal I27580: std_logic; attribute dont_touch of I27580: signal is true;
	signal I27581: std_logic; attribute dont_touch of I27581: signal is true;
	signal I27586: std_logic; attribute dont_touch of I27586: signal is true;
	signal I27587: std_logic; attribute dont_touch of I27587: signal is true;
	signal I27588: std_logic; attribute dont_touch of I27588: signal is true;
	signal I27593: std_logic; attribute dont_touch of I27593: signal is true;
	signal I27594: std_logic; attribute dont_touch of I27594: signal is true;
	signal I27595: std_logic; attribute dont_touch of I27595: signal is true;
	signal I27600: std_logic; attribute dont_touch of I27600: signal is true;
	signal I27601: std_logic; attribute dont_touch of I27601: signal is true;
	signal I27602: std_logic; attribute dont_touch of I27602: signal is true;
	signal I27607: std_logic; attribute dont_touch of I27607: signal is true;
	signal I27608: std_logic; attribute dont_touch of I27608: signal is true;
	signal I27609: std_logic; attribute dont_touch of I27609: signal is true;
	signal I27614: std_logic; attribute dont_touch of I27614: signal is true;
	signal I27615: std_logic; attribute dont_touch of I27615: signal is true;
	signal I27616: std_logic; attribute dont_touch of I27616: signal is true;
	signal I27621: std_logic; attribute dont_touch of I27621: signal is true;
	signal I27622: std_logic; attribute dont_touch of I27622: signal is true;
	signal I27623: std_logic; attribute dont_touch of I27623: signal is true;
	signal I27628: std_logic; attribute dont_touch of I27628: signal is true;
	signal I27629: std_logic; attribute dont_touch of I27629: signal is true;
	signal I27630: std_logic; attribute dont_touch of I27630: signal is true;
	signal I27635: std_logic; attribute dont_touch of I27635: signal is true;
	signal I27636: std_logic; attribute dont_touch of I27636: signal is true;
	signal I27637: std_logic; attribute dont_touch of I27637: signal is true;
	signal I27642: std_logic; attribute dont_touch of I27642: signal is true;
	signal I27643: std_logic; attribute dont_touch of I27643: signal is true;
	signal I27644: std_logic; attribute dont_touch of I27644: signal is true;
	signal I27649: std_logic; attribute dont_touch of I27649: signal is true;
	signal I27650: std_logic; attribute dont_touch of I27650: signal is true;
	signal I27651: std_logic; attribute dont_touch of I27651: signal is true;
	signal I27656: std_logic; attribute dont_touch of I27656: signal is true;
	signal I27657: std_logic; attribute dont_touch of I27657: signal is true;
	signal I27658: std_logic; attribute dont_touch of I27658: signal is true;
	signal I27663: std_logic; attribute dont_touch of I27663: signal is true;
	signal I27664: std_logic; attribute dont_touch of I27664: signal is true;
	signal I27665: std_logic; attribute dont_touch of I27665: signal is true;
	signal I27670: std_logic; attribute dont_touch of I27670: signal is true;
	signal I27671: std_logic; attribute dont_touch of I27671: signal is true;
	signal I27672: std_logic; attribute dont_touch of I27672: signal is true;
	signal I27677: std_logic; attribute dont_touch of I27677: signal is true;
	signal I27678: std_logic; attribute dont_touch of I27678: signal is true;
	signal I27679: std_logic; attribute dont_touch of I27679: signal is true;
	signal I27684: std_logic; attribute dont_touch of I27684: signal is true;
	signal I27685: std_logic; attribute dont_touch of I27685: signal is true;
	signal I27686: std_logic; attribute dont_touch of I27686: signal is true;
	signal I27691: std_logic; attribute dont_touch of I27691: signal is true;
	signal I27692: std_logic; attribute dont_touch of I27692: signal is true;
	signal I27693: std_logic; attribute dont_touch of I27693: signal is true;
	signal I27698: std_logic; attribute dont_touch of I27698: signal is true;
	signal I27699: std_logic; attribute dont_touch of I27699: signal is true;
	signal I27700: std_logic; attribute dont_touch of I27700: signal is true;
	signal I27705: std_logic; attribute dont_touch of I27705: signal is true;
	signal I27706: std_logic; attribute dont_touch of I27706: signal is true;
	signal I27707: std_logic; attribute dont_touch of I27707: signal is true;
	signal I27712: std_logic; attribute dont_touch of I27712: signal is true;
	signal I27713: std_logic; attribute dont_touch of I27713: signal is true;
	signal I27714: std_logic; attribute dont_touch of I27714: signal is true;
	signal I27719: std_logic; attribute dont_touch of I27719: signal is true;
	signal I27720: std_logic; attribute dont_touch of I27720: signal is true;
	signal I27721: std_logic; attribute dont_touch of I27721: signal is true;
	signal I27726: std_logic; attribute dont_touch of I27726: signal is true;
	signal I27727: std_logic; attribute dont_touch of I27727: signal is true;
	signal I27728: std_logic; attribute dont_touch of I27728: signal is true;
	signal I27733: std_logic; attribute dont_touch of I27733: signal is true;
	signal I27734: std_logic; attribute dont_touch of I27734: signal is true;
	signal I27735: std_logic; attribute dont_touch of I27735: signal is true;
	signal I27740: std_logic; attribute dont_touch of I27740: signal is true;
	signal I27741: std_logic; attribute dont_touch of I27741: signal is true;
	signal I27742: std_logic; attribute dont_touch of I27742: signal is true;
	signal I30021: std_logic; attribute dont_touch of I30021: signal is true;
	signal I30022: std_logic; attribute dont_touch of I30022: signal is true;
	signal I30023: std_logic; attribute dont_touch of I30023: signal is true;
	signal I30024: std_logic; attribute dont_touch of I30024: signal is true;
	signal I30025: std_logic; attribute dont_touch of I30025: signal is true;
	signal I30030: std_logic; attribute dont_touch of I30030: signal is true;
	signal I30031: std_logic; attribute dont_touch of I30031: signal is true;
	signal I30032: std_logic; attribute dont_touch of I30032: signal is true;
	signal I30037: std_logic; attribute dont_touch of I30037: signal is true;
	signal I30038: std_logic; attribute dont_touch of I30038: signal is true;
	signal I30039: std_logic; attribute dont_touch of I30039: signal is true;
	signal I30040: std_logic; attribute dont_touch of I30040: signal is true;
	signal I30045: std_logic; attribute dont_touch of I30045: signal is true;
	signal I30046: std_logic; attribute dont_touch of I30046: signal is true;
	signal I30047: std_logic; attribute dont_touch of I30047: signal is true;
	signal I30052: std_logic; attribute dont_touch of I30052: signal is true;
	signal I30053: std_logic; attribute dont_touch of I30053: signal is true;
	signal I30054: std_logic; attribute dont_touch of I30054: signal is true;
	signal I30055: std_logic; attribute dont_touch of I30055: signal is true;
	signal I30056: std_logic; attribute dont_touch of I30056: signal is true;
	signal I30061: std_logic; attribute dont_touch of I30061: signal is true;
	signal I30062: std_logic; attribute dont_touch of I30062: signal is true;
	signal I30063: std_logic; attribute dont_touch of I30063: signal is true;
	signal I30068: std_logic; attribute dont_touch of I30068: signal is true;
	signal I30069: std_logic; attribute dont_touch of I30069: signal is true;
	signal I30070: std_logic; attribute dont_touch of I30070: signal is true;
	signal I30071: std_logic; attribute dont_touch of I30071: signal is true;
	signal I30076: std_logic; attribute dont_touch of I30076: signal is true;
	signal I30077: std_logic; attribute dont_touch of I30077: signal is true;
	signal I30078: std_logic; attribute dont_touch of I30078: signal is true;
	signal I30083: std_logic; attribute dont_touch of I30083: signal is true;
	signal I30084: std_logic; attribute dont_touch of I30084: signal is true;
	signal I30085: std_logic; attribute dont_touch of I30085: signal is true;
	signal I30086: std_logic; attribute dont_touch of I30086: signal is true;
	signal I30087: std_logic; attribute dont_touch of I30087: signal is true;
	signal I30092: std_logic; attribute dont_touch of I30092: signal is true;
	signal I30093: std_logic; attribute dont_touch of I30093: signal is true;
	signal I30094: std_logic; attribute dont_touch of I30094: signal is true;
	signal I30099: std_logic; attribute dont_touch of I30099: signal is true;
	signal I30100: std_logic; attribute dont_touch of I30100: signal is true;
	signal I30101: std_logic; attribute dont_touch of I30101: signal is true;
	signal I30102: std_logic; attribute dont_touch of I30102: signal is true;
	signal I30107: std_logic; attribute dont_touch of I30107: signal is true;
	signal I30108: std_logic; attribute dont_touch of I30108: signal is true;
	signal I30109: std_logic; attribute dont_touch of I30109: signal is true;
	signal I30114: std_logic; attribute dont_touch of I30114: signal is true;
	signal I30115: std_logic; attribute dont_touch of I30115: signal is true;
	signal I30116: std_logic; attribute dont_touch of I30116: signal is true;
	signal I30117: std_logic; attribute dont_touch of I30117: signal is true;
	signal I30118: std_logic; attribute dont_touch of I30118: signal is true;
	signal I30123: std_logic; attribute dont_touch of I30123: signal is true;
	signal I30124: std_logic; attribute dont_touch of I30124: signal is true;
	signal I30125: std_logic; attribute dont_touch of I30125: signal is true;
	signal I30130: std_logic; attribute dont_touch of I30130: signal is true;
	signal I30131: std_logic; attribute dont_touch of I30131: signal is true;
	signal I30132: std_logic; attribute dont_touch of I30132: signal is true;
	signal I30133: std_logic; attribute dont_touch of I30133: signal is true;
	signal I30138: std_logic; attribute dont_touch of I30138: signal is true;
	signal I30139: std_logic; attribute dont_touch of I30139: signal is true;
	signal I30140: std_logic; attribute dont_touch of I30140: signal is true;
	signal I30145: std_logic; attribute dont_touch of I30145: signal is true;
	signal I30146: std_logic; attribute dont_touch of I30146: signal is true;
	signal I30147: std_logic; attribute dont_touch of I30147: signal is true;
	signal I30148: std_logic; attribute dont_touch of I30148: signal is true;
	signal I30149: std_logic; attribute dont_touch of I30149: signal is true;
	signal I30154: std_logic; attribute dont_touch of I30154: signal is true;
	signal I30155: std_logic; attribute dont_touch of I30155: signal is true;
	signal I30156: std_logic; attribute dont_touch of I30156: signal is true;
	signal I30161: std_logic; attribute dont_touch of I30161: signal is true;
	signal I30162: std_logic; attribute dont_touch of I30162: signal is true;
	signal I30163: std_logic; attribute dont_touch of I30163: signal is true;
	signal I30164: std_logic; attribute dont_touch of I30164: signal is true;
	signal I30169: std_logic; attribute dont_touch of I30169: signal is true;
	signal I30170: std_logic; attribute dont_touch of I30170: signal is true;
	signal I30171: std_logic; attribute dont_touch of I30171: signal is true;
	signal I30176: std_logic; attribute dont_touch of I30176: signal is true;
	signal I30177: std_logic; attribute dont_touch of I30177: signal is true;
	signal I30178: std_logic; attribute dont_touch of I30178: signal is true;
	signal I30179: std_logic; attribute dont_touch of I30179: signal is true;
	signal I30180: std_logic; attribute dont_touch of I30180: signal is true;
	signal I30185: std_logic; attribute dont_touch of I30185: signal is true;
	signal I30186: std_logic; attribute dont_touch of I30186: signal is true;
	signal I30187: std_logic; attribute dont_touch of I30187: signal is true;
	signal I30192: std_logic; attribute dont_touch of I30192: signal is true;
	signal I30193: std_logic; attribute dont_touch of I30193: signal is true;
	signal I30194: std_logic; attribute dont_touch of I30194: signal is true;
	signal I30195: std_logic; attribute dont_touch of I30195: signal is true;
	signal I30200: std_logic; attribute dont_touch of I30200: signal is true;
	signal I30201: std_logic; attribute dont_touch of I30201: signal is true;
	signal I30202: std_logic; attribute dont_touch of I30202: signal is true;
	signal I30207: std_logic; attribute dont_touch of I30207: signal is true;
	signal I30208: std_logic; attribute dont_touch of I30208: signal is true;
	signal I30209: std_logic; attribute dont_touch of I30209: signal is true;
	signal I30210: std_logic; attribute dont_touch of I30210: signal is true;
	signal I30211: std_logic; attribute dont_touch of I30211: signal is true;
	signal I30216: std_logic; attribute dont_touch of I30216: signal is true;
	signal I30217: std_logic; attribute dont_touch of I30217: signal is true;
	signal I30218: std_logic; attribute dont_touch of I30218: signal is true;
	signal I30223: std_logic; attribute dont_touch of I30223: signal is true;
	signal I30224: std_logic; attribute dont_touch of I30224: signal is true;
	signal I30225: std_logic; attribute dont_touch of I30225: signal is true;
	signal I30226: std_logic; attribute dont_touch of I30226: signal is true;
	signal I30231: std_logic; attribute dont_touch of I30231: signal is true;
	signal I30232: std_logic; attribute dont_touch of I30232: signal is true;
	signal I30233: std_logic; attribute dont_touch of I30233: signal is true;
	signal I30238: std_logic; attribute dont_touch of I30238: signal is true;
	signal I30239: std_logic; attribute dont_touch of I30239: signal is true;
	signal I30240: std_logic; attribute dont_touch of I30240: signal is true;
	signal I30241: std_logic; attribute dont_touch of I30241: signal is true;
	signal I30242: std_logic; attribute dont_touch of I30242: signal is true;
	signal I30247: std_logic; attribute dont_touch of I30247: signal is true;
	signal I30248: std_logic; attribute dont_touch of I30248: signal is true;
	signal I30249: std_logic; attribute dont_touch of I30249: signal is true;
	signal I30254: std_logic; attribute dont_touch of I30254: signal is true;
	signal I30255: std_logic; attribute dont_touch of I30255: signal is true;
	signal I30256: std_logic; attribute dont_touch of I30256: signal is true;
	signal I30257: std_logic; attribute dont_touch of I30257: signal is true;
	signal I30262: std_logic; attribute dont_touch of I30262: signal is true;
	signal I30263: std_logic; attribute dont_touch of I30263: signal is true;
	signal I30264: std_logic; attribute dont_touch of I30264: signal is true;
	signal I30269: std_logic; attribute dont_touch of I30269: signal is true;
	signal I30270: std_logic; attribute dont_touch of I30270: signal is true;
	signal I30271: std_logic; attribute dont_touch of I30271: signal is true;
	signal I30272: std_logic; attribute dont_touch of I30272: signal is true;
	signal I30273: std_logic; attribute dont_touch of I30273: signal is true;
	signal I30278: std_logic; attribute dont_touch of I30278: signal is true;
	signal I30279: std_logic; attribute dont_touch of I30279: signal is true;
	signal I30280: std_logic; attribute dont_touch of I30280: signal is true;
	signal I30285: std_logic; attribute dont_touch of I30285: signal is true;
	signal I30286: std_logic; attribute dont_touch of I30286: signal is true;
	signal I30287: std_logic; attribute dont_touch of I30287: signal is true;
	signal I30288: std_logic; attribute dont_touch of I30288: signal is true;
	signal I30293: std_logic; attribute dont_touch of I30293: signal is true;
	signal I30294: std_logic; attribute dont_touch of I30294: signal is true;
	signal I30295: std_logic; attribute dont_touch of I30295: signal is true;
	signal I30300: std_logic; attribute dont_touch of I30300: signal is true;
	signal I30301: std_logic; attribute dont_touch of I30301: signal is true;
	signal I30302: std_logic; attribute dont_touch of I30302: signal is true;
	signal I30303: std_logic; attribute dont_touch of I30303: signal is true;
	signal I30304: std_logic; attribute dont_touch of I30304: signal is true;
	signal I30309: std_logic; attribute dont_touch of I30309: signal is true;
	signal I30310: std_logic; attribute dont_touch of I30310: signal is true;
	signal I30311: std_logic; attribute dont_touch of I30311: signal is true;
	signal I30316: std_logic; attribute dont_touch of I30316: signal is true;
	signal I30317: std_logic; attribute dont_touch of I30317: signal is true;
	signal I30318: std_logic; attribute dont_touch of I30318: signal is true;
	signal I30319: std_logic; attribute dont_touch of I30319: signal is true;
	signal I30324: std_logic; attribute dont_touch of I30324: signal is true;
	signal I30325: std_logic; attribute dont_touch of I30325: signal is true;
	signal I30326: std_logic; attribute dont_touch of I30326: signal is true;
	signal I30331: std_logic; attribute dont_touch of I30331: signal is true;
	signal I30332: std_logic; attribute dont_touch of I30332: signal is true;
	signal I30333: std_logic; attribute dont_touch of I30333: signal is true;
	signal I30334: std_logic; attribute dont_touch of I30334: signal is true;
	signal I30335: std_logic; attribute dont_touch of I30335: signal is true;
	signal I30340: std_logic; attribute dont_touch of I30340: signal is true;
	signal I30341: std_logic; attribute dont_touch of I30341: signal is true;
	signal I30342: std_logic; attribute dont_touch of I30342: signal is true;
	signal I30347: std_logic; attribute dont_touch of I30347: signal is true;
	signal I30348: std_logic; attribute dont_touch of I30348: signal is true;
	signal I30349: std_logic; attribute dont_touch of I30349: signal is true;
	signal I30350: std_logic; attribute dont_touch of I30350: signal is true;
	signal I30355: std_logic; attribute dont_touch of I30355: signal is true;
	signal I30356: std_logic; attribute dont_touch of I30356: signal is true;
	signal I30357: std_logic; attribute dont_touch of I30357: signal is true;
	signal I30362: std_logic; attribute dont_touch of I30362: signal is true;
	signal I30363: std_logic; attribute dont_touch of I30363: signal is true;
	signal I30364: std_logic; attribute dont_touch of I30364: signal is true;
	signal I30365: std_logic; attribute dont_touch of I30365: signal is true;
	signal I30366: std_logic; attribute dont_touch of I30366: signal is true;
	signal I30371: std_logic; attribute dont_touch of I30371: signal is true;
	signal I30372: std_logic; attribute dont_touch of I30372: signal is true;
	signal I30373: std_logic; attribute dont_touch of I30373: signal is true;
	signal I30378: std_logic; attribute dont_touch of I30378: signal is true;
	signal I30379: std_logic; attribute dont_touch of I30379: signal is true;
	signal I30380: std_logic; attribute dont_touch of I30380: signal is true;
	signal I30381: std_logic; attribute dont_touch of I30381: signal is true;
	signal I30386: std_logic; attribute dont_touch of I30386: signal is true;
	signal I30387: std_logic; attribute dont_touch of I30387: signal is true;
	signal I30388: std_logic; attribute dont_touch of I30388: signal is true;
	signal I30393: std_logic; attribute dont_touch of I30393: signal is true;
	signal I30394: std_logic; attribute dont_touch of I30394: signal is true;
	signal I30395: std_logic; attribute dont_touch of I30395: signal is true;
	signal I30396: std_logic; attribute dont_touch of I30396: signal is true;
	signal I30397: std_logic; attribute dont_touch of I30397: signal is true;
	signal I30402: std_logic; attribute dont_touch of I30402: signal is true;
	signal I30403: std_logic; attribute dont_touch of I30403: signal is true;
	signal I30404: std_logic; attribute dont_touch of I30404: signal is true;
	signal I30409: std_logic; attribute dont_touch of I30409: signal is true;
	signal I30410: std_logic; attribute dont_touch of I30410: signal is true;
	signal I30411: std_logic; attribute dont_touch of I30411: signal is true;
	signal I30412: std_logic; attribute dont_touch of I30412: signal is true;
	signal I30417: std_logic; attribute dont_touch of I30417: signal is true;
	signal I30418: std_logic; attribute dont_touch of I30418: signal is true;
	signal I30419: std_logic; attribute dont_touch of I30419: signal is true;
	signal I30424: std_logic; attribute dont_touch of I30424: signal is true;
	signal I30425: std_logic; attribute dont_touch of I30425: signal is true;
	signal I30426: std_logic; attribute dont_touch of I30426: signal is true;
	signal I30427: std_logic; attribute dont_touch of I30427: signal is true;
	signal I30428: std_logic; attribute dont_touch of I30428: signal is true;
	signal I30433: std_logic; attribute dont_touch of I30433: signal is true;
	signal I30434: std_logic; attribute dont_touch of I30434: signal is true;
	signal I30435: std_logic; attribute dont_touch of I30435: signal is true;
	signal I30440: std_logic; attribute dont_touch of I30440: signal is true;
	signal I30441: std_logic; attribute dont_touch of I30441: signal is true;
	signal I30442: std_logic; attribute dont_touch of I30442: signal is true;
	signal I30443: std_logic; attribute dont_touch of I30443: signal is true;
	signal I30448: std_logic; attribute dont_touch of I30448: signal is true;
	signal I30449: std_logic; attribute dont_touch of I30449: signal is true;
	signal I30450: std_logic; attribute dont_touch of I30450: signal is true;
	signal I30455: std_logic; attribute dont_touch of I30455: signal is true;
	signal I30456: std_logic; attribute dont_touch of I30456: signal is true;
	signal I30457: std_logic; attribute dont_touch of I30457: signal is true;
	signal I30458: std_logic; attribute dont_touch of I30458: signal is true;
	signal I30459: std_logic; attribute dont_touch of I30459: signal is true;
	signal I30464: std_logic; attribute dont_touch of I30464: signal is true;
	signal I30465: std_logic; attribute dont_touch of I30465: signal is true;
	signal I30466: std_logic; attribute dont_touch of I30466: signal is true;
	signal I30471: std_logic; attribute dont_touch of I30471: signal is true;
	signal I30472: std_logic; attribute dont_touch of I30472: signal is true;
	signal I30473: std_logic; attribute dont_touch of I30473: signal is true;
	signal I30474: std_logic; attribute dont_touch of I30474: signal is true;
	signal I30479: std_logic; attribute dont_touch of I30479: signal is true;
	signal I30480: std_logic; attribute dont_touch of I30480: signal is true;
	signal I30481: std_logic; attribute dont_touch of I30481: signal is true;
	signal I30486: std_logic; attribute dont_touch of I30486: signal is true;
	signal I30487: std_logic; attribute dont_touch of I30487: signal is true;
	signal I30488: std_logic; attribute dont_touch of I30488: signal is true;
	signal I30489: std_logic; attribute dont_touch of I30489: signal is true;
	signal I30490: std_logic; attribute dont_touch of I30490: signal is true;
	signal I30495: std_logic; attribute dont_touch of I30495: signal is true;
	signal I30496: std_logic; attribute dont_touch of I30496: signal is true;
	signal I30497: std_logic; attribute dont_touch of I30497: signal is true;
	signal I30502: std_logic; attribute dont_touch of I30502: signal is true;
	signal I30503: std_logic; attribute dont_touch of I30503: signal is true;
	signal I30504: std_logic; attribute dont_touch of I30504: signal is true;
	signal I30505: std_logic; attribute dont_touch of I30505: signal is true;
	signal I30510: std_logic; attribute dont_touch of I30510: signal is true;
	signal I30511: std_logic; attribute dont_touch of I30511: signal is true;
	signal I30512: std_logic; attribute dont_touch of I30512: signal is true;
	signal I30517: std_logic; attribute dont_touch of I30517: signal is true;
	signal I30518: std_logic; attribute dont_touch of I30518: signal is true;
	signal I30519: std_logic; attribute dont_touch of I30519: signal is true;
	signal I30520: std_logic; attribute dont_touch of I30520: signal is true;
	signal I30521: std_logic; attribute dont_touch of I30521: signal is true;
	signal I30526: std_logic; attribute dont_touch of I30526: signal is true;
	signal I30527: std_logic; attribute dont_touch of I30527: signal is true;
	signal I30528: std_logic; attribute dont_touch of I30528: signal is true;
	signal I30533: std_logic; attribute dont_touch of I30533: signal is true;
	signal I30534: std_logic; attribute dont_touch of I30534: signal is true;
	signal I30535: std_logic; attribute dont_touch of I30535: signal is true;
	signal I30536: std_logic; attribute dont_touch of I30536: signal is true;
	signal I30541: std_logic; attribute dont_touch of I30541: signal is true;
	signal I30542: std_logic; attribute dont_touch of I30542: signal is true;
	signal I30543: std_logic; attribute dont_touch of I30543: signal is true;
	signal I30548: std_logic; attribute dont_touch of I30548: signal is true;
	signal I30549: std_logic; attribute dont_touch of I30549: signal is true;
	signal I30550: std_logic; attribute dont_touch of I30550: signal is true;
	signal I30551: std_logic; attribute dont_touch of I30551: signal is true;
	signal I30552: std_logic; attribute dont_touch of I30552: signal is true;
	signal I30557: std_logic; attribute dont_touch of I30557: signal is true;
	signal I30558: std_logic; attribute dont_touch of I30558: signal is true;
	signal I30559: std_logic; attribute dont_touch of I30559: signal is true;
	signal I30564: std_logic; attribute dont_touch of I30564: signal is true;
	signal I30565: std_logic; attribute dont_touch of I30565: signal is true;
	signal I30566: std_logic; attribute dont_touch of I30566: signal is true;
	signal I30567: std_logic; attribute dont_touch of I30567: signal is true;
	signal I30572: std_logic; attribute dont_touch of I30572: signal is true;
	signal I30573: std_logic; attribute dont_touch of I30573: signal is true;
	signal I30574: std_logic; attribute dont_touch of I30574: signal is true;
	signal I30579: std_logic; attribute dont_touch of I30579: signal is true;
	signal I30580: std_logic; attribute dont_touch of I30580: signal is true;
	signal I30581: std_logic; attribute dont_touch of I30581: signal is true;
	signal I30582: std_logic; attribute dont_touch of I30582: signal is true;
	signal I30583: std_logic; attribute dont_touch of I30583: signal is true;
	signal I30588: std_logic; attribute dont_touch of I30588: signal is true;
	signal I30589: std_logic; attribute dont_touch of I30589: signal is true;
	signal I30590: std_logic; attribute dont_touch of I30590: signal is true;
	signal I30595: std_logic; attribute dont_touch of I30595: signal is true;
	signal I30596: std_logic; attribute dont_touch of I30596: signal is true;
	signal I30597: std_logic; attribute dont_touch of I30597: signal is true;
	signal I30598: std_logic; attribute dont_touch of I30598: signal is true;
	signal I30603: std_logic; attribute dont_touch of I30603: signal is true;
	signal I30604: std_logic; attribute dont_touch of I30604: signal is true;
	signal I30605: std_logic; attribute dont_touch of I30605: signal is true;
	signal I30610: std_logic; attribute dont_touch of I30610: signal is true;
	signal I30611: std_logic; attribute dont_touch of I30611: signal is true;
	signal I30612: std_logic; attribute dont_touch of I30612: signal is true;
	signal I30613: std_logic; attribute dont_touch of I30613: signal is true;
	signal I30614: std_logic; attribute dont_touch of I30614: signal is true;
	signal I30619: std_logic; attribute dont_touch of I30619: signal is true;
	signal I30620: std_logic; attribute dont_touch of I30620: signal is true;
	signal I30621: std_logic; attribute dont_touch of I30621: signal is true;
	signal I30626: std_logic; attribute dont_touch of I30626: signal is true;
	signal I30627: std_logic; attribute dont_touch of I30627: signal is true;
	signal I30628: std_logic; attribute dont_touch of I30628: signal is true;
	signal I30629: std_logic; attribute dont_touch of I30629: signal is true;
	signal I30634: std_logic; attribute dont_touch of I30634: signal is true;
	signal I30635: std_logic; attribute dont_touch of I30635: signal is true;
	signal I30636: std_logic; attribute dont_touch of I30636: signal is true;
	signal I30641: std_logic; attribute dont_touch of I30641: signal is true;
	signal I30642: std_logic; attribute dont_touch of I30642: signal is true;
	signal I30643: std_logic; attribute dont_touch of I30643: signal is true;
	signal I30644: std_logic; attribute dont_touch of I30644: signal is true;
	signal I30645: std_logic; attribute dont_touch of I30645: signal is true;
	signal I30650: std_logic; attribute dont_touch of I30650: signal is true;
	signal I30651: std_logic; attribute dont_touch of I30651: signal is true;
	signal I30652: std_logic; attribute dont_touch of I30652: signal is true;
	signal I30657: std_logic; attribute dont_touch of I30657: signal is true;
	signal I30658: std_logic; attribute dont_touch of I30658: signal is true;
	signal I30659: std_logic; attribute dont_touch of I30659: signal is true;
	signal I30660: std_logic; attribute dont_touch of I30660: signal is true;
	signal I30665: std_logic; attribute dont_touch of I30665: signal is true;
	signal I30666: std_logic; attribute dont_touch of I30666: signal is true;
	signal I30667: std_logic; attribute dont_touch of I30667: signal is true;
	signal I30672: std_logic; attribute dont_touch of I30672: signal is true;
	signal I30673: std_logic; attribute dont_touch of I30673: signal is true;
	signal I30674: std_logic; attribute dont_touch of I30674: signal is true;
	signal I30675: std_logic; attribute dont_touch of I30675: signal is true;
	signal I30676: std_logic; attribute dont_touch of I30676: signal is true;
	signal I30681: std_logic; attribute dont_touch of I30681: signal is true;
	signal I30682: std_logic; attribute dont_touch of I30682: signal is true;
	signal I30683: std_logic; attribute dont_touch of I30683: signal is true;
	signal I30688: std_logic; attribute dont_touch of I30688: signal is true;
	signal I30689: std_logic; attribute dont_touch of I30689: signal is true;
	signal I30690: std_logic; attribute dont_touch of I30690: signal is true;
	signal I30691: std_logic; attribute dont_touch of I30691: signal is true;
	signal I30696: std_logic; attribute dont_touch of I30696: signal is true;
	signal I30697: std_logic; attribute dont_touch of I30697: signal is true;
	signal I30698: std_logic; attribute dont_touch of I30698: signal is true;
	signal I30703: std_logic; attribute dont_touch of I30703: signal is true;
	signal I30704: std_logic; attribute dont_touch of I30704: signal is true;
	signal I30705: std_logic; attribute dont_touch of I30705: signal is true;
	signal I30706: std_logic; attribute dont_touch of I30706: signal is true;
	signal I30707: std_logic; attribute dont_touch of I30707: signal is true;
	signal I30712: std_logic; attribute dont_touch of I30712: signal is true;
	signal I30713: std_logic; attribute dont_touch of I30713: signal is true;
	signal I30714: std_logic; attribute dont_touch of I30714: signal is true;
	signal I30719: std_logic; attribute dont_touch of I30719: signal is true;
	signal I30720: std_logic; attribute dont_touch of I30720: signal is true;
	signal I30721: std_logic; attribute dont_touch of I30721: signal is true;
	signal I30722: std_logic; attribute dont_touch of I30722: signal is true;
	signal I30727: std_logic; attribute dont_touch of I30727: signal is true;
	signal I30728: std_logic; attribute dont_touch of I30728: signal is true;
	signal I30729: std_logic; attribute dont_touch of I30729: signal is true;
	signal I30734: std_logic; attribute dont_touch of I30734: signal is true;
	signal I30735: std_logic; attribute dont_touch of I30735: signal is true;
	signal I30736: std_logic; attribute dont_touch of I30736: signal is true;
	signal I30737: std_logic; attribute dont_touch of I30737: signal is true;
	signal I30738: std_logic; attribute dont_touch of I30738: signal is true;
	signal I30743: std_logic; attribute dont_touch of I30743: signal is true;
	signal I30744: std_logic; attribute dont_touch of I30744: signal is true;
	signal I30745: std_logic; attribute dont_touch of I30745: signal is true;
	signal I30750: std_logic; attribute dont_touch of I30750: signal is true;
	signal I30751: std_logic; attribute dont_touch of I30751: signal is true;
	signal I30752: std_logic; attribute dont_touch of I30752: signal is true;
	signal I30753: std_logic; attribute dont_touch of I30753: signal is true;
	signal I30758: std_logic; attribute dont_touch of I30758: signal is true;
	signal I30759: std_logic; attribute dont_touch of I30759: signal is true;
	signal I30760: std_logic; attribute dont_touch of I30760: signal is true;
	signal I30765: std_logic; attribute dont_touch of I30765: signal is true;
	signal I30766: std_logic; attribute dont_touch of I30766: signal is true;
	signal I30767: std_logic; attribute dont_touch of I30767: signal is true;
	signal I30768: std_logic; attribute dont_touch of I30768: signal is true;
	signal I30769: std_logic; attribute dont_touch of I30769: signal is true;
	signal I30774: std_logic; attribute dont_touch of I30774: signal is true;
	signal I30775: std_logic; attribute dont_touch of I30775: signal is true;
	signal I30776: std_logic; attribute dont_touch of I30776: signal is true;
	signal I30781: std_logic; attribute dont_touch of I30781: signal is true;
	signal I30782: std_logic; attribute dont_touch of I30782: signal is true;
	signal I30783: std_logic; attribute dont_touch of I30783: signal is true;
	signal I30784: std_logic; attribute dont_touch of I30784: signal is true;
	signal I30789: std_logic; attribute dont_touch of I30789: signal is true;
	signal I30790: std_logic; attribute dont_touch of I30790: signal is true;
	signal I30791: std_logic; attribute dont_touch of I30791: signal is true;
	signal I30796: std_logic; attribute dont_touch of I30796: signal is true;
	signal I30797: std_logic; attribute dont_touch of I30797: signal is true;
	signal I30798: std_logic; attribute dont_touch of I30798: signal is true;
	signal I30799: std_logic; attribute dont_touch of I30799: signal is true;
	signal I30800: std_logic; attribute dont_touch of I30800: signal is true;
	signal I30805: std_logic; attribute dont_touch of I30805: signal is true;
	signal I30806: std_logic; attribute dont_touch of I30806: signal is true;
	signal I30807: std_logic; attribute dont_touch of I30807: signal is true;
	signal I30812: std_logic; attribute dont_touch of I30812: signal is true;
	signal I30813: std_logic; attribute dont_touch of I30813: signal is true;
	signal I30814: std_logic; attribute dont_touch of I30814: signal is true;
	signal I30815: std_logic; attribute dont_touch of I30815: signal is true;
	signal I30820: std_logic; attribute dont_touch of I30820: signal is true;
	signal I30821: std_logic; attribute dont_touch of I30821: signal is true;
	signal I30822: std_logic; attribute dont_touch of I30822: signal is true;
	signal I30827: std_logic; attribute dont_touch of I30827: signal is true;
	signal I30828: std_logic; attribute dont_touch of I30828: signal is true;
	signal I30829: std_logic; attribute dont_touch of I30829: signal is true;
	signal I30830: std_logic; attribute dont_touch of I30830: signal is true;
	signal I30831: std_logic; attribute dont_touch of I30831: signal is true;
	signal I30836: std_logic; attribute dont_touch of I30836: signal is true;
	signal I30837: std_logic; attribute dont_touch of I30837: signal is true;
	signal I30838: std_logic; attribute dont_touch of I30838: signal is true;
	signal I30843: std_logic; attribute dont_touch of I30843: signal is true;
	signal I30844: std_logic; attribute dont_touch of I30844: signal is true;
	signal I30845: std_logic; attribute dont_touch of I30845: signal is true;
	signal I30846: std_logic; attribute dont_touch of I30846: signal is true;
	signal I30851: std_logic; attribute dont_touch of I30851: signal is true;
	signal I30852: std_logic; attribute dont_touch of I30852: signal is true;
	signal I30853: std_logic; attribute dont_touch of I30853: signal is true;
	signal I30858: std_logic; attribute dont_touch of I30858: signal is true;
	signal I30859: std_logic; attribute dont_touch of I30859: signal is true;
	signal I30860: std_logic; attribute dont_touch of I30860: signal is true;
	signal I30861: std_logic; attribute dont_touch of I30861: signal is true;
	signal I30862: std_logic; attribute dont_touch of I30862: signal is true;
	signal I30867: std_logic; attribute dont_touch of I30867: signal is true;
	signal I30868: std_logic; attribute dont_touch of I30868: signal is true;
	signal I30869: std_logic; attribute dont_touch of I30869: signal is true;
	signal I30874: std_logic; attribute dont_touch of I30874: signal is true;
	signal I30875: std_logic; attribute dont_touch of I30875: signal is true;
	signal I30876: std_logic; attribute dont_touch of I30876: signal is true;
	signal I30877: std_logic; attribute dont_touch of I30877: signal is true;
	signal I30882: std_logic; attribute dont_touch of I30882: signal is true;
	signal I30883: std_logic; attribute dont_touch of I30883: signal is true;
	signal I30884: std_logic; attribute dont_touch of I30884: signal is true;
	signal I30889: std_logic; attribute dont_touch of I30889: signal is true;
	signal I30890: std_logic; attribute dont_touch of I30890: signal is true;
	signal I30891: std_logic; attribute dont_touch of I30891: signal is true;
	signal I30892: std_logic; attribute dont_touch of I30892: signal is true;
	signal I30893: std_logic; attribute dont_touch of I30893: signal is true;
	signal I30898: std_logic; attribute dont_touch of I30898: signal is true;
	signal I30899: std_logic; attribute dont_touch of I30899: signal is true;
	signal I30900: std_logic; attribute dont_touch of I30900: signal is true;
	signal I30905: std_logic; attribute dont_touch of I30905: signal is true;
	signal I30906: std_logic; attribute dont_touch of I30906: signal is true;
	signal I30907: std_logic; attribute dont_touch of I30907: signal is true;
	signal I30908: std_logic; attribute dont_touch of I30908: signal is true;
	signal I30913: std_logic; attribute dont_touch of I30913: signal is true;
	signal I30914: std_logic; attribute dont_touch of I30914: signal is true;
	signal I30915: std_logic; attribute dont_touch of I30915: signal is true;
	signal I30920: std_logic; attribute dont_touch of I30920: signal is true;
	signal I30921: std_logic; attribute dont_touch of I30921: signal is true;
	signal I30922: std_logic; attribute dont_touch of I30922: signal is true;
	signal I30923: std_logic; attribute dont_touch of I30923: signal is true;
	signal I30924: std_logic; attribute dont_touch of I30924: signal is true;
	signal I30929: std_logic; attribute dont_touch of I30929: signal is true;
	signal I30930: std_logic; attribute dont_touch of I30930: signal is true;
	signal I30931: std_logic; attribute dont_touch of I30931: signal is true;
	signal I30936: std_logic; attribute dont_touch of I30936: signal is true;
	signal I30937: std_logic; attribute dont_touch of I30937: signal is true;
	signal I30938: std_logic; attribute dont_touch of I30938: signal is true;
	signal I30939: std_logic; attribute dont_touch of I30939: signal is true;
	signal I30944: std_logic; attribute dont_touch of I30944: signal is true;
	signal I30945: std_logic; attribute dont_touch of I30945: signal is true;
	signal I30946: std_logic; attribute dont_touch of I30946: signal is true;
	signal I30951: std_logic; attribute dont_touch of I30951: signal is true;
	signal I30952: std_logic; attribute dont_touch of I30952: signal is true;
	signal I30953: std_logic; attribute dont_touch of I30953: signal is true;
	signal I30954: std_logic; attribute dont_touch of I30954: signal is true;
	signal I30955: std_logic; attribute dont_touch of I30955: signal is true;
	signal I30960: std_logic; attribute dont_touch of I30960: signal is true;
	signal I30961: std_logic; attribute dont_touch of I30961: signal is true;
	signal I30962: std_logic; attribute dont_touch of I30962: signal is true;
	signal I30967: std_logic; attribute dont_touch of I30967: signal is true;
	signal I30968: std_logic; attribute dont_touch of I30968: signal is true;
	signal I30969: std_logic; attribute dont_touch of I30969: signal is true;
	signal I30970: std_logic; attribute dont_touch of I30970: signal is true;
	signal I30975: std_logic; attribute dont_touch of I30975: signal is true;
	signal I30976: std_logic; attribute dont_touch of I30976: signal is true;
	signal I30977: std_logic; attribute dont_touch of I30977: signal is true;
	signal I30982: std_logic; attribute dont_touch of I30982: signal is true;
	signal I30983: std_logic; attribute dont_touch of I30983: signal is true;
	signal I30984: std_logic; attribute dont_touch of I30984: signal is true;
	signal I30985: std_logic; attribute dont_touch of I30985: signal is true;
	signal I30986: std_logic; attribute dont_touch of I30986: signal is true;
	signal I30991: std_logic; attribute dont_touch of I30991: signal is true;
	signal I30992: std_logic; attribute dont_touch of I30992: signal is true;
	signal I30993: std_logic; attribute dont_touch of I30993: signal is true;
	signal I30998: std_logic; attribute dont_touch of I30998: signal is true;
	signal I30999: std_logic; attribute dont_touch of I30999: signal is true;
	signal I31000: std_logic; attribute dont_touch of I31000: signal is true;
	signal I31001: std_logic; attribute dont_touch of I31001: signal is true;
	signal I31006: std_logic; attribute dont_touch of I31006: signal is true;
	signal I31007: std_logic; attribute dont_touch of I31007: signal is true;
	signal I31008: std_logic; attribute dont_touch of I31008: signal is true;
	signal I31087: std_logic; attribute dont_touch of I31087: signal is true;
	signal I31088: std_logic; attribute dont_touch of I31088: signal is true;
	signal I31089: std_logic; attribute dont_touch of I31089: signal is true;
	signal I31100: std_logic; attribute dont_touch of I31100: signal is true;
	signal I31101: std_logic; attribute dont_touch of I31101: signal is true;
	signal I31102: std_logic; attribute dont_touch of I31102: signal is true;
	signal I31113: std_logic; attribute dont_touch of I31113: signal is true;
	signal I31114: std_logic; attribute dont_touch of I31114: signal is true;
	signal I31115: std_logic; attribute dont_touch of I31115: signal is true;
	signal I31126: std_logic; attribute dont_touch of I31126: signal is true;
	signal I31127: std_logic; attribute dont_touch of I31127: signal is true;
	signal I31128: std_logic; attribute dont_touch of I31128: signal is true;
	signal I31139: std_logic; attribute dont_touch of I31139: signal is true;
	signal I31140: std_logic; attribute dont_touch of I31140: signal is true;
	signal I31141: std_logic; attribute dont_touch of I31141: signal is true;
	signal I31152: std_logic; attribute dont_touch of I31152: signal is true;
	signal I31153: std_logic; attribute dont_touch of I31153: signal is true;
	signal I31154: std_logic; attribute dont_touch of I31154: signal is true;
	signal I31165: std_logic; attribute dont_touch of I31165: signal is true;
	signal I31166: std_logic; attribute dont_touch of I31166: signal is true;
	signal I31167: std_logic; attribute dont_touch of I31167: signal is true;
	signal I31178: std_logic; attribute dont_touch of I31178: signal is true;
	signal I31179: std_logic; attribute dont_touch of I31179: signal is true;
	signal I31180: std_logic; attribute dont_touch of I31180: signal is true;
	signal I31191: std_logic; attribute dont_touch of I31191: signal is true;
	signal I31192: std_logic; attribute dont_touch of I31192: signal is true;
	signal I31193: std_logic; attribute dont_touch of I31193: signal is true;
	signal I31204: std_logic; attribute dont_touch of I31204: signal is true;
	signal I31205: std_logic; attribute dont_touch of I31205: signal is true;
	signal I31206: std_logic; attribute dont_touch of I31206: signal is true;
	signal I31217: std_logic; attribute dont_touch of I31217: signal is true;
	signal I31218: std_logic; attribute dont_touch of I31218: signal is true;
	signal I31219: std_logic; attribute dont_touch of I31219: signal is true;
	signal I31230: std_logic; attribute dont_touch of I31230: signal is true;
	signal I31231: std_logic; attribute dont_touch of I31231: signal is true;
	signal I31232: std_logic; attribute dont_touch of I31232: signal is true;
	signal I31243: std_logic; attribute dont_touch of I31243: signal is true;
	signal I31244: std_logic; attribute dont_touch of I31244: signal is true;
	signal I31245: std_logic; attribute dont_touch of I31245: signal is true;
	signal I31256: std_logic; attribute dont_touch of I31256: signal is true;
	signal I31257: std_logic; attribute dont_touch of I31257: signal is true;
	signal I31258: std_logic; attribute dont_touch of I31258: signal is true;
	signal I31269: std_logic; attribute dont_touch of I31269: signal is true;
	signal I31270: std_logic; attribute dont_touch of I31270: signal is true;
	signal I31271: std_logic; attribute dont_touch of I31271: signal is true;
	signal I31282: std_logic; attribute dont_touch of I31282: signal is true;
	signal I31283: std_logic; attribute dont_touch of I31283: signal is true;
	signal I31284: std_logic; attribute dont_touch of I31284: signal is true;
	signal I31295: std_logic; attribute dont_touch of I31295: signal is true;
	signal I31296: std_logic; attribute dont_touch of I31296: signal is true;
	signal I31297: std_logic; attribute dont_touch of I31297: signal is true;
	signal I31308: std_logic; attribute dont_touch of I31308: signal is true;
	signal I31309: std_logic; attribute dont_touch of I31309: signal is true;
	signal I31310: std_logic; attribute dont_touch of I31310: signal is true;
	signal I31321: std_logic; attribute dont_touch of I31321: signal is true;
	signal I31322: std_logic; attribute dont_touch of I31322: signal is true;
	signal I31323: std_logic; attribute dont_touch of I31323: signal is true;
	signal I31334: std_logic; attribute dont_touch of I31334: signal is true;
	signal I31335: std_logic; attribute dont_touch of I31335: signal is true;
	signal I31336: std_logic; attribute dont_touch of I31336: signal is true;
	signal I31347: std_logic; attribute dont_touch of I31347: signal is true;
	signal I31348: std_logic; attribute dont_touch of I31348: signal is true;
	signal I31349: std_logic; attribute dont_touch of I31349: signal is true;
	signal I31360: std_logic; attribute dont_touch of I31360: signal is true;
	signal I31361: std_logic; attribute dont_touch of I31361: signal is true;
	signal I31362: std_logic; attribute dont_touch of I31362: signal is true;
	signal I31373: std_logic; attribute dont_touch of I31373: signal is true;
	signal I31374: std_logic; attribute dont_touch of I31374: signal is true;
	signal I31375: std_logic; attribute dont_touch of I31375: signal is true;
	signal I31386: std_logic; attribute dont_touch of I31386: signal is true;
	signal I31387: std_logic; attribute dont_touch of I31387: signal is true;
	signal I31388: std_logic; attribute dont_touch of I31388: signal is true;
	signal I31399: std_logic; attribute dont_touch of I31399: signal is true;
	signal I31400: std_logic; attribute dont_touch of I31400: signal is true;
	signal I31401: std_logic; attribute dont_touch of I31401: signal is true;
	signal I31412: std_logic; attribute dont_touch of I31412: signal is true;
	signal I31413: std_logic; attribute dont_touch of I31413: signal is true;
	signal I31414: std_logic; attribute dont_touch of I31414: signal is true;
	signal I31425: std_logic; attribute dont_touch of I31425: signal is true;
	signal I31426: std_logic; attribute dont_touch of I31426: signal is true;
	signal I31427: std_logic; attribute dont_touch of I31427: signal is true;
	signal I31438: std_logic; attribute dont_touch of I31438: signal is true;
	signal I31439: std_logic; attribute dont_touch of I31439: signal is true;
	signal I31440: std_logic; attribute dont_touch of I31440: signal is true;
	signal I31451: std_logic; attribute dont_touch of I31451: signal is true;
	signal I31452: std_logic; attribute dont_touch of I31452: signal is true;
	signal I31453: std_logic; attribute dont_touch of I31453: signal is true;
	signal I31464: std_logic; attribute dont_touch of I31464: signal is true;
	signal I31465: std_logic; attribute dont_touch of I31465: signal is true;
	signal I31466: std_logic; attribute dont_touch of I31466: signal is true;
	signal I31477: std_logic; attribute dont_touch of I31477: signal is true;
	signal I31478: std_logic; attribute dont_touch of I31478: signal is true;
	signal I31479: std_logic; attribute dont_touch of I31479: signal is true;
	signal I31490: std_logic; attribute dont_touch of I31490: signal is true;
	signal I31491: std_logic; attribute dont_touch of I31491: signal is true;
	signal I31492: std_logic; attribute dont_touch of I31492: signal is true;
	signal I31504: std_logic; attribute dont_touch of I31504: signal is true;
	signal I31505: std_logic; attribute dont_touch of I31505: signal is true;
	signal I31506: std_logic; attribute dont_touch of I31506: signal is true;
	signal I31507: std_logic; attribute dont_touch of I31507: signal is true;
	signal I31512: std_logic; attribute dont_touch of I31512: signal is true;
	signal I31513: std_logic; attribute dont_touch of I31513: signal is true;
	signal I31514: std_logic; attribute dont_touch of I31514: signal is true;
	signal I31519: std_logic; attribute dont_touch of I31519: signal is true;
	signal I31520: std_logic; attribute dont_touch of I31520: signal is true;
	signal I31521: std_logic; attribute dont_touch of I31521: signal is true;
	signal I31522: std_logic; attribute dont_touch of I31522: signal is true;
	signal I31527: std_logic; attribute dont_touch of I31527: signal is true;
	signal I31528: std_logic; attribute dont_touch of I31528: signal is true;
	signal I31529: std_logic; attribute dont_touch of I31529: signal is true;
	signal I31534: std_logic; attribute dont_touch of I31534: signal is true;
	signal I31535: std_logic; attribute dont_touch of I31535: signal is true;
	signal I31536: std_logic; attribute dont_touch of I31536: signal is true;
	signal I31537: std_logic; attribute dont_touch of I31537: signal is true;
	signal I31542: std_logic; attribute dont_touch of I31542: signal is true;
	signal I31543: std_logic; attribute dont_touch of I31543: signal is true;
	signal I31544: std_logic; attribute dont_touch of I31544: signal is true;
	signal I31549: std_logic; attribute dont_touch of I31549: signal is true;
	signal I31550: std_logic; attribute dont_touch of I31550: signal is true;
	signal I31551: std_logic; attribute dont_touch of I31551: signal is true;
	signal I31556: std_logic; attribute dont_touch of I31556: signal is true;
	signal I31557: std_logic; attribute dont_touch of I31557: signal is true;
	signal I31558: std_logic; attribute dont_touch of I31558: signal is true;
	signal I31563: std_logic; attribute dont_touch of I31563: signal is true;
	signal I31564: std_logic; attribute dont_touch of I31564: signal is true;
	signal I31565: std_logic; attribute dont_touch of I31565: signal is true;
	signal I31570: std_logic; attribute dont_touch of I31570: signal is true;
	signal I31571: std_logic; attribute dont_touch of I31571: signal is true;
	signal I31572: std_logic; attribute dont_touch of I31572: signal is true;
	signal I31577: std_logic; attribute dont_touch of I31577: signal is true;
	signal I31578: std_logic; attribute dont_touch of I31578: signal is true;
	signal I31579: std_logic; attribute dont_touch of I31579: signal is true;
	signal I31584: std_logic; attribute dont_touch of I31584: signal is true;
	signal I31585: std_logic; attribute dont_touch of I31585: signal is true;
	signal I31586: std_logic; attribute dont_touch of I31586: signal is true;
	signal I31591: std_logic; attribute dont_touch of I31591: signal is true;
	signal I31592: std_logic; attribute dont_touch of I31592: signal is true;
	signal I31593: std_logic; attribute dont_touch of I31593: signal is true;
	signal I31598: std_logic; attribute dont_touch of I31598: signal is true;
	signal I31599: std_logic; attribute dont_touch of I31599: signal is true;
	signal I31600: std_logic; attribute dont_touch of I31600: signal is true;
	signal I31605: std_logic; attribute dont_touch of I31605: signal is true;
	signal I31606: std_logic; attribute dont_touch of I31606: signal is true;
	signal I31607: std_logic; attribute dont_touch of I31607: signal is true;
	signal I31612: std_logic; attribute dont_touch of I31612: signal is true;
	signal I31613: std_logic; attribute dont_touch of I31613: signal is true;
	signal I31614: std_logic; attribute dont_touch of I31614: signal is true;
	signal I31619: std_logic; attribute dont_touch of I31619: signal is true;
	signal I31620: std_logic; attribute dont_touch of I31620: signal is true;
	signal I31621: std_logic; attribute dont_touch of I31621: signal is true;
	signal I31626: std_logic; attribute dont_touch of I31626: signal is true;
	signal I31627: std_logic; attribute dont_touch of I31627: signal is true;
	signal I31628: std_logic; attribute dont_touch of I31628: signal is true;
	signal I31633: std_logic; attribute dont_touch of I31633: signal is true;
	signal I31634: std_logic; attribute dont_touch of I31634: signal is true;
	signal I31635: std_logic; attribute dont_touch of I31635: signal is true;
	signal I31640: std_logic; attribute dont_touch of I31640: signal is true;
	signal I31641: std_logic; attribute dont_touch of I31641: signal is true;
	signal I31642: std_logic; attribute dont_touch of I31642: signal is true;
	signal I31647: std_logic; attribute dont_touch of I31647: signal is true;
	signal I31648: std_logic; attribute dont_touch of I31648: signal is true;
	signal I31649: std_logic; attribute dont_touch of I31649: signal is true;
	signal I31654: std_logic; attribute dont_touch of I31654: signal is true;
	signal I31655: std_logic; attribute dont_touch of I31655: signal is true;
	signal I31656: std_logic; attribute dont_touch of I31656: signal is true;
	signal I31661: std_logic; attribute dont_touch of I31661: signal is true;
	signal I31662: std_logic; attribute dont_touch of I31662: signal is true;
	signal I31663: std_logic; attribute dont_touch of I31663: signal is true;
	signal I31668: std_logic; attribute dont_touch of I31668: signal is true;
	signal I31669: std_logic; attribute dont_touch of I31669: signal is true;
	signal I31670: std_logic; attribute dont_touch of I31670: signal is true;
	signal I31675: std_logic; attribute dont_touch of I31675: signal is true;
	signal I31676: std_logic; attribute dont_touch of I31676: signal is true;
	signal I31677: std_logic; attribute dont_touch of I31677: signal is true;
	signal I31682: std_logic; attribute dont_touch of I31682: signal is true;
	signal I31683: std_logic; attribute dont_touch of I31683: signal is true;
	signal I31684: std_logic; attribute dont_touch of I31684: signal is true;
	signal I31689: std_logic; attribute dont_touch of I31689: signal is true;
	signal I31690: std_logic; attribute dont_touch of I31690: signal is true;
	signal I31691: std_logic; attribute dont_touch of I31691: signal is true;
	signal I31696: std_logic; attribute dont_touch of I31696: signal is true;
	signal I31697: std_logic; attribute dont_touch of I31697: signal is true;
	signal I31698: std_logic; attribute dont_touch of I31698: signal is true;
	signal I31703: std_logic; attribute dont_touch of I31703: signal is true;
	signal I31704: std_logic; attribute dont_touch of I31704: signal is true;
	signal I31705: std_logic; attribute dont_touch of I31705: signal is true;
	signal I31710: std_logic; attribute dont_touch of I31710: signal is true;
	signal I31711: std_logic; attribute dont_touch of I31711: signal is true;
	signal I31712: std_logic; attribute dont_touch of I31712: signal is true;
	signal I31717: std_logic; attribute dont_touch of I31717: signal is true;
	signal I31718: std_logic; attribute dont_touch of I31718: signal is true;
	signal I31719: std_logic; attribute dont_touch of I31719: signal is true;
	signal I31724: std_logic; attribute dont_touch of I31724: signal is true;
	signal I31725: std_logic; attribute dont_touch of I31725: signal is true;
	signal I31726: std_logic; attribute dont_touch of I31726: signal is true;
	signal I31731: std_logic; attribute dont_touch of I31731: signal is true;
	signal I31732: std_logic; attribute dont_touch of I31732: signal is true;
	signal I31733: std_logic; attribute dont_touch of I31733: signal is true;
	signal I31738: std_logic; attribute dont_touch of I31738: signal is true;
	signal I31739: std_logic; attribute dont_touch of I31739: signal is true;
	signal I31740: std_logic; attribute dont_touch of I31740: signal is true;
	signal I31745: std_logic; attribute dont_touch of I31745: signal is true;
	signal I31746: std_logic; attribute dont_touch of I31746: signal is true;
	signal I31747: std_logic; attribute dont_touch of I31747: signal is true;
	signal I34026: std_logic; attribute dont_touch of I34026: signal is true;
	signal I34027: std_logic; attribute dont_touch of I34027: signal is true;
	signal I34028: std_logic; attribute dont_touch of I34028: signal is true;
	signal I34029: std_logic; attribute dont_touch of I34029: signal is true;
	signal I34030: std_logic; attribute dont_touch of I34030: signal is true;
	signal I34035: std_logic; attribute dont_touch of I34035: signal is true;
	signal I34036: std_logic; attribute dont_touch of I34036: signal is true;
	signal I34037: std_logic; attribute dont_touch of I34037: signal is true;
	signal I34042: std_logic; attribute dont_touch of I34042: signal is true;
	signal I34043: std_logic; attribute dont_touch of I34043: signal is true;
	signal I34044: std_logic; attribute dont_touch of I34044: signal is true;
	signal I34045: std_logic; attribute dont_touch of I34045: signal is true;
	signal I34050: std_logic; attribute dont_touch of I34050: signal is true;
	signal I34051: std_logic; attribute dont_touch of I34051: signal is true;
	signal I34052: std_logic; attribute dont_touch of I34052: signal is true;
	signal I34057: std_logic; attribute dont_touch of I34057: signal is true;
	signal I34058: std_logic; attribute dont_touch of I34058: signal is true;
	signal I34059: std_logic; attribute dont_touch of I34059: signal is true;
	signal I34060: std_logic; attribute dont_touch of I34060: signal is true;
	signal I34061: std_logic; attribute dont_touch of I34061: signal is true;
	signal I34066: std_logic; attribute dont_touch of I34066: signal is true;
	signal I34067: std_logic; attribute dont_touch of I34067: signal is true;
	signal I34068: std_logic; attribute dont_touch of I34068: signal is true;
	signal I34073: std_logic; attribute dont_touch of I34073: signal is true;
	signal I34074: std_logic; attribute dont_touch of I34074: signal is true;
	signal I34075: std_logic; attribute dont_touch of I34075: signal is true;
	signal I34076: std_logic; attribute dont_touch of I34076: signal is true;
	signal I34081: std_logic; attribute dont_touch of I34081: signal is true;
	signal I34082: std_logic; attribute dont_touch of I34082: signal is true;
	signal I34083: std_logic; attribute dont_touch of I34083: signal is true;
	signal I34088: std_logic; attribute dont_touch of I34088: signal is true;
	signal I34089: std_logic; attribute dont_touch of I34089: signal is true;
	signal I34090: std_logic; attribute dont_touch of I34090: signal is true;
	signal I34091: std_logic; attribute dont_touch of I34091: signal is true;
	signal I34092: std_logic; attribute dont_touch of I34092: signal is true;
	signal I34097: std_logic; attribute dont_touch of I34097: signal is true;
	signal I34098: std_logic; attribute dont_touch of I34098: signal is true;
	signal I34099: std_logic; attribute dont_touch of I34099: signal is true;
	signal I34104: std_logic; attribute dont_touch of I34104: signal is true;
	signal I34105: std_logic; attribute dont_touch of I34105: signal is true;
	signal I34106: std_logic; attribute dont_touch of I34106: signal is true;
	signal I34107: std_logic; attribute dont_touch of I34107: signal is true;
	signal I34112: std_logic; attribute dont_touch of I34112: signal is true;
	signal I34113: std_logic; attribute dont_touch of I34113: signal is true;
	signal I34114: std_logic; attribute dont_touch of I34114: signal is true;
	signal I34119: std_logic; attribute dont_touch of I34119: signal is true;
	signal I34120: std_logic; attribute dont_touch of I34120: signal is true;
	signal I34121: std_logic; attribute dont_touch of I34121: signal is true;
	signal I34122: std_logic; attribute dont_touch of I34122: signal is true;
	signal I34123: std_logic; attribute dont_touch of I34123: signal is true;
	signal I34128: std_logic; attribute dont_touch of I34128: signal is true;
	signal I34129: std_logic; attribute dont_touch of I34129: signal is true;
	signal I34130: std_logic; attribute dont_touch of I34130: signal is true;
	signal I34135: std_logic; attribute dont_touch of I34135: signal is true;
	signal I34136: std_logic; attribute dont_touch of I34136: signal is true;
	signal I34137: std_logic; attribute dont_touch of I34137: signal is true;
	signal I34138: std_logic; attribute dont_touch of I34138: signal is true;
	signal I34143: std_logic; attribute dont_touch of I34143: signal is true;
	signal I34144: std_logic; attribute dont_touch of I34144: signal is true;
	signal I34145: std_logic; attribute dont_touch of I34145: signal is true;
	signal I34150: std_logic; attribute dont_touch of I34150: signal is true;
	signal I34151: std_logic; attribute dont_touch of I34151: signal is true;
	signal I34152: std_logic; attribute dont_touch of I34152: signal is true;
	signal I34153: std_logic; attribute dont_touch of I34153: signal is true;
	signal I34154: std_logic; attribute dont_touch of I34154: signal is true;
	signal I34159: std_logic; attribute dont_touch of I34159: signal is true;
	signal I34160: std_logic; attribute dont_touch of I34160: signal is true;
	signal I34161: std_logic; attribute dont_touch of I34161: signal is true;
	signal I34166: std_logic; attribute dont_touch of I34166: signal is true;
	signal I34167: std_logic; attribute dont_touch of I34167: signal is true;
	signal I34168: std_logic; attribute dont_touch of I34168: signal is true;
	signal I34169: std_logic; attribute dont_touch of I34169: signal is true;
	signal I34174: std_logic; attribute dont_touch of I34174: signal is true;
	signal I34175: std_logic; attribute dont_touch of I34175: signal is true;
	signal I34176: std_logic; attribute dont_touch of I34176: signal is true;
	signal I34181: std_logic; attribute dont_touch of I34181: signal is true;
	signal I34182: std_logic; attribute dont_touch of I34182: signal is true;
	signal I34183: std_logic; attribute dont_touch of I34183: signal is true;
	signal I34184: std_logic; attribute dont_touch of I34184: signal is true;
	signal I34185: std_logic; attribute dont_touch of I34185: signal is true;
	signal I34190: std_logic; attribute dont_touch of I34190: signal is true;
	signal I34191: std_logic; attribute dont_touch of I34191: signal is true;
	signal I34192: std_logic; attribute dont_touch of I34192: signal is true;
	signal I34197: std_logic; attribute dont_touch of I34197: signal is true;
	signal I34198: std_logic; attribute dont_touch of I34198: signal is true;
	signal I34199: std_logic; attribute dont_touch of I34199: signal is true;
	signal I34200: std_logic; attribute dont_touch of I34200: signal is true;
	signal I34205: std_logic; attribute dont_touch of I34205: signal is true;
	signal I34206: std_logic; attribute dont_touch of I34206: signal is true;
	signal I34207: std_logic; attribute dont_touch of I34207: signal is true;
	signal I34212: std_logic; attribute dont_touch of I34212: signal is true;
	signal I34213: std_logic; attribute dont_touch of I34213: signal is true;
	signal I34214: std_logic; attribute dont_touch of I34214: signal is true;
	signal I34215: std_logic; attribute dont_touch of I34215: signal is true;
	signal I34216: std_logic; attribute dont_touch of I34216: signal is true;
	signal I34221: std_logic; attribute dont_touch of I34221: signal is true;
	signal I34222: std_logic; attribute dont_touch of I34222: signal is true;
	signal I34223: std_logic; attribute dont_touch of I34223: signal is true;
	signal I34228: std_logic; attribute dont_touch of I34228: signal is true;
	signal I34229: std_logic; attribute dont_touch of I34229: signal is true;
	signal I34230: std_logic; attribute dont_touch of I34230: signal is true;
	signal I34231: std_logic; attribute dont_touch of I34231: signal is true;
	signal I34236: std_logic; attribute dont_touch of I34236: signal is true;
	signal I34237: std_logic; attribute dont_touch of I34237: signal is true;
	signal I34238: std_logic; attribute dont_touch of I34238: signal is true;
	signal I34243: std_logic; attribute dont_touch of I34243: signal is true;
	signal I34244: std_logic; attribute dont_touch of I34244: signal is true;
	signal I34245: std_logic; attribute dont_touch of I34245: signal is true;
	signal I34246: std_logic; attribute dont_touch of I34246: signal is true;
	signal I34247: std_logic; attribute dont_touch of I34247: signal is true;
	signal I34252: std_logic; attribute dont_touch of I34252: signal is true;
	signal I34253: std_logic; attribute dont_touch of I34253: signal is true;
	signal I34254: std_logic; attribute dont_touch of I34254: signal is true;
	signal I34259: std_logic; attribute dont_touch of I34259: signal is true;
	signal I34260: std_logic; attribute dont_touch of I34260: signal is true;
	signal I34261: std_logic; attribute dont_touch of I34261: signal is true;
	signal I34262: std_logic; attribute dont_touch of I34262: signal is true;
	signal I34267: std_logic; attribute dont_touch of I34267: signal is true;
	signal I34268: std_logic; attribute dont_touch of I34268: signal is true;
	signal I34269: std_logic; attribute dont_touch of I34269: signal is true;
	signal I34274: std_logic; attribute dont_touch of I34274: signal is true;
	signal I34275: std_logic; attribute dont_touch of I34275: signal is true;
	signal I34276: std_logic; attribute dont_touch of I34276: signal is true;
	signal I34277: std_logic; attribute dont_touch of I34277: signal is true;
	signal I34278: std_logic; attribute dont_touch of I34278: signal is true;
	signal I34283: std_logic; attribute dont_touch of I34283: signal is true;
	signal I34284: std_logic; attribute dont_touch of I34284: signal is true;
	signal I34285: std_logic; attribute dont_touch of I34285: signal is true;
	signal I34290: std_logic; attribute dont_touch of I34290: signal is true;
	signal I34291: std_logic; attribute dont_touch of I34291: signal is true;
	signal I34292: std_logic; attribute dont_touch of I34292: signal is true;
	signal I34293: std_logic; attribute dont_touch of I34293: signal is true;
	signal I34298: std_logic; attribute dont_touch of I34298: signal is true;
	signal I34299: std_logic; attribute dont_touch of I34299: signal is true;
	signal I34300: std_logic; attribute dont_touch of I34300: signal is true;
	signal I34305: std_logic; attribute dont_touch of I34305: signal is true;
	signal I34306: std_logic; attribute dont_touch of I34306: signal is true;
	signal I34307: std_logic; attribute dont_touch of I34307: signal is true;
	signal I34308: std_logic; attribute dont_touch of I34308: signal is true;
	signal I34309: std_logic; attribute dont_touch of I34309: signal is true;
	signal I34314: std_logic; attribute dont_touch of I34314: signal is true;
	signal I34315: std_logic; attribute dont_touch of I34315: signal is true;
	signal I34316: std_logic; attribute dont_touch of I34316: signal is true;
	signal I34321: std_logic; attribute dont_touch of I34321: signal is true;
	signal I34322: std_logic; attribute dont_touch of I34322: signal is true;
	signal I34323: std_logic; attribute dont_touch of I34323: signal is true;
	signal I34324: std_logic; attribute dont_touch of I34324: signal is true;
	signal I34329: std_logic; attribute dont_touch of I34329: signal is true;
	signal I34330: std_logic; attribute dont_touch of I34330: signal is true;
	signal I34331: std_logic; attribute dont_touch of I34331: signal is true;
	signal I34336: std_logic; attribute dont_touch of I34336: signal is true;
	signal I34337: std_logic; attribute dont_touch of I34337: signal is true;
	signal I34338: std_logic; attribute dont_touch of I34338: signal is true;
	signal I34339: std_logic; attribute dont_touch of I34339: signal is true;
	signal I34340: std_logic; attribute dont_touch of I34340: signal is true;
	signal I34345: std_logic; attribute dont_touch of I34345: signal is true;
	signal I34346: std_logic; attribute dont_touch of I34346: signal is true;
	signal I34347: std_logic; attribute dont_touch of I34347: signal is true;
	signal I34352: std_logic; attribute dont_touch of I34352: signal is true;
	signal I34353: std_logic; attribute dont_touch of I34353: signal is true;
	signal I34354: std_logic; attribute dont_touch of I34354: signal is true;
	signal I34355: std_logic; attribute dont_touch of I34355: signal is true;
	signal I34360: std_logic; attribute dont_touch of I34360: signal is true;
	signal I34361: std_logic; attribute dont_touch of I34361: signal is true;
	signal I34362: std_logic; attribute dont_touch of I34362: signal is true;
	signal I34367: std_logic; attribute dont_touch of I34367: signal is true;
	signal I34368: std_logic; attribute dont_touch of I34368: signal is true;
	signal I34369: std_logic; attribute dont_touch of I34369: signal is true;
	signal I34370: std_logic; attribute dont_touch of I34370: signal is true;
	signal I34371: std_logic; attribute dont_touch of I34371: signal is true;
	signal I34376: std_logic; attribute dont_touch of I34376: signal is true;
	signal I34377: std_logic; attribute dont_touch of I34377: signal is true;
	signal I34378: std_logic; attribute dont_touch of I34378: signal is true;
	signal I34383: std_logic; attribute dont_touch of I34383: signal is true;
	signal I34384: std_logic; attribute dont_touch of I34384: signal is true;
	signal I34385: std_logic; attribute dont_touch of I34385: signal is true;
	signal I34386: std_logic; attribute dont_touch of I34386: signal is true;
	signal I34391: std_logic; attribute dont_touch of I34391: signal is true;
	signal I34392: std_logic; attribute dont_touch of I34392: signal is true;
	signal I34393: std_logic; attribute dont_touch of I34393: signal is true;
	signal I34398: std_logic; attribute dont_touch of I34398: signal is true;
	signal I34399: std_logic; attribute dont_touch of I34399: signal is true;
	signal I34400: std_logic; attribute dont_touch of I34400: signal is true;
	signal I34401: std_logic; attribute dont_touch of I34401: signal is true;
	signal I34402: std_logic; attribute dont_touch of I34402: signal is true;
	signal I34407: std_logic; attribute dont_touch of I34407: signal is true;
	signal I34408: std_logic; attribute dont_touch of I34408: signal is true;
	signal I34409: std_logic; attribute dont_touch of I34409: signal is true;
	signal I34414: std_logic; attribute dont_touch of I34414: signal is true;
	signal I34415: std_logic; attribute dont_touch of I34415: signal is true;
	signal I34416: std_logic; attribute dont_touch of I34416: signal is true;
	signal I34417: std_logic; attribute dont_touch of I34417: signal is true;
	signal I34422: std_logic; attribute dont_touch of I34422: signal is true;
	signal I34423: std_logic; attribute dont_touch of I34423: signal is true;
	signal I34424: std_logic; attribute dont_touch of I34424: signal is true;
	signal I34429: std_logic; attribute dont_touch of I34429: signal is true;
	signal I34430: std_logic; attribute dont_touch of I34430: signal is true;
	signal I34431: std_logic; attribute dont_touch of I34431: signal is true;
	signal I34432: std_logic; attribute dont_touch of I34432: signal is true;
	signal I34433: std_logic; attribute dont_touch of I34433: signal is true;
	signal I34438: std_logic; attribute dont_touch of I34438: signal is true;
	signal I34439: std_logic; attribute dont_touch of I34439: signal is true;
	signal I34440: std_logic; attribute dont_touch of I34440: signal is true;
	signal I34445: std_logic; attribute dont_touch of I34445: signal is true;
	signal I34446: std_logic; attribute dont_touch of I34446: signal is true;
	signal I34447: std_logic; attribute dont_touch of I34447: signal is true;
	signal I34448: std_logic; attribute dont_touch of I34448: signal is true;
	signal I34453: std_logic; attribute dont_touch of I34453: signal is true;
	signal I34454: std_logic; attribute dont_touch of I34454: signal is true;
	signal I34455: std_logic; attribute dont_touch of I34455: signal is true;
	signal I34460: std_logic; attribute dont_touch of I34460: signal is true;
	signal I34461: std_logic; attribute dont_touch of I34461: signal is true;
	signal I34462: std_logic; attribute dont_touch of I34462: signal is true;
	signal I34463: std_logic; attribute dont_touch of I34463: signal is true;
	signal I34464: std_logic; attribute dont_touch of I34464: signal is true;
	signal I34469: std_logic; attribute dont_touch of I34469: signal is true;
	signal I34470: std_logic; attribute dont_touch of I34470: signal is true;
	signal I34471: std_logic; attribute dont_touch of I34471: signal is true;
	signal I34476: std_logic; attribute dont_touch of I34476: signal is true;
	signal I34477: std_logic; attribute dont_touch of I34477: signal is true;
	signal I34478: std_logic; attribute dont_touch of I34478: signal is true;
	signal I34479: std_logic; attribute dont_touch of I34479: signal is true;
	signal I34484: std_logic; attribute dont_touch of I34484: signal is true;
	signal I34485: std_logic; attribute dont_touch of I34485: signal is true;
	signal I34486: std_logic; attribute dont_touch of I34486: signal is true;
	signal I34491: std_logic; attribute dont_touch of I34491: signal is true;
	signal I34492: std_logic; attribute dont_touch of I34492: signal is true;
	signal I34493: std_logic; attribute dont_touch of I34493: signal is true;
	signal I34494: std_logic; attribute dont_touch of I34494: signal is true;
	signal I34495: std_logic; attribute dont_touch of I34495: signal is true;
	signal I34500: std_logic; attribute dont_touch of I34500: signal is true;
	signal I34501: std_logic; attribute dont_touch of I34501: signal is true;
	signal I34502: std_logic; attribute dont_touch of I34502: signal is true;
	signal I34507: std_logic; attribute dont_touch of I34507: signal is true;
	signal I34508: std_logic; attribute dont_touch of I34508: signal is true;
	signal I34509: std_logic; attribute dont_touch of I34509: signal is true;
	signal I34510: std_logic; attribute dont_touch of I34510: signal is true;
	signal I34515: std_logic; attribute dont_touch of I34515: signal is true;
	signal I34516: std_logic; attribute dont_touch of I34516: signal is true;
	signal I34517: std_logic; attribute dont_touch of I34517: signal is true;
	signal I34522: std_logic; attribute dont_touch of I34522: signal is true;
	signal I34523: std_logic; attribute dont_touch of I34523: signal is true;
	signal I34524: std_logic; attribute dont_touch of I34524: signal is true;
	signal I34525: std_logic; attribute dont_touch of I34525: signal is true;
	signal I34526: std_logic; attribute dont_touch of I34526: signal is true;
	signal I34531: std_logic; attribute dont_touch of I34531: signal is true;
	signal I34532: std_logic; attribute dont_touch of I34532: signal is true;
	signal I34533: std_logic; attribute dont_touch of I34533: signal is true;
	signal I34538: std_logic; attribute dont_touch of I34538: signal is true;
	signal I34539: std_logic; attribute dont_touch of I34539: signal is true;
	signal I34540: std_logic; attribute dont_touch of I34540: signal is true;
	signal I34541: std_logic; attribute dont_touch of I34541: signal is true;
	signal I34546: std_logic; attribute dont_touch of I34546: signal is true;
	signal I34547: std_logic; attribute dont_touch of I34547: signal is true;
	signal I34548: std_logic; attribute dont_touch of I34548: signal is true;
	signal I34553: std_logic; attribute dont_touch of I34553: signal is true;
	signal I34554: std_logic; attribute dont_touch of I34554: signal is true;
	signal I34555: std_logic; attribute dont_touch of I34555: signal is true;
	signal I34556: std_logic; attribute dont_touch of I34556: signal is true;
	signal I34557: std_logic; attribute dont_touch of I34557: signal is true;
	signal I34562: std_logic; attribute dont_touch of I34562: signal is true;
	signal I34563: std_logic; attribute dont_touch of I34563: signal is true;
	signal I34564: std_logic; attribute dont_touch of I34564: signal is true;
	signal I34569: std_logic; attribute dont_touch of I34569: signal is true;
	signal I34570: std_logic; attribute dont_touch of I34570: signal is true;
	signal I34571: std_logic; attribute dont_touch of I34571: signal is true;
	signal I34572: std_logic; attribute dont_touch of I34572: signal is true;
	signal I34577: std_logic; attribute dont_touch of I34577: signal is true;
	signal I34578: std_logic; attribute dont_touch of I34578: signal is true;
	signal I34579: std_logic; attribute dont_touch of I34579: signal is true;
	signal I34584: std_logic; attribute dont_touch of I34584: signal is true;
	signal I34585: std_logic; attribute dont_touch of I34585: signal is true;
	signal I34586: std_logic; attribute dont_touch of I34586: signal is true;
	signal I34587: std_logic; attribute dont_touch of I34587: signal is true;
	signal I34588: std_logic; attribute dont_touch of I34588: signal is true;
	signal I34593: std_logic; attribute dont_touch of I34593: signal is true;
	signal I34594: std_logic; attribute dont_touch of I34594: signal is true;
	signal I34595: std_logic; attribute dont_touch of I34595: signal is true;
	signal I34600: std_logic; attribute dont_touch of I34600: signal is true;
	signal I34601: std_logic; attribute dont_touch of I34601: signal is true;
	signal I34602: std_logic; attribute dont_touch of I34602: signal is true;
	signal I34603: std_logic; attribute dont_touch of I34603: signal is true;
	signal I34608: std_logic; attribute dont_touch of I34608: signal is true;
	signal I34609: std_logic; attribute dont_touch of I34609: signal is true;
	signal I34610: std_logic; attribute dont_touch of I34610: signal is true;
	signal I34615: std_logic; attribute dont_touch of I34615: signal is true;
	signal I34616: std_logic; attribute dont_touch of I34616: signal is true;
	signal I34617: std_logic; attribute dont_touch of I34617: signal is true;
	signal I34618: std_logic; attribute dont_touch of I34618: signal is true;
	signal I34619: std_logic; attribute dont_touch of I34619: signal is true;
	signal I34624: std_logic; attribute dont_touch of I34624: signal is true;
	signal I34625: std_logic; attribute dont_touch of I34625: signal is true;
	signal I34626: std_logic; attribute dont_touch of I34626: signal is true;
	signal I34631: std_logic; attribute dont_touch of I34631: signal is true;
	signal I34632: std_logic; attribute dont_touch of I34632: signal is true;
	signal I34633: std_logic; attribute dont_touch of I34633: signal is true;
	signal I34634: std_logic; attribute dont_touch of I34634: signal is true;
	signal I34639: std_logic; attribute dont_touch of I34639: signal is true;
	signal I34640: std_logic; attribute dont_touch of I34640: signal is true;
	signal I34641: std_logic; attribute dont_touch of I34641: signal is true;
	signal I34646: std_logic; attribute dont_touch of I34646: signal is true;
	signal I34647: std_logic; attribute dont_touch of I34647: signal is true;
	signal I34648: std_logic; attribute dont_touch of I34648: signal is true;
	signal I34649: std_logic; attribute dont_touch of I34649: signal is true;
	signal I34650: std_logic; attribute dont_touch of I34650: signal is true;
	signal I34655: std_logic; attribute dont_touch of I34655: signal is true;
	signal I34656: std_logic; attribute dont_touch of I34656: signal is true;
	signal I34657: std_logic; attribute dont_touch of I34657: signal is true;
	signal I34662: std_logic; attribute dont_touch of I34662: signal is true;
	signal I34663: std_logic; attribute dont_touch of I34663: signal is true;
	signal I34664: std_logic; attribute dont_touch of I34664: signal is true;
	signal I34665: std_logic; attribute dont_touch of I34665: signal is true;
	signal I34670: std_logic; attribute dont_touch of I34670: signal is true;
	signal I34671: std_logic; attribute dont_touch of I34671: signal is true;
	signal I34672: std_logic; attribute dont_touch of I34672: signal is true;
	signal I34677: std_logic; attribute dont_touch of I34677: signal is true;
	signal I34678: std_logic; attribute dont_touch of I34678: signal is true;
	signal I34679: std_logic; attribute dont_touch of I34679: signal is true;
	signal I34680: std_logic; attribute dont_touch of I34680: signal is true;
	signal I34681: std_logic; attribute dont_touch of I34681: signal is true;
	signal I34686: std_logic; attribute dont_touch of I34686: signal is true;
	signal I34687: std_logic; attribute dont_touch of I34687: signal is true;
	signal I34688: std_logic; attribute dont_touch of I34688: signal is true;
	signal I34693: std_logic; attribute dont_touch of I34693: signal is true;
	signal I34694: std_logic; attribute dont_touch of I34694: signal is true;
	signal I34695: std_logic; attribute dont_touch of I34695: signal is true;
	signal I34696: std_logic; attribute dont_touch of I34696: signal is true;
	signal I34701: std_logic; attribute dont_touch of I34701: signal is true;
	signal I34702: std_logic; attribute dont_touch of I34702: signal is true;
	signal I34703: std_logic; attribute dont_touch of I34703: signal is true;
	signal I34708: std_logic; attribute dont_touch of I34708: signal is true;
	signal I34709: std_logic; attribute dont_touch of I34709: signal is true;
	signal I34710: std_logic; attribute dont_touch of I34710: signal is true;
	signal I34711: std_logic; attribute dont_touch of I34711: signal is true;
	signal I34712: std_logic; attribute dont_touch of I34712: signal is true;
	signal I34717: std_logic; attribute dont_touch of I34717: signal is true;
	signal I34718: std_logic; attribute dont_touch of I34718: signal is true;
	signal I34719: std_logic; attribute dont_touch of I34719: signal is true;
	signal I34724: std_logic; attribute dont_touch of I34724: signal is true;
	signal I34725: std_logic; attribute dont_touch of I34725: signal is true;
	signal I34726: std_logic; attribute dont_touch of I34726: signal is true;
	signal I34727: std_logic; attribute dont_touch of I34727: signal is true;
	signal I34732: std_logic; attribute dont_touch of I34732: signal is true;
	signal I34733: std_logic; attribute dont_touch of I34733: signal is true;
	signal I34734: std_logic; attribute dont_touch of I34734: signal is true;
	signal I34739: std_logic; attribute dont_touch of I34739: signal is true;
	signal I34740: std_logic; attribute dont_touch of I34740: signal is true;
	signal I34741: std_logic; attribute dont_touch of I34741: signal is true;
	signal I34742: std_logic; attribute dont_touch of I34742: signal is true;
	signal I34743: std_logic; attribute dont_touch of I34743: signal is true;
	signal I34748: std_logic; attribute dont_touch of I34748: signal is true;
	signal I34749: std_logic; attribute dont_touch of I34749: signal is true;
	signal I34750: std_logic; attribute dont_touch of I34750: signal is true;
	signal I34755: std_logic; attribute dont_touch of I34755: signal is true;
	signal I34756: std_logic; attribute dont_touch of I34756: signal is true;
	signal I34757: std_logic; attribute dont_touch of I34757: signal is true;
	signal I34758: std_logic; attribute dont_touch of I34758: signal is true;
	signal I34763: std_logic; attribute dont_touch of I34763: signal is true;
	signal I34764: std_logic; attribute dont_touch of I34764: signal is true;
	signal I34765: std_logic; attribute dont_touch of I34765: signal is true;
	signal I34770: std_logic; attribute dont_touch of I34770: signal is true;
	signal I34771: std_logic; attribute dont_touch of I34771: signal is true;
	signal I34772: std_logic; attribute dont_touch of I34772: signal is true;
	signal I34773: std_logic; attribute dont_touch of I34773: signal is true;
	signal I34774: std_logic; attribute dont_touch of I34774: signal is true;
	signal I34779: std_logic; attribute dont_touch of I34779: signal is true;
	signal I34780: std_logic; attribute dont_touch of I34780: signal is true;
	signal I34781: std_logic; attribute dont_touch of I34781: signal is true;
	signal I34786: std_logic; attribute dont_touch of I34786: signal is true;
	signal I34787: std_logic; attribute dont_touch of I34787: signal is true;
	signal I34788: std_logic; attribute dont_touch of I34788: signal is true;
	signal I34789: std_logic; attribute dont_touch of I34789: signal is true;
	signal I34794: std_logic; attribute dont_touch of I34794: signal is true;
	signal I34795: std_logic; attribute dont_touch of I34795: signal is true;
	signal I34796: std_logic; attribute dont_touch of I34796: signal is true;
	signal I34801: std_logic; attribute dont_touch of I34801: signal is true;
	signal I34802: std_logic; attribute dont_touch of I34802: signal is true;
	signal I34803: std_logic; attribute dont_touch of I34803: signal is true;
	signal I34804: std_logic; attribute dont_touch of I34804: signal is true;
	signal I34805: std_logic; attribute dont_touch of I34805: signal is true;
	signal I34810: std_logic; attribute dont_touch of I34810: signal is true;
	signal I34811: std_logic; attribute dont_touch of I34811: signal is true;
	signal I34812: std_logic; attribute dont_touch of I34812: signal is true;
	signal I34817: std_logic; attribute dont_touch of I34817: signal is true;
	signal I34818: std_logic; attribute dont_touch of I34818: signal is true;
	signal I34819: std_logic; attribute dont_touch of I34819: signal is true;
	signal I34820: std_logic; attribute dont_touch of I34820: signal is true;
	signal I34825: std_logic; attribute dont_touch of I34825: signal is true;
	signal I34826: std_logic; attribute dont_touch of I34826: signal is true;
	signal I34827: std_logic; attribute dont_touch of I34827: signal is true;
	signal I34832: std_logic; attribute dont_touch of I34832: signal is true;
	signal I34833: std_logic; attribute dont_touch of I34833: signal is true;
	signal I34834: std_logic; attribute dont_touch of I34834: signal is true;
	signal I34835: std_logic; attribute dont_touch of I34835: signal is true;
	signal I34836: std_logic; attribute dont_touch of I34836: signal is true;
	signal I34841: std_logic; attribute dont_touch of I34841: signal is true;
	signal I34842: std_logic; attribute dont_touch of I34842: signal is true;
	signal I34843: std_logic; attribute dont_touch of I34843: signal is true;
	signal I34848: std_logic; attribute dont_touch of I34848: signal is true;
	signal I34849: std_logic; attribute dont_touch of I34849: signal is true;
	signal I34850: std_logic; attribute dont_touch of I34850: signal is true;
	signal I34851: std_logic; attribute dont_touch of I34851: signal is true;
	signal I34856: std_logic; attribute dont_touch of I34856: signal is true;
	signal I34857: std_logic; attribute dont_touch of I34857: signal is true;
	signal I34858: std_logic; attribute dont_touch of I34858: signal is true;
	signal I34863: std_logic; attribute dont_touch of I34863: signal is true;
	signal I34864: std_logic; attribute dont_touch of I34864: signal is true;
	signal I34865: std_logic; attribute dont_touch of I34865: signal is true;
	signal I34866: std_logic; attribute dont_touch of I34866: signal is true;
	signal I34867: std_logic; attribute dont_touch of I34867: signal is true;
	signal I34872: std_logic; attribute dont_touch of I34872: signal is true;
	signal I34873: std_logic; attribute dont_touch of I34873: signal is true;
	signal I34874: std_logic; attribute dont_touch of I34874: signal is true;
	signal I34879: std_logic; attribute dont_touch of I34879: signal is true;
	signal I34880: std_logic; attribute dont_touch of I34880: signal is true;
	signal I34881: std_logic; attribute dont_touch of I34881: signal is true;
	signal I34882: std_logic; attribute dont_touch of I34882: signal is true;
	signal I34887: std_logic; attribute dont_touch of I34887: signal is true;
	signal I34888: std_logic; attribute dont_touch of I34888: signal is true;
	signal I34889: std_logic; attribute dont_touch of I34889: signal is true;
	signal I34894: std_logic; attribute dont_touch of I34894: signal is true;
	signal I34895: std_logic; attribute dont_touch of I34895: signal is true;
	signal I34896: std_logic; attribute dont_touch of I34896: signal is true;
	signal I34897: std_logic; attribute dont_touch of I34897: signal is true;
	signal I34898: std_logic; attribute dont_touch of I34898: signal is true;
	signal I34903: std_logic; attribute dont_touch of I34903: signal is true;
	signal I34904: std_logic; attribute dont_touch of I34904: signal is true;
	signal I34905: std_logic; attribute dont_touch of I34905: signal is true;
	signal I34910: std_logic; attribute dont_touch of I34910: signal is true;
	signal I34911: std_logic; attribute dont_touch of I34911: signal is true;
	signal I34912: std_logic; attribute dont_touch of I34912: signal is true;
	signal I34913: std_logic; attribute dont_touch of I34913: signal is true;
	signal I34918: std_logic; attribute dont_touch of I34918: signal is true;
	signal I34919: std_logic; attribute dont_touch of I34919: signal is true;
	signal I34920: std_logic; attribute dont_touch of I34920: signal is true;
	signal I34925: std_logic; attribute dont_touch of I34925: signal is true;
	signal I34926: std_logic; attribute dont_touch of I34926: signal is true;
	signal I34927: std_logic; attribute dont_touch of I34927: signal is true;
	signal I34928: std_logic; attribute dont_touch of I34928: signal is true;
	signal I34929: std_logic; attribute dont_touch of I34929: signal is true;
	signal I34934: std_logic; attribute dont_touch of I34934: signal is true;
	signal I34935: std_logic; attribute dont_touch of I34935: signal is true;
	signal I34936: std_logic; attribute dont_touch of I34936: signal is true;
	signal I34941: std_logic; attribute dont_touch of I34941: signal is true;
	signal I34942: std_logic; attribute dont_touch of I34942: signal is true;
	signal I34943: std_logic; attribute dont_touch of I34943: signal is true;
	signal I34944: std_logic; attribute dont_touch of I34944: signal is true;
	signal I34949: std_logic; attribute dont_touch of I34949: signal is true;
	signal I34950: std_logic; attribute dont_touch of I34950: signal is true;
	signal I34951: std_logic; attribute dont_touch of I34951: signal is true;
	signal I34956: std_logic; attribute dont_touch of I34956: signal is true;
	signal I34957: std_logic; attribute dont_touch of I34957: signal is true;
	signal I34958: std_logic; attribute dont_touch of I34958: signal is true;
	signal I34959: std_logic; attribute dont_touch of I34959: signal is true;
	signal I34960: std_logic; attribute dont_touch of I34960: signal is true;
	signal I34965: std_logic; attribute dont_touch of I34965: signal is true;
	signal I34966: std_logic; attribute dont_touch of I34966: signal is true;
	signal I34967: std_logic; attribute dont_touch of I34967: signal is true;
	signal I34972: std_logic; attribute dont_touch of I34972: signal is true;
	signal I34973: std_logic; attribute dont_touch of I34973: signal is true;
	signal I34974: std_logic; attribute dont_touch of I34974: signal is true;
	signal I34975: std_logic; attribute dont_touch of I34975: signal is true;
	signal I34980: std_logic; attribute dont_touch of I34980: signal is true;
	signal I34981: std_logic; attribute dont_touch of I34981: signal is true;
	signal I34982: std_logic; attribute dont_touch of I34982: signal is true;
	signal I34987: std_logic; attribute dont_touch of I34987: signal is true;
	signal I34988: std_logic; attribute dont_touch of I34988: signal is true;
	signal I34989: std_logic; attribute dont_touch of I34989: signal is true;
	signal I34990: std_logic; attribute dont_touch of I34990: signal is true;
	signal I34991: std_logic; attribute dont_touch of I34991: signal is true;
	signal I34996: std_logic; attribute dont_touch of I34996: signal is true;
	signal I34997: std_logic; attribute dont_touch of I34997: signal is true;
	signal I34998: std_logic; attribute dont_touch of I34998: signal is true;
	signal I35003: std_logic; attribute dont_touch of I35003: signal is true;
	signal I35004: std_logic; attribute dont_touch of I35004: signal is true;
	signal I35005: std_logic; attribute dont_touch of I35005: signal is true;
	signal I35006: std_logic; attribute dont_touch of I35006: signal is true;
	signal I35011: std_logic; attribute dont_touch of I35011: signal is true;
	signal I35012: std_logic; attribute dont_touch of I35012: signal is true;
	signal I35013: std_logic; attribute dont_touch of I35013: signal is true;
	signal I35092: std_logic; attribute dont_touch of I35092: signal is true;
	signal I35093: std_logic; attribute dont_touch of I35093: signal is true;
	signal I35094: std_logic; attribute dont_touch of I35094: signal is true;
	signal I35105: std_logic; attribute dont_touch of I35105: signal is true;
	signal I35106: std_logic; attribute dont_touch of I35106: signal is true;
	signal I35107: std_logic; attribute dont_touch of I35107: signal is true;
	signal I35118: std_logic; attribute dont_touch of I35118: signal is true;
	signal I35119: std_logic; attribute dont_touch of I35119: signal is true;
	signal I35120: std_logic; attribute dont_touch of I35120: signal is true;
	signal I35131: std_logic; attribute dont_touch of I35131: signal is true;
	signal I35132: std_logic; attribute dont_touch of I35132: signal is true;
	signal I35133: std_logic; attribute dont_touch of I35133: signal is true;
	signal I35144: std_logic; attribute dont_touch of I35144: signal is true;
	signal I35145: std_logic; attribute dont_touch of I35145: signal is true;
	signal I35146: std_logic; attribute dont_touch of I35146: signal is true;
	signal I35157: std_logic; attribute dont_touch of I35157: signal is true;
	signal I35158: std_logic; attribute dont_touch of I35158: signal is true;
	signal I35159: std_logic; attribute dont_touch of I35159: signal is true;
	signal I35170: std_logic; attribute dont_touch of I35170: signal is true;
	signal I35171: std_logic; attribute dont_touch of I35171: signal is true;
	signal I35172: std_logic; attribute dont_touch of I35172: signal is true;
	signal I35183: std_logic; attribute dont_touch of I35183: signal is true;
	signal I35184: std_logic; attribute dont_touch of I35184: signal is true;
	signal I35185: std_logic; attribute dont_touch of I35185: signal is true;
	signal I35196: std_logic; attribute dont_touch of I35196: signal is true;
	signal I35197: std_logic; attribute dont_touch of I35197: signal is true;
	signal I35198: std_logic; attribute dont_touch of I35198: signal is true;
	signal I35209: std_logic; attribute dont_touch of I35209: signal is true;
	signal I35210: std_logic; attribute dont_touch of I35210: signal is true;
	signal I35211: std_logic; attribute dont_touch of I35211: signal is true;
	signal I35222: std_logic; attribute dont_touch of I35222: signal is true;
	signal I35223: std_logic; attribute dont_touch of I35223: signal is true;
	signal I35224: std_logic; attribute dont_touch of I35224: signal is true;
	signal I35235: std_logic; attribute dont_touch of I35235: signal is true;
	signal I35236: std_logic; attribute dont_touch of I35236: signal is true;
	signal I35237: std_logic; attribute dont_touch of I35237: signal is true;
	signal I35248: std_logic; attribute dont_touch of I35248: signal is true;
	signal I35249: std_logic; attribute dont_touch of I35249: signal is true;
	signal I35250: std_logic; attribute dont_touch of I35250: signal is true;
	signal I35261: std_logic; attribute dont_touch of I35261: signal is true;
	signal I35262: std_logic; attribute dont_touch of I35262: signal is true;
	signal I35263: std_logic; attribute dont_touch of I35263: signal is true;
	signal I35274: std_logic; attribute dont_touch of I35274: signal is true;
	signal I35275: std_logic; attribute dont_touch of I35275: signal is true;
	signal I35276: std_logic; attribute dont_touch of I35276: signal is true;
	signal I35287: std_logic; attribute dont_touch of I35287: signal is true;
	signal I35288: std_logic; attribute dont_touch of I35288: signal is true;
	signal I35289: std_logic; attribute dont_touch of I35289: signal is true;
	signal I35300: std_logic; attribute dont_touch of I35300: signal is true;
	signal I35301: std_logic; attribute dont_touch of I35301: signal is true;
	signal I35302: std_logic; attribute dont_touch of I35302: signal is true;
	signal I35313: std_logic; attribute dont_touch of I35313: signal is true;
	signal I35314: std_logic; attribute dont_touch of I35314: signal is true;
	signal I35315: std_logic; attribute dont_touch of I35315: signal is true;
	signal I35326: std_logic; attribute dont_touch of I35326: signal is true;
	signal I35327: std_logic; attribute dont_touch of I35327: signal is true;
	signal I35328: std_logic; attribute dont_touch of I35328: signal is true;
	signal I35339: std_logic; attribute dont_touch of I35339: signal is true;
	signal I35340: std_logic; attribute dont_touch of I35340: signal is true;
	signal I35341: std_logic; attribute dont_touch of I35341: signal is true;
	signal I35352: std_logic; attribute dont_touch of I35352: signal is true;
	signal I35353: std_logic; attribute dont_touch of I35353: signal is true;
	signal I35354: std_logic; attribute dont_touch of I35354: signal is true;
	signal I35365: std_logic; attribute dont_touch of I35365: signal is true;
	signal I35366: std_logic; attribute dont_touch of I35366: signal is true;
	signal I35367: std_logic; attribute dont_touch of I35367: signal is true;
	signal I35378: std_logic; attribute dont_touch of I35378: signal is true;
	signal I35379: std_logic; attribute dont_touch of I35379: signal is true;
	signal I35380: std_logic; attribute dont_touch of I35380: signal is true;
	signal I35391: std_logic; attribute dont_touch of I35391: signal is true;
	signal I35392: std_logic; attribute dont_touch of I35392: signal is true;
	signal I35393: std_logic; attribute dont_touch of I35393: signal is true;
	signal I35404: std_logic; attribute dont_touch of I35404: signal is true;
	signal I35405: std_logic; attribute dont_touch of I35405: signal is true;
	signal I35406: std_logic; attribute dont_touch of I35406: signal is true;
	signal I35417: std_logic; attribute dont_touch of I35417: signal is true;
	signal I35418: std_logic; attribute dont_touch of I35418: signal is true;
	signal I35419: std_logic; attribute dont_touch of I35419: signal is true;
	signal I35430: std_logic; attribute dont_touch of I35430: signal is true;
	signal I35431: std_logic; attribute dont_touch of I35431: signal is true;
	signal I35432: std_logic; attribute dont_touch of I35432: signal is true;
	signal I35443: std_logic; attribute dont_touch of I35443: signal is true;
	signal I35444: std_logic; attribute dont_touch of I35444: signal is true;
	signal I35445: std_logic; attribute dont_touch of I35445: signal is true;
	signal I35456: std_logic; attribute dont_touch of I35456: signal is true;
	signal I35457: std_logic; attribute dont_touch of I35457: signal is true;
	signal I35458: std_logic; attribute dont_touch of I35458: signal is true;
	signal I35469: std_logic; attribute dont_touch of I35469: signal is true;
	signal I35470: std_logic; attribute dont_touch of I35470: signal is true;
	signal I35471: std_logic; attribute dont_touch of I35471: signal is true;
	signal I35482: std_logic; attribute dont_touch of I35482: signal is true;
	signal I35483: std_logic; attribute dont_touch of I35483: signal is true;
	signal I35484: std_logic; attribute dont_touch of I35484: signal is true;
	signal I35495: std_logic; attribute dont_touch of I35495: signal is true;
	signal I35496: std_logic; attribute dont_touch of I35496: signal is true;
	signal I35497: std_logic; attribute dont_touch of I35497: signal is true;
	signal I35509: std_logic; attribute dont_touch of I35509: signal is true;
	signal I35510: std_logic; attribute dont_touch of I35510: signal is true;
	signal I35511: std_logic; attribute dont_touch of I35511: signal is true;
	signal I35512: std_logic; attribute dont_touch of I35512: signal is true;
	signal I35517: std_logic; attribute dont_touch of I35517: signal is true;
	signal I35518: std_logic; attribute dont_touch of I35518: signal is true;
	signal I35519: std_logic; attribute dont_touch of I35519: signal is true;
	signal I35524: std_logic; attribute dont_touch of I35524: signal is true;
	signal I35525: std_logic; attribute dont_touch of I35525: signal is true;
	signal I35526: std_logic; attribute dont_touch of I35526: signal is true;
	signal I35527: std_logic; attribute dont_touch of I35527: signal is true;
	signal I35532: std_logic; attribute dont_touch of I35532: signal is true;
	signal I35533: std_logic; attribute dont_touch of I35533: signal is true;
	signal I35534: std_logic; attribute dont_touch of I35534: signal is true;
	signal I35539: std_logic; attribute dont_touch of I35539: signal is true;
	signal I35540: std_logic; attribute dont_touch of I35540: signal is true;
	signal I35541: std_logic; attribute dont_touch of I35541: signal is true;
	signal I35542: std_logic; attribute dont_touch of I35542: signal is true;
	signal I35547: std_logic; attribute dont_touch of I35547: signal is true;
	signal I35548: std_logic; attribute dont_touch of I35548: signal is true;
	signal I35549: std_logic; attribute dont_touch of I35549: signal is true;
	signal I35554: std_logic; attribute dont_touch of I35554: signal is true;
	signal I35555: std_logic; attribute dont_touch of I35555: signal is true;
	signal I35556: std_logic; attribute dont_touch of I35556: signal is true;
	signal I35561: std_logic; attribute dont_touch of I35561: signal is true;
	signal I35562: std_logic; attribute dont_touch of I35562: signal is true;
	signal I35563: std_logic; attribute dont_touch of I35563: signal is true;
	signal I35568: std_logic; attribute dont_touch of I35568: signal is true;
	signal I35569: std_logic; attribute dont_touch of I35569: signal is true;
	signal I35570: std_logic; attribute dont_touch of I35570: signal is true;
	signal I35575: std_logic; attribute dont_touch of I35575: signal is true;
	signal I35576: std_logic; attribute dont_touch of I35576: signal is true;
	signal I35577: std_logic; attribute dont_touch of I35577: signal is true;
	signal I35582: std_logic; attribute dont_touch of I35582: signal is true;
	signal I35583: std_logic; attribute dont_touch of I35583: signal is true;
	signal I35584: std_logic; attribute dont_touch of I35584: signal is true;
	signal I35589: std_logic; attribute dont_touch of I35589: signal is true;
	signal I35590: std_logic; attribute dont_touch of I35590: signal is true;
	signal I35591: std_logic; attribute dont_touch of I35591: signal is true;
	signal I35596: std_logic; attribute dont_touch of I35596: signal is true;
	signal I35597: std_logic; attribute dont_touch of I35597: signal is true;
	signal I35598: std_logic; attribute dont_touch of I35598: signal is true;
	signal I35603: std_logic; attribute dont_touch of I35603: signal is true;
	signal I35604: std_logic; attribute dont_touch of I35604: signal is true;
	signal I35605: std_logic; attribute dont_touch of I35605: signal is true;
	signal I35610: std_logic; attribute dont_touch of I35610: signal is true;
	signal I35611: std_logic; attribute dont_touch of I35611: signal is true;
	signal I35612: std_logic; attribute dont_touch of I35612: signal is true;
	signal I35617: std_logic; attribute dont_touch of I35617: signal is true;
	signal I35618: std_logic; attribute dont_touch of I35618: signal is true;
	signal I35619: std_logic; attribute dont_touch of I35619: signal is true;
	signal I35624: std_logic; attribute dont_touch of I35624: signal is true;
	signal I35625: std_logic; attribute dont_touch of I35625: signal is true;
	signal I35626: std_logic; attribute dont_touch of I35626: signal is true;
	signal I35631: std_logic; attribute dont_touch of I35631: signal is true;
	signal I35632: std_logic; attribute dont_touch of I35632: signal is true;
	signal I35633: std_logic; attribute dont_touch of I35633: signal is true;
	signal I35638: std_logic; attribute dont_touch of I35638: signal is true;
	signal I35639: std_logic; attribute dont_touch of I35639: signal is true;
	signal I35640: std_logic; attribute dont_touch of I35640: signal is true;
	signal I35645: std_logic; attribute dont_touch of I35645: signal is true;
	signal I35646: std_logic; attribute dont_touch of I35646: signal is true;
	signal I35647: std_logic; attribute dont_touch of I35647: signal is true;
	signal I35652: std_logic; attribute dont_touch of I35652: signal is true;
	signal I35653: std_logic; attribute dont_touch of I35653: signal is true;
	signal I35654: std_logic; attribute dont_touch of I35654: signal is true;
	signal I35659: std_logic; attribute dont_touch of I35659: signal is true;
	signal I35660: std_logic; attribute dont_touch of I35660: signal is true;
	signal I35661: std_logic; attribute dont_touch of I35661: signal is true;
	signal I35666: std_logic; attribute dont_touch of I35666: signal is true;
	signal I35667: std_logic; attribute dont_touch of I35667: signal is true;
	signal I35668: std_logic; attribute dont_touch of I35668: signal is true;
	signal I35673: std_logic; attribute dont_touch of I35673: signal is true;
	signal I35674: std_logic; attribute dont_touch of I35674: signal is true;
	signal I35675: std_logic; attribute dont_touch of I35675: signal is true;
	signal I35680: std_logic; attribute dont_touch of I35680: signal is true;
	signal I35681: std_logic; attribute dont_touch of I35681: signal is true;
	signal I35682: std_logic; attribute dont_touch of I35682: signal is true;
	signal I35687: std_logic; attribute dont_touch of I35687: signal is true;
	signal I35688: std_logic; attribute dont_touch of I35688: signal is true;
	signal I35689: std_logic; attribute dont_touch of I35689: signal is true;
	signal I35694: std_logic; attribute dont_touch of I35694: signal is true;
	signal I35695: std_logic; attribute dont_touch of I35695: signal is true;
	signal I35696: std_logic; attribute dont_touch of I35696: signal is true;
	signal I35701: std_logic; attribute dont_touch of I35701: signal is true;
	signal I35702: std_logic; attribute dont_touch of I35702: signal is true;
	signal I35703: std_logic; attribute dont_touch of I35703: signal is true;
	signal I35708: std_logic; attribute dont_touch of I35708: signal is true;
	signal I35709: std_logic; attribute dont_touch of I35709: signal is true;
	signal I35710: std_logic; attribute dont_touch of I35710: signal is true;
	signal I35715: std_logic; attribute dont_touch of I35715: signal is true;
	signal I35716: std_logic; attribute dont_touch of I35716: signal is true;
	signal I35717: std_logic; attribute dont_touch of I35717: signal is true;
	signal I35722: std_logic; attribute dont_touch of I35722: signal is true;
	signal I35723: std_logic; attribute dont_touch of I35723: signal is true;
	signal I35724: std_logic; attribute dont_touch of I35724: signal is true;
	signal I35729: std_logic; attribute dont_touch of I35729: signal is true;
	signal I35730: std_logic; attribute dont_touch of I35730: signal is true;
	signal I35731: std_logic; attribute dont_touch of I35731: signal is true;
	signal I35736: std_logic; attribute dont_touch of I35736: signal is true;
	signal I35737: std_logic; attribute dont_touch of I35737: signal is true;
	signal I35738: std_logic; attribute dont_touch of I35738: signal is true;
	signal I35743: std_logic; attribute dont_touch of I35743: signal is true;
	signal I35744: std_logic; attribute dont_touch of I35744: signal is true;
	signal I35745: std_logic; attribute dont_touch of I35745: signal is true;
	signal I35750: std_logic; attribute dont_touch of I35750: signal is true;
	signal I35751: std_logic; attribute dont_touch of I35751: signal is true;
	signal I35752: std_logic; attribute dont_touch of I35752: signal is true;
	signal WX35: std_logic; attribute dont_touch of WX35: signal is true;
	signal WX36: std_logic; attribute dont_touch of WX36: signal is true;
	signal WX37: std_logic; attribute dont_touch of WX37: signal is true;
	signal WX38: std_logic; attribute dont_touch of WX38: signal is true;
	signal WX39: std_logic; attribute dont_touch of WX39: signal is true;
	signal WX40: std_logic; attribute dont_touch of WX40: signal is true;
	signal WX41: std_logic; attribute dont_touch of WX41: signal is true;
	signal WX42: std_logic; attribute dont_touch of WX42: signal is true;
	signal WX43: std_logic; attribute dont_touch of WX43: signal is true;
	signal WX44: std_logic; attribute dont_touch of WX44: signal is true;
	signal WX45: std_logic; attribute dont_touch of WX45: signal is true;
	signal WX46: std_logic; attribute dont_touch of WX46: signal is true;
	signal WX47: std_logic; attribute dont_touch of WX47: signal is true;
	signal WX48: std_logic; attribute dont_touch of WX48: signal is true;
	signal WX49: std_logic; attribute dont_touch of WX49: signal is true;
	signal WX50: std_logic; attribute dont_touch of WX50: signal is true;
	signal WX51: std_logic; attribute dont_touch of WX51: signal is true;
	signal WX52: std_logic; attribute dont_touch of WX52: signal is true;
	signal WX53: std_logic; attribute dont_touch of WX53: signal is true;
	signal WX54: std_logic; attribute dont_touch of WX54: signal is true;
	signal WX55: std_logic; attribute dont_touch of WX55: signal is true;
	signal WX56: std_logic; attribute dont_touch of WX56: signal is true;
	signal WX57: std_logic; attribute dont_touch of WX57: signal is true;
	signal WX58: std_logic; attribute dont_touch of WX58: signal is true;
	signal WX59: std_logic; attribute dont_touch of WX59: signal is true;
	signal WX60: std_logic; attribute dont_touch of WX60: signal is true;
	signal WX61: std_logic; attribute dont_touch of WX61: signal is true;
	signal WX62: std_logic; attribute dont_touch of WX62: signal is true;
	signal WX63: std_logic; attribute dont_touch of WX63: signal is true;
	signal WX64: std_logic; attribute dont_touch of WX64: signal is true;
	signal WX65: std_logic; attribute dont_touch of WX65: signal is true;
	signal WX66: std_logic; attribute dont_touch of WX66: signal is true;
	signal WX67: std_logic; attribute dont_touch of WX67: signal is true;
	signal WX68: std_logic; attribute dont_touch of WX68: signal is true;
	signal WX69: std_logic; attribute dont_touch of WX69: signal is true;
	signal WX70: std_logic; attribute dont_touch of WX70: signal is true;
	signal WX71: std_logic; attribute dont_touch of WX71: signal is true;
	signal WX72: std_logic; attribute dont_touch of WX72: signal is true;
	signal WX73: std_logic; attribute dont_touch of WX73: signal is true;
	signal WX74: std_logic; attribute dont_touch of WX74: signal is true;
	signal WX75: std_logic; attribute dont_touch of WX75: signal is true;
	signal WX76: std_logic; attribute dont_touch of WX76: signal is true;
	signal WX77: std_logic; attribute dont_touch of WX77: signal is true;
	signal WX78: std_logic; attribute dont_touch of WX78: signal is true;
	signal WX79: std_logic; attribute dont_touch of WX79: signal is true;
	signal WX80: std_logic; attribute dont_touch of WX80: signal is true;
	signal WX81: std_logic; attribute dont_touch of WX81: signal is true;
	signal WX82: std_logic; attribute dont_touch of WX82: signal is true;
	signal WX83: std_logic; attribute dont_touch of WX83: signal is true;
	signal WX84: std_logic; attribute dont_touch of WX84: signal is true;
	signal WX85: std_logic; attribute dont_touch of WX85: signal is true;
	signal WX86: std_logic; attribute dont_touch of WX86: signal is true;
	signal WX87: std_logic; attribute dont_touch of WX87: signal is true;
	signal WX88: std_logic; attribute dont_touch of WX88: signal is true;
	signal WX89: std_logic; attribute dont_touch of WX89: signal is true;
	signal WX90: std_logic; attribute dont_touch of WX90: signal is true;
	signal WX91: std_logic; attribute dont_touch of WX91: signal is true;
	signal WX92: std_logic; attribute dont_touch of WX92: signal is true;
	signal WX93: std_logic; attribute dont_touch of WX93: signal is true;
	signal WX94: std_logic; attribute dont_touch of WX94: signal is true;
	signal WX95: std_logic; attribute dont_touch of WX95: signal is true;
	signal WX96: std_logic; attribute dont_touch of WX96: signal is true;
	signal WX97: std_logic; attribute dont_touch of WX97: signal is true;
	signal WX98: std_logic; attribute dont_touch of WX98: signal is true;
	signal WX99: std_logic; attribute dont_touch of WX99: signal is true;
	signal WX100: std_logic; attribute dont_touch of WX100: signal is true;
	signal WX101: std_logic; attribute dont_touch of WX101: signal is true;
	signal WX102: std_logic; attribute dont_touch of WX102: signal is true;
	signal WX103: std_logic; attribute dont_touch of WX103: signal is true;
	signal WX104: std_logic; attribute dont_touch of WX104: signal is true;
	signal WX105: std_logic; attribute dont_touch of WX105: signal is true;
	signal WX106: std_logic; attribute dont_touch of WX106: signal is true;
	signal WX107: std_logic; attribute dont_touch of WX107: signal is true;
	signal WX108: std_logic; attribute dont_touch of WX108: signal is true;
	signal WX109: std_logic; attribute dont_touch of WX109: signal is true;
	signal WX110: std_logic; attribute dont_touch of WX110: signal is true;
	signal WX111: std_logic; attribute dont_touch of WX111: signal is true;
	signal WX112: std_logic; attribute dont_touch of WX112: signal is true;
	signal WX113: std_logic; attribute dont_touch of WX113: signal is true;
	signal WX114: std_logic; attribute dont_touch of WX114: signal is true;
	signal WX115: std_logic; attribute dont_touch of WX115: signal is true;
	signal WX116: std_logic; attribute dont_touch of WX116: signal is true;
	signal WX117: std_logic; attribute dont_touch of WX117: signal is true;
	signal WX118: std_logic; attribute dont_touch of WX118: signal is true;
	signal WX119: std_logic; attribute dont_touch of WX119: signal is true;
	signal WX120: std_logic; attribute dont_touch of WX120: signal is true;
	signal WX121: std_logic; attribute dont_touch of WX121: signal is true;
	signal WX122: std_logic; attribute dont_touch of WX122: signal is true;
	signal WX123: std_logic; attribute dont_touch of WX123: signal is true;
	signal WX124: std_logic; attribute dont_touch of WX124: signal is true;
	signal WX125: std_logic; attribute dont_touch of WX125: signal is true;
	signal WX126: std_logic; attribute dont_touch of WX126: signal is true;
	signal WX127: std_logic; attribute dont_touch of WX127: signal is true;
	signal WX128: std_logic; attribute dont_touch of WX128: signal is true;
	signal WX129: std_logic; attribute dont_touch of WX129: signal is true;
	signal WX130: std_logic; attribute dont_touch of WX130: signal is true;
	signal WX131: std_logic; attribute dont_touch of WX131: signal is true;
	signal WX132: std_logic; attribute dont_touch of WX132: signal is true;
	signal WX133: std_logic; attribute dont_touch of WX133: signal is true;
	signal WX134: std_logic; attribute dont_touch of WX134: signal is true;
	signal WX135: std_logic; attribute dont_touch of WX135: signal is true;
	signal WX136: std_logic; attribute dont_touch of WX136: signal is true;
	signal WX137: std_logic; attribute dont_touch of WX137: signal is true;
	signal WX138: std_logic; attribute dont_touch of WX138: signal is true;
	signal WX139: std_logic; attribute dont_touch of WX139: signal is true;
	signal WX140: std_logic; attribute dont_touch of WX140: signal is true;
	signal WX141: std_logic; attribute dont_touch of WX141: signal is true;
	signal WX142: std_logic; attribute dont_touch of WX142: signal is true;
	signal WX143: std_logic; attribute dont_touch of WX143: signal is true;
	signal WX144: std_logic; attribute dont_touch of WX144: signal is true;
	signal WX145: std_logic; attribute dont_touch of WX145: signal is true;
	signal WX146: std_logic; attribute dont_touch of WX146: signal is true;
	signal WX147: std_logic; attribute dont_touch of WX147: signal is true;
	signal WX148: std_logic; attribute dont_touch of WX148: signal is true;
	signal WX149: std_logic; attribute dont_touch of WX149: signal is true;
	signal WX150: std_logic; attribute dont_touch of WX150: signal is true;
	signal WX151: std_logic; attribute dont_touch of WX151: signal is true;
	signal WX152: std_logic; attribute dont_touch of WX152: signal is true;
	signal WX153: std_logic; attribute dont_touch of WX153: signal is true;
	signal WX154: std_logic; attribute dont_touch of WX154: signal is true;
	signal WX155: std_logic; attribute dont_touch of WX155: signal is true;
	signal WX156: std_logic; attribute dont_touch of WX156: signal is true;
	signal WX157: std_logic; attribute dont_touch of WX157: signal is true;
	signal WX158: std_logic; attribute dont_touch of WX158: signal is true;
	signal WX159: std_logic; attribute dont_touch of WX159: signal is true;
	signal WX160: std_logic; attribute dont_touch of WX160: signal is true;
	signal WX161: std_logic; attribute dont_touch of WX161: signal is true;
	signal WX162: std_logic; attribute dont_touch of WX162: signal is true;
	signal WX163: std_logic; attribute dont_touch of WX163: signal is true;
	signal WX164: std_logic; attribute dont_touch of WX164: signal is true;
	signal WX165: std_logic; attribute dont_touch of WX165: signal is true;
	signal WX166: std_logic; attribute dont_touch of WX166: signal is true;
	signal WX167: std_logic; attribute dont_touch of WX167: signal is true;
	signal WX168: std_logic; attribute dont_touch of WX168: signal is true;
	signal WX169: std_logic; attribute dont_touch of WX169: signal is true;
	signal WX170: std_logic; attribute dont_touch of WX170: signal is true;
	signal WX171: std_logic; attribute dont_touch of WX171: signal is true;
	signal WX172: std_logic; attribute dont_touch of WX172: signal is true;
	signal WX173: std_logic; attribute dont_touch of WX173: signal is true;
	signal WX174: std_logic; attribute dont_touch of WX174: signal is true;
	signal WX175: std_logic; attribute dont_touch of WX175: signal is true;
	signal WX176: std_logic; attribute dont_touch of WX176: signal is true;
	signal WX177: std_logic; attribute dont_touch of WX177: signal is true;
	signal WX178: std_logic; attribute dont_touch of WX178: signal is true;
	signal WX179: std_logic; attribute dont_touch of WX179: signal is true;
	signal WX180: std_logic; attribute dont_touch of WX180: signal is true;
	signal WX181: std_logic; attribute dont_touch of WX181: signal is true;
	signal WX182: std_logic; attribute dont_touch of WX182: signal is true;
	signal WX183: std_logic; attribute dont_touch of WX183: signal is true;
	signal WX184: std_logic; attribute dont_touch of WX184: signal is true;
	signal WX185: std_logic; attribute dont_touch of WX185: signal is true;
	signal WX186: std_logic; attribute dont_touch of WX186: signal is true;
	signal WX187: std_logic; attribute dont_touch of WX187: signal is true;
	signal WX188: std_logic; attribute dont_touch of WX188: signal is true;
	signal WX189: std_logic; attribute dont_touch of WX189: signal is true;
	signal WX190: std_logic; attribute dont_touch of WX190: signal is true;
	signal WX191: std_logic; attribute dont_touch of WX191: signal is true;
	signal WX192: std_logic; attribute dont_touch of WX192: signal is true;
	signal WX193: std_logic; attribute dont_touch of WX193: signal is true;
	signal WX194: std_logic; attribute dont_touch of WX194: signal is true;
	signal WX195: std_logic; attribute dont_touch of WX195: signal is true;
	signal WX196: std_logic; attribute dont_touch of WX196: signal is true;
	signal WX197: std_logic; attribute dont_touch of WX197: signal is true;
	signal WX198: std_logic; attribute dont_touch of WX198: signal is true;
	signal WX199: std_logic; attribute dont_touch of WX199: signal is true;
	signal WX200: std_logic; attribute dont_touch of WX200: signal is true;
	signal WX201: std_logic; attribute dont_touch of WX201: signal is true;
	signal WX202: std_logic; attribute dont_touch of WX202: signal is true;
	signal WX203: std_logic; attribute dont_touch of WX203: signal is true;
	signal WX204: std_logic; attribute dont_touch of WX204: signal is true;
	signal WX205: std_logic; attribute dont_touch of WX205: signal is true;
	signal WX206: std_logic; attribute dont_touch of WX206: signal is true;
	signal WX207: std_logic; attribute dont_touch of WX207: signal is true;
	signal WX208: std_logic; attribute dont_touch of WX208: signal is true;
	signal WX209: std_logic; attribute dont_touch of WX209: signal is true;
	signal WX210: std_logic; attribute dont_touch of WX210: signal is true;
	signal WX211: std_logic; attribute dont_touch of WX211: signal is true;
	signal WX212: std_logic; attribute dont_touch of WX212: signal is true;
	signal WX213: std_logic; attribute dont_touch of WX213: signal is true;
	signal WX214: std_logic; attribute dont_touch of WX214: signal is true;
	signal WX215: std_logic; attribute dont_touch of WX215: signal is true;
	signal WX216: std_logic; attribute dont_touch of WX216: signal is true;
	signal WX217: std_logic; attribute dont_touch of WX217: signal is true;
	signal WX218: std_logic; attribute dont_touch of WX218: signal is true;
	signal WX219: std_logic; attribute dont_touch of WX219: signal is true;
	signal WX220: std_logic; attribute dont_touch of WX220: signal is true;
	signal WX221: std_logic; attribute dont_touch of WX221: signal is true;
	signal WX222: std_logic; attribute dont_touch of WX222: signal is true;
	signal WX223: std_logic; attribute dont_touch of WX223: signal is true;
	signal WX224: std_logic; attribute dont_touch of WX224: signal is true;
	signal WX225: std_logic; attribute dont_touch of WX225: signal is true;
	signal WX226: std_logic; attribute dont_touch of WX226: signal is true;
	signal WX227: std_logic; attribute dont_touch of WX227: signal is true;
	signal WX228: std_logic; attribute dont_touch of WX228: signal is true;
	signal WX229: std_logic; attribute dont_touch of WX229: signal is true;
	signal WX230: std_logic; attribute dont_touch of WX230: signal is true;
	signal WX231: std_logic; attribute dont_touch of WX231: signal is true;
	signal WX232: std_logic; attribute dont_touch of WX232: signal is true;
	signal WX233: std_logic; attribute dont_touch of WX233: signal is true;
	signal WX234: std_logic; attribute dont_touch of WX234: signal is true;
	signal WX235: std_logic; attribute dont_touch of WX235: signal is true;
	signal WX236: std_logic; attribute dont_touch of WX236: signal is true;
	signal WX237: std_logic; attribute dont_touch of WX237: signal is true;
	signal WX238: std_logic; attribute dont_touch of WX238: signal is true;
	signal WX239: std_logic; attribute dont_touch of WX239: signal is true;
	signal WX240: std_logic; attribute dont_touch of WX240: signal is true;
	signal WX241: std_logic; attribute dont_touch of WX241: signal is true;
	signal WX242: std_logic; attribute dont_touch of WX242: signal is true;
	signal WX243: std_logic; attribute dont_touch of WX243: signal is true;
	signal WX244: std_logic; attribute dont_touch of WX244: signal is true;
	signal WX245: std_logic; attribute dont_touch of WX245: signal is true;
	signal WX246: std_logic; attribute dont_touch of WX246: signal is true;
	signal WX247: std_logic; attribute dont_touch of WX247: signal is true;
	signal WX248: std_logic; attribute dont_touch of WX248: signal is true;
	signal WX249: std_logic; attribute dont_touch of WX249: signal is true;
	signal WX250: std_logic; attribute dont_touch of WX250: signal is true;
	signal WX251: std_logic; attribute dont_touch of WX251: signal is true;
	signal WX252: std_logic; attribute dont_touch of WX252: signal is true;
	signal WX253: std_logic; attribute dont_touch of WX253: signal is true;
	signal WX254: std_logic; attribute dont_touch of WX254: signal is true;
	signal WX255: std_logic; attribute dont_touch of WX255: signal is true;
	signal WX256: std_logic; attribute dont_touch of WX256: signal is true;
	signal WX257: std_logic; attribute dont_touch of WX257: signal is true;
	signal WX258: std_logic; attribute dont_touch of WX258: signal is true;
	signal WX259: std_logic; attribute dont_touch of WX259: signal is true;
	signal WX260: std_logic; attribute dont_touch of WX260: signal is true;
	signal WX261: std_logic; attribute dont_touch of WX261: signal is true;
	signal WX262: std_logic; attribute dont_touch of WX262: signal is true;
	signal WX263: std_logic; attribute dont_touch of WX263: signal is true;
	signal WX264: std_logic; attribute dont_touch of WX264: signal is true;
	signal WX265: std_logic; attribute dont_touch of WX265: signal is true;
	signal WX266: std_logic; attribute dont_touch of WX266: signal is true;
	signal WX267: std_logic; attribute dont_touch of WX267: signal is true;
	signal WX268: std_logic; attribute dont_touch of WX268: signal is true;
	signal WX269: std_logic; attribute dont_touch of WX269: signal is true;
	signal WX270: std_logic; attribute dont_touch of WX270: signal is true;
	signal WX271: std_logic; attribute dont_touch of WX271: signal is true;
	signal WX272: std_logic; attribute dont_touch of WX272: signal is true;
	signal WX273: std_logic; attribute dont_touch of WX273: signal is true;
	signal WX274: std_logic; attribute dont_touch of WX274: signal is true;
	signal WX275: std_logic; attribute dont_touch of WX275: signal is true;
	signal WX276: std_logic; attribute dont_touch of WX276: signal is true;
	signal WX277: std_logic; attribute dont_touch of WX277: signal is true;
	signal WX278: std_logic; attribute dont_touch of WX278: signal is true;
	signal WX279: std_logic; attribute dont_touch of WX279: signal is true;
	signal WX280: std_logic; attribute dont_touch of WX280: signal is true;
	signal WX281: std_logic; attribute dont_touch of WX281: signal is true;
	signal WX282: std_logic; attribute dont_touch of WX282: signal is true;
	signal WX283: std_logic; attribute dont_touch of WX283: signal is true;
	signal WX284: std_logic; attribute dont_touch of WX284: signal is true;
	signal WX285: std_logic; attribute dont_touch of WX285: signal is true;
	signal WX286: std_logic; attribute dont_touch of WX286: signal is true;
	signal WX287: std_logic; attribute dont_touch of WX287: signal is true;
	signal WX288: std_logic; attribute dont_touch of WX288: signal is true;
	signal WX289: std_logic; attribute dont_touch of WX289: signal is true;
	signal WX290: std_logic; attribute dont_touch of WX290: signal is true;
	signal WX291: std_logic; attribute dont_touch of WX291: signal is true;
	signal WX292: std_logic; attribute dont_touch of WX292: signal is true;
	signal WX293: std_logic; attribute dont_touch of WX293: signal is true;
	signal WX294: std_logic; attribute dont_touch of WX294: signal is true;
	signal WX295: std_logic; attribute dont_touch of WX295: signal is true;
	signal WX296: std_logic; attribute dont_touch of WX296: signal is true;
	signal WX297: std_logic; attribute dont_touch of WX297: signal is true;
	signal WX298: std_logic; attribute dont_touch of WX298: signal is true;
	signal WX299: std_logic; attribute dont_touch of WX299: signal is true;
	signal WX300: std_logic; attribute dont_touch of WX300: signal is true;
	signal WX301: std_logic; attribute dont_touch of WX301: signal is true;
	signal WX302: std_logic; attribute dont_touch of WX302: signal is true;
	signal WX303: std_logic; attribute dont_touch of WX303: signal is true;
	signal WX304: std_logic; attribute dont_touch of WX304: signal is true;
	signal WX305: std_logic; attribute dont_touch of WX305: signal is true;
	signal WX306: std_logic; attribute dont_touch of WX306: signal is true;
	signal WX307: std_logic; attribute dont_touch of WX307: signal is true;
	signal WX308: std_logic; attribute dont_touch of WX308: signal is true;
	signal WX309: std_logic; attribute dont_touch of WX309: signal is true;
	signal WX310: std_logic; attribute dont_touch of WX310: signal is true;
	signal WX311: std_logic; attribute dont_touch of WX311: signal is true;
	signal WX312: std_logic; attribute dont_touch of WX312: signal is true;
	signal WX313: std_logic; attribute dont_touch of WX313: signal is true;
	signal WX314: std_logic; attribute dont_touch of WX314: signal is true;
	signal WX315: std_logic; attribute dont_touch of WX315: signal is true;
	signal WX316: std_logic; attribute dont_touch of WX316: signal is true;
	signal WX317: std_logic; attribute dont_touch of WX317: signal is true;
	signal WX318: std_logic; attribute dont_touch of WX318: signal is true;
	signal WX319: std_logic; attribute dont_touch of WX319: signal is true;
	signal WX320: std_logic; attribute dont_touch of WX320: signal is true;
	signal WX321: std_logic; attribute dont_touch of WX321: signal is true;
	signal WX322: std_logic; attribute dont_touch of WX322: signal is true;
	signal WX323: std_logic; attribute dont_touch of WX323: signal is true;
	signal WX324: std_logic; attribute dont_touch of WX324: signal is true;
	signal WX325: std_logic; attribute dont_touch of WX325: signal is true;
	signal WX326: std_logic; attribute dont_touch of WX326: signal is true;
	signal WX327: std_logic; attribute dont_touch of WX327: signal is true;
	signal WX328: std_logic; attribute dont_touch of WX328: signal is true;
	signal WX329: std_logic; attribute dont_touch of WX329: signal is true;
	signal WX330: std_logic; attribute dont_touch of WX330: signal is true;
	signal WX331: std_logic; attribute dont_touch of WX331: signal is true;
	signal WX332: std_logic; attribute dont_touch of WX332: signal is true;
	signal WX333: std_logic; attribute dont_touch of WX333: signal is true;
	signal WX334: std_logic; attribute dont_touch of WX334: signal is true;
	signal WX335: std_logic; attribute dont_touch of WX335: signal is true;
	signal WX336: std_logic; attribute dont_touch of WX336: signal is true;
	signal WX337: std_logic; attribute dont_touch of WX337: signal is true;
	signal WX338: std_logic; attribute dont_touch of WX338: signal is true;
	signal WX339: std_logic; attribute dont_touch of WX339: signal is true;
	signal WX340: std_logic; attribute dont_touch of WX340: signal is true;
	signal WX341: std_logic; attribute dont_touch of WX341: signal is true;
	signal WX342: std_logic; attribute dont_touch of WX342: signal is true;
	signal WX343: std_logic; attribute dont_touch of WX343: signal is true;
	signal WX344: std_logic; attribute dont_touch of WX344: signal is true;
	signal WX345: std_logic; attribute dont_touch of WX345: signal is true;
	signal WX346: std_logic; attribute dont_touch of WX346: signal is true;
	signal WX347: std_logic; attribute dont_touch of WX347: signal is true;
	signal WX348: std_logic; attribute dont_touch of WX348: signal is true;
	signal WX349: std_logic; attribute dont_touch of WX349: signal is true;
	signal WX350: std_logic; attribute dont_touch of WX350: signal is true;
	signal WX351: std_logic; attribute dont_touch of WX351: signal is true;
	signal WX352: std_logic; attribute dont_touch of WX352: signal is true;
	signal WX353: std_logic; attribute dont_touch of WX353: signal is true;
	signal WX354: std_logic; attribute dont_touch of WX354: signal is true;
	signal WX355: std_logic; attribute dont_touch of WX355: signal is true;
	signal WX356: std_logic; attribute dont_touch of WX356: signal is true;
	signal WX357: std_logic; attribute dont_touch of WX357: signal is true;
	signal WX358: std_logic; attribute dont_touch of WX358: signal is true;
	signal WX359: std_logic; attribute dont_touch of WX359: signal is true;
	signal WX360: std_logic; attribute dont_touch of WX360: signal is true;
	signal WX361: std_logic; attribute dont_touch of WX361: signal is true;
	signal WX362: std_logic; attribute dont_touch of WX362: signal is true;
	signal WX363: std_logic; attribute dont_touch of WX363: signal is true;
	signal WX364: std_logic; attribute dont_touch of WX364: signal is true;
	signal WX365: std_logic; attribute dont_touch of WX365: signal is true;
	signal WX366: std_logic; attribute dont_touch of WX366: signal is true;
	signal WX367: std_logic; attribute dont_touch of WX367: signal is true;
	signal WX368: std_logic; attribute dont_touch of WX368: signal is true;
	signal WX369: std_logic; attribute dont_touch of WX369: signal is true;
	signal WX370: std_logic; attribute dont_touch of WX370: signal is true;
	signal WX371: std_logic; attribute dont_touch of WX371: signal is true;
	signal WX372: std_logic; attribute dont_touch of WX372: signal is true;
	signal WX373: std_logic; attribute dont_touch of WX373: signal is true;
	signal WX374: std_logic; attribute dont_touch of WX374: signal is true;
	signal WX375: std_logic; attribute dont_touch of WX375: signal is true;
	signal WX376: std_logic; attribute dont_touch of WX376: signal is true;
	signal WX377: std_logic; attribute dont_touch of WX377: signal is true;
	signal WX378: std_logic; attribute dont_touch of WX378: signal is true;
	signal WX379: std_logic; attribute dont_touch of WX379: signal is true;
	signal WX380: std_logic; attribute dont_touch of WX380: signal is true;
	signal WX381: std_logic; attribute dont_touch of WX381: signal is true;
	signal WX382: std_logic; attribute dont_touch of WX382: signal is true;
	signal WX383: std_logic; attribute dont_touch of WX383: signal is true;
	signal WX384: std_logic; attribute dont_touch of WX384: signal is true;
	signal WX385: std_logic; attribute dont_touch of WX385: signal is true;
	signal WX386: std_logic; attribute dont_touch of WX386: signal is true;
	signal WX387: std_logic; attribute dont_touch of WX387: signal is true;
	signal WX388: std_logic; attribute dont_touch of WX388: signal is true;
	signal WX389: std_logic; attribute dont_touch of WX389: signal is true;
	signal WX390: std_logic; attribute dont_touch of WX390: signal is true;
	signal WX391: std_logic; attribute dont_touch of WX391: signal is true;
	signal WX392: std_logic; attribute dont_touch of WX392: signal is true;
	signal WX393: std_logic; attribute dont_touch of WX393: signal is true;
	signal WX394: std_logic; attribute dont_touch of WX394: signal is true;
	signal WX395: std_logic; attribute dont_touch of WX395: signal is true;
	signal WX396: std_logic; attribute dont_touch of WX396: signal is true;
	signal WX397: std_logic; attribute dont_touch of WX397: signal is true;
	signal WX398: std_logic; attribute dont_touch of WX398: signal is true;
	signal WX399: std_logic; attribute dont_touch of WX399: signal is true;
	signal WX400: std_logic; attribute dont_touch of WX400: signal is true;
	signal WX401: std_logic; attribute dont_touch of WX401: signal is true;
	signal WX402: std_logic; attribute dont_touch of WX402: signal is true;
	signal WX403: std_logic; attribute dont_touch of WX403: signal is true;
	signal WX404: std_logic; attribute dont_touch of WX404: signal is true;
	signal WX405: std_logic; attribute dont_touch of WX405: signal is true;
	signal WX406: std_logic; attribute dont_touch of WX406: signal is true;
	signal WX407: std_logic; attribute dont_touch of WX407: signal is true;
	signal WX408: std_logic; attribute dont_touch of WX408: signal is true;
	signal WX409: std_logic; attribute dont_touch of WX409: signal is true;
	signal WX410: std_logic; attribute dont_touch of WX410: signal is true;
	signal WX411: std_logic; attribute dont_touch of WX411: signal is true;
	signal WX412: std_logic; attribute dont_touch of WX412: signal is true;
	signal WX413: std_logic; attribute dont_touch of WX413: signal is true;
	signal WX414: std_logic; attribute dont_touch of WX414: signal is true;
	signal WX415: std_logic; attribute dont_touch of WX415: signal is true;
	signal WX416: std_logic; attribute dont_touch of WX416: signal is true;
	signal WX417: std_logic; attribute dont_touch of WX417: signal is true;
	signal WX418: std_logic; attribute dont_touch of WX418: signal is true;
	signal WX419: std_logic; attribute dont_touch of WX419: signal is true;
	signal WX420: std_logic; attribute dont_touch of WX420: signal is true;
	signal WX421: std_logic; attribute dont_touch of WX421: signal is true;
	signal WX422: std_logic; attribute dont_touch of WX422: signal is true;
	signal WX423: std_logic; attribute dont_touch of WX423: signal is true;
	signal WX424: std_logic; attribute dont_touch of WX424: signal is true;
	signal WX425: std_logic; attribute dont_touch of WX425: signal is true;
	signal WX426: std_logic; attribute dont_touch of WX426: signal is true;
	signal WX427: std_logic; attribute dont_touch of WX427: signal is true;
	signal WX428: std_logic; attribute dont_touch of WX428: signal is true;
	signal WX429: std_logic; attribute dont_touch of WX429: signal is true;
	signal WX430: std_logic; attribute dont_touch of WX430: signal is true;
	signal WX431: std_logic; attribute dont_touch of WX431: signal is true;
	signal WX432: std_logic; attribute dont_touch of WX432: signal is true;
	signal WX433: std_logic; attribute dont_touch of WX433: signal is true;
	signal WX434: std_logic; attribute dont_touch of WX434: signal is true;
	signal WX435: std_logic; attribute dont_touch of WX435: signal is true;
	signal WX436: std_logic; attribute dont_touch of WX436: signal is true;
	signal WX437: std_logic; attribute dont_touch of WX437: signal is true;
	signal WX438: std_logic; attribute dont_touch of WX438: signal is true;
	signal WX439: std_logic; attribute dont_touch of WX439: signal is true;
	signal WX440: std_logic; attribute dont_touch of WX440: signal is true;
	signal WX441: std_logic; attribute dont_touch of WX441: signal is true;
	signal WX442: std_logic; attribute dont_touch of WX442: signal is true;
	signal WX443: std_logic; attribute dont_touch of WX443: signal is true;
	signal WX444: std_logic; attribute dont_touch of WX444: signal is true;
	signal WX445: std_logic; attribute dont_touch of WX445: signal is true;
	signal WX446: std_logic; attribute dont_touch of WX446: signal is true;
	signal WX447: std_logic; attribute dont_touch of WX447: signal is true;
	signal WX448: std_logic; attribute dont_touch of WX448: signal is true;
	signal WX449: std_logic; attribute dont_touch of WX449: signal is true;
	signal WX450: std_logic; attribute dont_touch of WX450: signal is true;
	signal WX451: std_logic; attribute dont_touch of WX451: signal is true;
	signal WX452: std_logic; attribute dont_touch of WX452: signal is true;
	signal WX453: std_logic; attribute dont_touch of WX453: signal is true;
	signal WX454: std_logic; attribute dont_touch of WX454: signal is true;
	signal WX455: std_logic; attribute dont_touch of WX455: signal is true;
	signal WX456: std_logic; attribute dont_touch of WX456: signal is true;
	signal WX457: std_logic; attribute dont_touch of WX457: signal is true;
	signal WX458: std_logic; attribute dont_touch of WX458: signal is true;
	signal WX459: std_logic; attribute dont_touch of WX459: signal is true;
	signal WX460: std_logic; attribute dont_touch of WX460: signal is true;
	signal WX461: std_logic; attribute dont_touch of WX461: signal is true;
	signal WX462: std_logic; attribute dont_touch of WX462: signal is true;
	signal WX463: std_logic; attribute dont_touch of WX463: signal is true;
	signal WX464: std_logic; attribute dont_touch of WX464: signal is true;
	signal WX465: std_logic; attribute dont_touch of WX465: signal is true;
	signal WX466: std_logic; attribute dont_touch of WX466: signal is true;
	signal WX467: std_logic; attribute dont_touch of WX467: signal is true;
	signal WX468: std_logic; attribute dont_touch of WX468: signal is true;
	signal WX469: std_logic; attribute dont_touch of WX469: signal is true;
	signal WX470: std_logic; attribute dont_touch of WX470: signal is true;
	signal WX471: std_logic; attribute dont_touch of WX471: signal is true;
	signal WX472: std_logic; attribute dont_touch of WX472: signal is true;
	signal WX473: std_logic; attribute dont_touch of WX473: signal is true;
	signal WX474: std_logic; attribute dont_touch of WX474: signal is true;
	signal WX475: std_logic; attribute dont_touch of WX475: signal is true;
	signal WX476: std_logic; attribute dont_touch of WX476: signal is true;
	signal WX477: std_logic; attribute dont_touch of WX477: signal is true;
	signal WX478: std_logic; attribute dont_touch of WX478: signal is true;
	signal WX479: std_logic; attribute dont_touch of WX479: signal is true;
	signal WX480: std_logic; attribute dont_touch of WX480: signal is true;
	signal WX481: std_logic; attribute dont_touch of WX481: signal is true;
	signal WX482: std_logic; attribute dont_touch of WX482: signal is true;
	signal WX483: std_logic; attribute dont_touch of WX483: signal is true;
	signal WX484: std_logic; attribute dont_touch of WX484: signal is true;
	signal WX485: std_logic; attribute dont_touch of WX485: signal is true;
	signal WX486: std_logic; attribute dont_touch of WX486: signal is true;
	signal WX487: std_logic; attribute dont_touch of WX487: signal is true;
	signal WX488: std_logic; attribute dont_touch of WX488: signal is true;
	signal WX489: std_logic; attribute dont_touch of WX489: signal is true;
	signal WX490: std_logic; attribute dont_touch of WX490: signal is true;
	signal WX491: std_logic; attribute dont_touch of WX491: signal is true;
	signal WX492: std_logic; attribute dont_touch of WX492: signal is true;
	signal WX493: std_logic; attribute dont_touch of WX493: signal is true;
	signal WX494: std_logic; attribute dont_touch of WX494: signal is true;
	signal WX495: std_logic; attribute dont_touch of WX495: signal is true;
	signal WX496: std_logic; attribute dont_touch of WX496: signal is true;
	signal WX497: std_logic; attribute dont_touch of WX497: signal is true;
	signal WX498: std_logic; attribute dont_touch of WX498: signal is true;
	signal WX499: std_logic; attribute dont_touch of WX499: signal is true;
	signal WX500: std_logic; attribute dont_touch of WX500: signal is true;
	signal WX501: std_logic; attribute dont_touch of WX501: signal is true;
	signal WX502: std_logic; attribute dont_touch of WX502: signal is true;
	signal WX503: std_logic; attribute dont_touch of WX503: signal is true;
	signal WX504: std_logic; attribute dont_touch of WX504: signal is true;
	signal WX505: std_logic; attribute dont_touch of WX505: signal is true;
	signal WX506: std_logic; attribute dont_touch of WX506: signal is true;
	signal WX507: std_logic; attribute dont_touch of WX507: signal is true;
	signal WX508: std_logic; attribute dont_touch of WX508: signal is true;
	signal WX509: std_logic; attribute dont_touch of WX509: signal is true;
	signal WX510: std_logic; attribute dont_touch of WX510: signal is true;
	signal WX511: std_logic; attribute dont_touch of WX511: signal is true;
	signal WX512: std_logic; attribute dont_touch of WX512: signal is true;
	signal WX513: std_logic; attribute dont_touch of WX513: signal is true;
	signal WX514: std_logic; attribute dont_touch of WX514: signal is true;
	signal WX515: std_logic; attribute dont_touch of WX515: signal is true;
	signal WX516: std_logic; attribute dont_touch of WX516: signal is true;
	signal WX517: std_logic; attribute dont_touch of WX517: signal is true;
	signal WX518: std_logic; attribute dont_touch of WX518: signal is true;
	signal WX519: std_logic; attribute dont_touch of WX519: signal is true;
	signal WX520: std_logic; attribute dont_touch of WX520: signal is true;
	signal WX521: std_logic; attribute dont_touch of WX521: signal is true;
	signal WX522: std_logic; attribute dont_touch of WX522: signal is true;
	signal WX523: std_logic; attribute dont_touch of WX523: signal is true;
	signal WX524: std_logic; attribute dont_touch of WX524: signal is true;
	signal WX525: std_logic; attribute dont_touch of WX525: signal is true;
	signal WX526: std_logic; attribute dont_touch of WX526: signal is true;
	signal WX527: std_logic; attribute dont_touch of WX527: signal is true;
	signal WX528: std_logic; attribute dont_touch of WX528: signal is true;
	signal WX529: std_logic; attribute dont_touch of WX529: signal is true;
	signal WX530: std_logic; attribute dont_touch of WX530: signal is true;
	signal WX531: std_logic; attribute dont_touch of WX531: signal is true;
	signal WX532: std_logic; attribute dont_touch of WX532: signal is true;
	signal WX533: std_logic; attribute dont_touch of WX533: signal is true;
	signal WX534: std_logic; attribute dont_touch of WX534: signal is true;
	signal WX535: std_logic; attribute dont_touch of WX535: signal is true;
	signal WX536: std_logic; attribute dont_touch of WX536: signal is true;
	signal WX537: std_logic; attribute dont_touch of WX537: signal is true;
	signal WX538: std_logic; attribute dont_touch of WX538: signal is true;
	signal WX539: std_logic; attribute dont_touch of WX539: signal is true;
	signal WX540: std_logic; attribute dont_touch of WX540: signal is true;
	signal WX541: std_logic; attribute dont_touch of WX541: signal is true;
	signal WX542: std_logic; attribute dont_touch of WX542: signal is true;
	signal WX543: std_logic; attribute dont_touch of WX543: signal is true;
	signal WX544: std_logic; attribute dont_touch of WX544: signal is true;
	signal WX545: std_logic; attribute dont_touch of WX545: signal is true;
	signal WX546: std_logic; attribute dont_touch of WX546: signal is true;
	signal WX547: std_logic; attribute dont_touch of WX547: signal is true;
	signal WX548: std_logic; attribute dont_touch of WX548: signal is true;
	signal WX549: std_logic; attribute dont_touch of WX549: signal is true;
	signal WX550: std_logic; attribute dont_touch of WX550: signal is true;
	signal WX551: std_logic; attribute dont_touch of WX551: signal is true;
	signal WX552: std_logic; attribute dont_touch of WX552: signal is true;
	signal WX553: std_logic; attribute dont_touch of WX553: signal is true;
	signal WX554: std_logic; attribute dont_touch of WX554: signal is true;
	signal WX555: std_logic; attribute dont_touch of WX555: signal is true;
	signal WX556: std_logic; attribute dont_touch of WX556: signal is true;
	signal WX557: std_logic; attribute dont_touch of WX557: signal is true;
	signal WX558: std_logic; attribute dont_touch of WX558: signal is true;
	signal WX559: std_logic; attribute dont_touch of WX559: signal is true;
	signal WX560: std_logic; attribute dont_touch of WX560: signal is true;
	signal WX561: std_logic; attribute dont_touch of WX561: signal is true;
	signal WX562: std_logic; attribute dont_touch of WX562: signal is true;
	signal WX563: std_logic; attribute dont_touch of WX563: signal is true;
	signal WX564: std_logic; attribute dont_touch of WX564: signal is true;
	signal WX565: std_logic; attribute dont_touch of WX565: signal is true;
	signal WX566: std_logic; attribute dont_touch of WX566: signal is true;
	signal WX567: std_logic; attribute dont_touch of WX567: signal is true;
	signal WX568: std_logic; attribute dont_touch of WX568: signal is true;
	signal WX569: std_logic; attribute dont_touch of WX569: signal is true;
	signal WX570: std_logic; attribute dont_touch of WX570: signal is true;
	signal WX571: std_logic; attribute dont_touch of WX571: signal is true;
	signal WX572: std_logic; attribute dont_touch of WX572: signal is true;
	signal WX573: std_logic; attribute dont_touch of WX573: signal is true;
	signal WX574: std_logic; attribute dont_touch of WX574: signal is true;
	signal WX575: std_logic; attribute dont_touch of WX575: signal is true;
	signal WX576: std_logic; attribute dont_touch of WX576: signal is true;
	signal WX577: std_logic; attribute dont_touch of WX577: signal is true;
	signal WX578: std_logic; attribute dont_touch of WX578: signal is true;
	signal WX579: std_logic; attribute dont_touch of WX579: signal is true;
	signal WX580: std_logic; attribute dont_touch of WX580: signal is true;
	signal WX581: std_logic; attribute dont_touch of WX581: signal is true;
	signal WX582: std_logic; attribute dont_touch of WX582: signal is true;
	signal WX583: std_logic; attribute dont_touch of WX583: signal is true;
	signal WX584: std_logic; attribute dont_touch of WX584: signal is true;
	signal WX585: std_logic; attribute dont_touch of WX585: signal is true;
	signal WX586: std_logic; attribute dont_touch of WX586: signal is true;
	signal WX587: std_logic; attribute dont_touch of WX587: signal is true;
	signal WX588: std_logic; attribute dont_touch of WX588: signal is true;
	signal WX589: std_logic; attribute dont_touch of WX589: signal is true;
	signal WX590: std_logic; attribute dont_touch of WX590: signal is true;
	signal WX591: std_logic; attribute dont_touch of WX591: signal is true;
	signal WX592: std_logic; attribute dont_touch of WX592: signal is true;
	signal WX593: std_logic; attribute dont_touch of WX593: signal is true;
	signal WX594: std_logic; attribute dont_touch of WX594: signal is true;
	signal WX595: std_logic; attribute dont_touch of WX595: signal is true;
	signal WX596: std_logic; attribute dont_touch of WX596: signal is true;
	signal WX597: std_logic; attribute dont_touch of WX597: signal is true;
	signal WX598: std_logic; attribute dont_touch of WX598: signal is true;
	signal WX599: std_logic; attribute dont_touch of WX599: signal is true;
	signal WX600: std_logic; attribute dont_touch of WX600: signal is true;
	signal WX601: std_logic; attribute dont_touch of WX601: signal is true;
	signal WX602: std_logic; attribute dont_touch of WX602: signal is true;
	signal WX603: std_logic; attribute dont_touch of WX603: signal is true;
	signal WX604: std_logic; attribute dont_touch of WX604: signal is true;
	signal WX605: std_logic; attribute dont_touch of WX605: signal is true;
	signal WX606: std_logic; attribute dont_touch of WX606: signal is true;
	signal WX607: std_logic; attribute dont_touch of WX607: signal is true;
	signal WX608: std_logic; attribute dont_touch of WX608: signal is true;
	signal WX609: std_logic; attribute dont_touch of WX609: signal is true;
	signal WX610: std_logic; attribute dont_touch of WX610: signal is true;
	signal WX611: std_logic; attribute dont_touch of WX611: signal is true;
	signal WX612: std_logic; attribute dont_touch of WX612: signal is true;
	signal WX613: std_logic; attribute dont_touch of WX613: signal is true;
	signal WX614: std_logic; attribute dont_touch of WX614: signal is true;
	signal WX615: std_logic; attribute dont_touch of WX615: signal is true;
	signal WX616: std_logic; attribute dont_touch of WX616: signal is true;
	signal WX617: std_logic; attribute dont_touch of WX617: signal is true;
	signal WX618: std_logic; attribute dont_touch of WX618: signal is true;
	signal WX619: std_logic; attribute dont_touch of WX619: signal is true;
	signal WX620: std_logic; attribute dont_touch of WX620: signal is true;
	signal WX621: std_logic; attribute dont_touch of WX621: signal is true;
	signal WX622: std_logic; attribute dont_touch of WX622: signal is true;
	signal WX623: std_logic; attribute dont_touch of WX623: signal is true;
	signal WX624: std_logic; attribute dont_touch of WX624: signal is true;
	signal WX625: std_logic; attribute dont_touch of WX625: signal is true;
	signal WX626: std_logic; attribute dont_touch of WX626: signal is true;
	signal WX627: std_logic; attribute dont_touch of WX627: signal is true;
	signal WX628: std_logic; attribute dont_touch of WX628: signal is true;
	signal WX629: std_logic; attribute dont_touch of WX629: signal is true;
	signal WX630: std_logic; attribute dont_touch of WX630: signal is true;
	signal WX631: std_logic; attribute dont_touch of WX631: signal is true;
	signal WX632: std_logic; attribute dont_touch of WX632: signal is true;
	signal WX633: std_logic; attribute dont_touch of WX633: signal is true;
	signal WX634: std_logic; attribute dont_touch of WX634: signal is true;
	signal WX635: std_logic; attribute dont_touch of WX635: signal is true;
	signal WX636: std_logic; attribute dont_touch of WX636: signal is true;
	signal WX637: std_logic; attribute dont_touch of WX637: signal is true;
	signal WX638: std_logic; attribute dont_touch of WX638: signal is true;
	signal WX639: std_logic; attribute dont_touch of WX639: signal is true;
	signal WX640: std_logic; attribute dont_touch of WX640: signal is true;
	signal WX641: std_logic; attribute dont_touch of WX641: signal is true;
	signal WX642: std_logic; attribute dont_touch of WX642: signal is true;
	signal WX643: std_logic; attribute dont_touch of WX643: signal is true;
	signal WX644: std_logic; attribute dont_touch of WX644: signal is true;
	signal WX645: std_logic; attribute dont_touch of WX645: signal is true;
	signal WX646: std_logic; attribute dont_touch of WX646: signal is true;
	signal WX647: std_logic; attribute dont_touch of WX647: signal is true;
	signal WX648: std_logic; attribute dont_touch of WX648: signal is true;
	signal WX649: std_logic; attribute dont_touch of WX649: signal is true;
	signal WX650: std_logic; attribute dont_touch of WX650: signal is true;
	signal WX651: std_logic; attribute dont_touch of WX651: signal is true;
	signal WX652: std_logic; attribute dont_touch of WX652: signal is true;
	signal WX653: std_logic; attribute dont_touch of WX653: signal is true;
	signal WX654: std_logic; attribute dont_touch of WX654: signal is true;
	signal WX655: std_logic; attribute dont_touch of WX655: signal is true;
	signal WX656: std_logic; attribute dont_touch of WX656: signal is true;
	signal WX657: std_logic; attribute dont_touch of WX657: signal is true;
	signal WX658: std_logic; attribute dont_touch of WX658: signal is true;
	signal WX659: std_logic; attribute dont_touch of WX659: signal is true;
	signal WX660: std_logic; attribute dont_touch of WX660: signal is true;
	signal WX661: std_logic; attribute dont_touch of WX661: signal is true;
	signal WX662: std_logic; attribute dont_touch of WX662: signal is true;
	signal WX663: std_logic; attribute dont_touch of WX663: signal is true;
	signal WX664: std_logic; attribute dont_touch of WX664: signal is true;
	signal WX665: std_logic; attribute dont_touch of WX665: signal is true;
	signal WX666: std_logic; attribute dont_touch of WX666: signal is true;
	signal WX667: std_logic; attribute dont_touch of WX667: signal is true;
	signal WX668: std_logic; attribute dont_touch of WX668: signal is true;
	signal WX669: std_logic; attribute dont_touch of WX669: signal is true;
	signal WX670: std_logic; attribute dont_touch of WX670: signal is true;
	signal WX671: std_logic; attribute dont_touch of WX671: signal is true;
	signal WX672: std_logic; attribute dont_touch of WX672: signal is true;
	signal WX673: std_logic; attribute dont_touch of WX673: signal is true;
	signal WX674: std_logic; attribute dont_touch of WX674: signal is true;
	signal WX675: std_logic; attribute dont_touch of WX675: signal is true;
	signal WX676: std_logic; attribute dont_touch of WX676: signal is true;
	signal WX677: std_logic; attribute dont_touch of WX677: signal is true;
	signal WX678: std_logic; attribute dont_touch of WX678: signal is true;
	signal WX679: std_logic; attribute dont_touch of WX679: signal is true;
	signal WX680: std_logic; attribute dont_touch of WX680: signal is true;
	signal WX681: std_logic; attribute dont_touch of WX681: signal is true;
	signal WX682: std_logic; attribute dont_touch of WX682: signal is true;
	signal WX683: std_logic; attribute dont_touch of WX683: signal is true;
	signal WX684: std_logic; attribute dont_touch of WX684: signal is true;
	signal WX685: std_logic; attribute dont_touch of WX685: signal is true;
	signal WX686: std_logic; attribute dont_touch of WX686: signal is true;
	signal WX687: std_logic; attribute dont_touch of WX687: signal is true;
	signal WX688: std_logic; attribute dont_touch of WX688: signal is true;
	signal WX689: std_logic; attribute dont_touch of WX689: signal is true;
	signal WX690: std_logic; attribute dont_touch of WX690: signal is true;
	signal WX691: std_logic; attribute dont_touch of WX691: signal is true;
	signal WX692: std_logic; attribute dont_touch of WX692: signal is true;
	signal WX693: std_logic; attribute dont_touch of WX693: signal is true;
	signal WX694: std_logic; attribute dont_touch of WX694: signal is true;
	signal WX695: std_logic; attribute dont_touch of WX695: signal is true;
	signal WX696: std_logic; attribute dont_touch of WX696: signal is true;
	signal WX697: std_logic; attribute dont_touch of WX697: signal is true;
	signal WX698: std_logic; attribute dont_touch of WX698: signal is true;
	signal WX699: std_logic; attribute dont_touch of WX699: signal is true;
	signal WX700: std_logic; attribute dont_touch of WX700: signal is true;
	signal WX701: std_logic; attribute dont_touch of WX701: signal is true;
	signal WX702: std_logic; attribute dont_touch of WX702: signal is true;
	signal WX703: std_logic; attribute dont_touch of WX703: signal is true;
	signal WX704: std_logic; attribute dont_touch of WX704: signal is true;
	signal WX705: std_logic; attribute dont_touch of WX705: signal is true;
	signal WX706: std_logic; attribute dont_touch of WX706: signal is true;
	signal WX707: std_logic; attribute dont_touch of WX707: signal is true;
	signal WX708: std_logic; attribute dont_touch of WX708: signal is true;
	signal WX709: std_logic; attribute dont_touch of WX709: signal is true;
	signal WX710: std_logic; attribute dont_touch of WX710: signal is true;
	signal WX711: std_logic; attribute dont_touch of WX711: signal is true;
	signal WX712: std_logic; attribute dont_touch of WX712: signal is true;
	signal WX713: std_logic; attribute dont_touch of WX713: signal is true;
	signal WX714: std_logic; attribute dont_touch of WX714: signal is true;
	signal WX715: std_logic; attribute dont_touch of WX715: signal is true;
	signal WX716: std_logic; attribute dont_touch of WX716: signal is true;
	signal WX717: std_logic; attribute dont_touch of WX717: signal is true;
	signal WX718: std_logic; attribute dont_touch of WX718: signal is true;
	signal WX719: std_logic; attribute dont_touch of WX719: signal is true;
	signal WX720: std_logic; attribute dont_touch of WX720: signal is true;
	signal WX721: std_logic; attribute dont_touch of WX721: signal is true;
	signal WX722: std_logic; attribute dont_touch of WX722: signal is true;
	signal WX723: std_logic; attribute dont_touch of WX723: signal is true;
	signal WX724: std_logic; attribute dont_touch of WX724: signal is true;
	signal WX725: std_logic; attribute dont_touch of WX725: signal is true;
	signal WX726: std_logic; attribute dont_touch of WX726: signal is true;
	signal WX727: std_logic; attribute dont_touch of WX727: signal is true;
	signal WX728: std_logic; attribute dont_touch of WX728: signal is true;
	signal WX729: std_logic; attribute dont_touch of WX729: signal is true;
	signal WX730: std_logic; attribute dont_touch of WX730: signal is true;
	signal WX731: std_logic; attribute dont_touch of WX731: signal is true;
	signal WX732: std_logic; attribute dont_touch of WX732: signal is true;
	signal WX733: std_logic; attribute dont_touch of WX733: signal is true;
	signal WX734: std_logic; attribute dont_touch of WX734: signal is true;
	signal WX735: std_logic; attribute dont_touch of WX735: signal is true;
	signal WX736: std_logic; attribute dont_touch of WX736: signal is true;
	signal WX737: std_logic; attribute dont_touch of WX737: signal is true;
	signal WX738: std_logic; attribute dont_touch of WX738: signal is true;
	signal WX739: std_logic; attribute dont_touch of WX739: signal is true;
	signal WX740: std_logic; attribute dont_touch of WX740: signal is true;
	signal WX741: std_logic; attribute dont_touch of WX741: signal is true;
	signal WX742: std_logic; attribute dont_touch of WX742: signal is true;
	signal WX743: std_logic; attribute dont_touch of WX743: signal is true;
	signal WX744: std_logic; attribute dont_touch of WX744: signal is true;
	signal WX745: std_logic; attribute dont_touch of WX745: signal is true;
	signal WX746: std_logic; attribute dont_touch of WX746: signal is true;
	signal WX747: std_logic; attribute dont_touch of WX747: signal is true;
	signal WX748: std_logic; attribute dont_touch of WX748: signal is true;
	signal WX749: std_logic; attribute dont_touch of WX749: signal is true;
	signal WX750: std_logic; attribute dont_touch of WX750: signal is true;
	signal WX751: std_logic; attribute dont_touch of WX751: signal is true;
	signal WX752: std_logic; attribute dont_touch of WX752: signal is true;
	signal WX753: std_logic; attribute dont_touch of WX753: signal is true;
	signal WX754: std_logic; attribute dont_touch of WX754: signal is true;
	signal WX755: std_logic; attribute dont_touch of WX755: signal is true;
	signal WX756: std_logic; attribute dont_touch of WX756: signal is true;
	signal WX757: std_logic; attribute dont_touch of WX757: signal is true;
	signal WX758: std_logic; attribute dont_touch of WX758: signal is true;
	signal WX759: std_logic; attribute dont_touch of WX759: signal is true;
	signal WX760: std_logic; attribute dont_touch of WX760: signal is true;
	signal WX761: std_logic; attribute dont_touch of WX761: signal is true;
	signal WX762: std_logic; attribute dont_touch of WX762: signal is true;
	signal WX763: std_logic; attribute dont_touch of WX763: signal is true;
	signal WX764: std_logic; attribute dont_touch of WX764: signal is true;
	signal WX765: std_logic; attribute dont_touch of WX765: signal is true;
	signal WX766: std_logic; attribute dont_touch of WX766: signal is true;
	signal WX767: std_logic; attribute dont_touch of WX767: signal is true;
	signal WX768: std_logic; attribute dont_touch of WX768: signal is true;
	signal WX769: std_logic; attribute dont_touch of WX769: signal is true;
	signal WX770: std_logic; attribute dont_touch of WX770: signal is true;
	signal WX771: std_logic; attribute dont_touch of WX771: signal is true;
	signal WX772: std_logic; attribute dont_touch of WX772: signal is true;
	signal WX773: std_logic; attribute dont_touch of WX773: signal is true;
	signal WX774: std_logic; attribute dont_touch of WX774: signal is true;
	signal WX775: std_logic; attribute dont_touch of WX775: signal is true;
	signal WX776: std_logic; attribute dont_touch of WX776: signal is true;
	signal WX777: std_logic; attribute dont_touch of WX777: signal is true;
	signal WX778: std_logic; attribute dont_touch of WX778: signal is true;
	signal WX779: std_logic; attribute dont_touch of WX779: signal is true;
	signal WX780: std_logic; attribute dont_touch of WX780: signal is true;
	signal WX781: std_logic; attribute dont_touch of WX781: signal is true;
	signal WX782: std_logic; attribute dont_touch of WX782: signal is true;
	signal WX783: std_logic; attribute dont_touch of WX783: signal is true;
	signal WX784: std_logic; attribute dont_touch of WX784: signal is true;
	signal WX785: std_logic; attribute dont_touch of WX785: signal is true;
	signal WX786: std_logic; attribute dont_touch of WX786: signal is true;
	signal WX787: std_logic; attribute dont_touch of WX787: signal is true;
	signal WX788: std_logic; attribute dont_touch of WX788: signal is true;
	signal WX789: std_logic; attribute dont_touch of WX789: signal is true;
	signal WX790: std_logic; attribute dont_touch of WX790: signal is true;
	signal WX791: std_logic; attribute dont_touch of WX791: signal is true;
	signal WX792: std_logic; attribute dont_touch of WX792: signal is true;
	signal WX793: std_logic; attribute dont_touch of WX793: signal is true;
	signal WX794: std_logic; attribute dont_touch of WX794: signal is true;
	signal WX795: std_logic; attribute dont_touch of WX795: signal is true;
	signal WX796: std_logic; attribute dont_touch of WX796: signal is true;
	signal WX797: std_logic; attribute dont_touch of WX797: signal is true;
	signal WX798: std_logic; attribute dont_touch of WX798: signal is true;
	signal WX799: std_logic; attribute dont_touch of WX799: signal is true;
	signal WX800: std_logic; attribute dont_touch of WX800: signal is true;
	signal WX801: std_logic; attribute dont_touch of WX801: signal is true;
	signal WX802: std_logic; attribute dont_touch of WX802: signal is true;
	signal WX803: std_logic; attribute dont_touch of WX803: signal is true;
	signal WX804: std_logic; attribute dont_touch of WX804: signal is true;
	signal WX805: std_logic; attribute dont_touch of WX805: signal is true;
	signal WX806: std_logic; attribute dont_touch of WX806: signal is true;
	signal WX807: std_logic; attribute dont_touch of WX807: signal is true;
	signal WX808: std_logic; attribute dont_touch of WX808: signal is true;
	signal WX809: std_logic; attribute dont_touch of WX809: signal is true;
	signal WX810: std_logic; attribute dont_touch of WX810: signal is true;
	signal WX811: std_logic; attribute dont_touch of WX811: signal is true;
	signal WX812: std_logic; attribute dont_touch of WX812: signal is true;
	signal WX813: std_logic; attribute dont_touch of WX813: signal is true;
	signal WX814: std_logic; attribute dont_touch of WX814: signal is true;
	signal WX815: std_logic; attribute dont_touch of WX815: signal is true;
	signal WX816: std_logic; attribute dont_touch of WX816: signal is true;
	signal WX817: std_logic; attribute dont_touch of WX817: signal is true;
	signal WX818: std_logic; attribute dont_touch of WX818: signal is true;
	signal WX819: std_logic; attribute dont_touch of WX819: signal is true;
	signal WX820: std_logic; attribute dont_touch of WX820: signal is true;
	signal WX821: std_logic; attribute dont_touch of WX821: signal is true;
	signal WX822: std_logic; attribute dont_touch of WX822: signal is true;
	signal WX823: std_logic; attribute dont_touch of WX823: signal is true;
	signal WX824: std_logic; attribute dont_touch of WX824: signal is true;
	signal WX825: std_logic; attribute dont_touch of WX825: signal is true;
	signal WX826: std_logic; attribute dont_touch of WX826: signal is true;
	signal WX827: std_logic; attribute dont_touch of WX827: signal is true;
	signal WX828: std_logic; attribute dont_touch of WX828: signal is true;
	signal WX829: std_logic; attribute dont_touch of WX829: signal is true;
	signal WX830: std_logic; attribute dont_touch of WX830: signal is true;
	signal WX831: std_logic; attribute dont_touch of WX831: signal is true;
	signal WX832: std_logic; attribute dont_touch of WX832: signal is true;
	signal WX833: std_logic; attribute dont_touch of WX833: signal is true;
	signal WX834: std_logic; attribute dont_touch of WX834: signal is true;
	signal WX835: std_logic; attribute dont_touch of WX835: signal is true;
	signal WX836: std_logic; attribute dont_touch of WX836: signal is true;
	signal WX837: std_logic; attribute dont_touch of WX837: signal is true;
	signal WX838: std_logic; attribute dont_touch of WX838: signal is true;
	signal WX839: std_logic; attribute dont_touch of WX839: signal is true;
	signal WX840: std_logic; attribute dont_touch of WX840: signal is true;
	signal WX841: std_logic; attribute dont_touch of WX841: signal is true;
	signal WX842: std_logic; attribute dont_touch of WX842: signal is true;
	signal WX843: std_logic; attribute dont_touch of WX843: signal is true;
	signal WX844: std_logic; attribute dont_touch of WX844: signal is true;
	signal WX845: std_logic; attribute dont_touch of WX845: signal is true;
	signal WX846: std_logic; attribute dont_touch of WX846: signal is true;
	signal WX847: std_logic; attribute dont_touch of WX847: signal is true;
	signal WX848: std_logic; attribute dont_touch of WX848: signal is true;
	signal WX849: std_logic; attribute dont_touch of WX849: signal is true;
	signal WX850: std_logic; attribute dont_touch of WX850: signal is true;
	signal WX851: std_logic; attribute dont_touch of WX851: signal is true;
	signal WX852: std_logic; attribute dont_touch of WX852: signal is true;
	signal WX853: std_logic; attribute dont_touch of WX853: signal is true;
	signal WX854: std_logic; attribute dont_touch of WX854: signal is true;
	signal WX855: std_logic; attribute dont_touch of WX855: signal is true;
	signal WX856: std_logic; attribute dont_touch of WX856: signal is true;
	signal WX857: std_logic; attribute dont_touch of WX857: signal is true;
	signal WX858: std_logic; attribute dont_touch of WX858: signal is true;
	signal WX859: std_logic; attribute dont_touch of WX859: signal is true;
	signal WX860: std_logic; attribute dont_touch of WX860: signal is true;
	signal WX861: std_logic; attribute dont_touch of WX861: signal is true;
	signal WX862: std_logic; attribute dont_touch of WX862: signal is true;
	signal WX863: std_logic; attribute dont_touch of WX863: signal is true;
	signal WX864: std_logic; attribute dont_touch of WX864: signal is true;
	signal WX865: std_logic; attribute dont_touch of WX865: signal is true;
	signal WX866: std_logic; attribute dont_touch of WX866: signal is true;
	signal WX867: std_logic; attribute dont_touch of WX867: signal is true;
	signal WX868: std_logic; attribute dont_touch of WX868: signal is true;
	signal WX869: std_logic; attribute dont_touch of WX869: signal is true;
	signal WX870: std_logic; attribute dont_touch of WX870: signal is true;
	signal WX871: std_logic; attribute dont_touch of WX871: signal is true;
	signal WX872: std_logic; attribute dont_touch of WX872: signal is true;
	signal WX873: std_logic; attribute dont_touch of WX873: signal is true;
	signal WX874: std_logic; attribute dont_touch of WX874: signal is true;
	signal WX875: std_logic; attribute dont_touch of WX875: signal is true;
	signal WX876: std_logic; attribute dont_touch of WX876: signal is true;
	signal WX877: std_logic; attribute dont_touch of WX877: signal is true;
	signal WX878: std_logic; attribute dont_touch of WX878: signal is true;
	signal WX879: std_logic; attribute dont_touch of WX879: signal is true;
	signal WX880: std_logic; attribute dont_touch of WX880: signal is true;
	signal WX881: std_logic; attribute dont_touch of WX881: signal is true;
	signal WX882: std_logic; attribute dont_touch of WX882: signal is true;
	signal WX883: std_logic; attribute dont_touch of WX883: signal is true;
	signal WX884: std_logic; attribute dont_touch of WX884: signal is true;
	signal WX885: std_logic; attribute dont_touch of WX885: signal is true;
	signal WX886: std_logic; attribute dont_touch of WX886: signal is true;
	signal WX887: std_logic; attribute dont_touch of WX887: signal is true;
	signal WX888: std_logic; attribute dont_touch of WX888: signal is true;
	signal WX889: std_logic; attribute dont_touch of WX889: signal is true;
	signal WX890: std_logic; attribute dont_touch of WX890: signal is true;
	signal WX891: std_logic; attribute dont_touch of WX891: signal is true;
	signal WX892: std_logic; attribute dont_touch of WX892: signal is true;
	signal WX893: std_logic; attribute dont_touch of WX893: signal is true;
	signal WX894: std_logic; attribute dont_touch of WX894: signal is true;
	signal WX895: std_logic; attribute dont_touch of WX895: signal is true;
	signal WX896: std_logic; attribute dont_touch of WX896: signal is true;
	signal WX897: std_logic; attribute dont_touch of WX897: signal is true;
	signal WX898: std_logic; attribute dont_touch of WX898: signal is true;
	signal WX899: std_logic; attribute dont_touch of WX899: signal is true;
	signal WX900: std_logic; attribute dont_touch of WX900: signal is true;
	signal WX901: std_logic; attribute dont_touch of WX901: signal is true;
	signal WX902: std_logic; attribute dont_touch of WX902: signal is true;
	signal WX903: std_logic; attribute dont_touch of WX903: signal is true;
	signal WX904: std_logic; attribute dont_touch of WX904: signal is true;
	signal WX905: std_logic; attribute dont_touch of WX905: signal is true;
	signal WX906: std_logic; attribute dont_touch of WX906: signal is true;
	signal WX907: std_logic; attribute dont_touch of WX907: signal is true;
	signal WX908: std_logic; attribute dont_touch of WX908: signal is true;
	signal WX909: std_logic; attribute dont_touch of WX909: signal is true;
	signal WX910: std_logic; attribute dont_touch of WX910: signal is true;
	signal WX911: std_logic; attribute dont_touch of WX911: signal is true;
	signal WX912: std_logic; attribute dont_touch of WX912: signal is true;
	signal WX913: std_logic; attribute dont_touch of WX913: signal is true;
	signal WX914: std_logic; attribute dont_touch of WX914: signal is true;
	signal WX915: std_logic; attribute dont_touch of WX915: signal is true;
	signal WX916: std_logic; attribute dont_touch of WX916: signal is true;
	signal WX917: std_logic; attribute dont_touch of WX917: signal is true;
	signal WX918: std_logic; attribute dont_touch of WX918: signal is true;
	signal WX919: std_logic; attribute dont_touch of WX919: signal is true;
	signal WX920: std_logic; attribute dont_touch of WX920: signal is true;
	signal WX921: std_logic; attribute dont_touch of WX921: signal is true;
	signal WX922: std_logic; attribute dont_touch of WX922: signal is true;
	signal WX923: std_logic; attribute dont_touch of WX923: signal is true;
	signal WX924: std_logic; attribute dont_touch of WX924: signal is true;
	signal WX925: std_logic; attribute dont_touch of WX925: signal is true;
	signal WX926: std_logic; attribute dont_touch of WX926: signal is true;
	signal WX927: std_logic; attribute dont_touch of WX927: signal is true;
	signal WX928: std_logic; attribute dont_touch of WX928: signal is true;
	signal WX929: std_logic; attribute dont_touch of WX929: signal is true;
	signal WX930: std_logic; attribute dont_touch of WX930: signal is true;
	signal WX931: std_logic; attribute dont_touch of WX931: signal is true;
	signal WX932: std_logic; attribute dont_touch of WX932: signal is true;
	signal WX933: std_logic; attribute dont_touch of WX933: signal is true;
	signal WX934: std_logic; attribute dont_touch of WX934: signal is true;
	signal WX935: std_logic; attribute dont_touch of WX935: signal is true;
	signal WX936: std_logic; attribute dont_touch of WX936: signal is true;
	signal WX937: std_logic; attribute dont_touch of WX937: signal is true;
	signal WX938: std_logic; attribute dont_touch of WX938: signal is true;
	signal WX939: std_logic; attribute dont_touch of WX939: signal is true;
	signal WX940: std_logic; attribute dont_touch of WX940: signal is true;
	signal WX941: std_logic; attribute dont_touch of WX941: signal is true;
	signal WX942: std_logic; attribute dont_touch of WX942: signal is true;
	signal WX943: std_logic; attribute dont_touch of WX943: signal is true;
	signal WX944: std_logic; attribute dont_touch of WX944: signal is true;
	signal WX945: std_logic; attribute dont_touch of WX945: signal is true;
	signal WX946: std_logic; attribute dont_touch of WX946: signal is true;
	signal WX947: std_logic; attribute dont_touch of WX947: signal is true;
	signal WX948: std_logic; attribute dont_touch of WX948: signal is true;
	signal WX949: std_logic; attribute dont_touch of WX949: signal is true;
	signal WX950: std_logic; attribute dont_touch of WX950: signal is true;
	signal WX951: std_logic; attribute dont_touch of WX951: signal is true;
	signal WX952: std_logic; attribute dont_touch of WX952: signal is true;
	signal WX953: std_logic; attribute dont_touch of WX953: signal is true;
	signal WX954: std_logic; attribute dont_touch of WX954: signal is true;
	signal WX955: std_logic; attribute dont_touch of WX955: signal is true;
	signal WX956: std_logic; attribute dont_touch of WX956: signal is true;
	signal WX957: std_logic; attribute dont_touch of WX957: signal is true;
	signal WX958: std_logic; attribute dont_touch of WX958: signal is true;
	signal WX959: std_logic; attribute dont_touch of WX959: signal is true;
	signal WX960: std_logic; attribute dont_touch of WX960: signal is true;
	signal WX961: std_logic; attribute dont_touch of WX961: signal is true;
	signal WX962: std_logic; attribute dont_touch of WX962: signal is true;
	signal WX963: std_logic; attribute dont_touch of WX963: signal is true;
	signal WX964: std_logic; attribute dont_touch of WX964: signal is true;
	signal WX965: std_logic; attribute dont_touch of WX965: signal is true;
	signal WX966: std_logic; attribute dont_touch of WX966: signal is true;
	signal WX967: std_logic; attribute dont_touch of WX967: signal is true;
	signal WX968: std_logic; attribute dont_touch of WX968: signal is true;
	signal WX969: std_logic; attribute dont_touch of WX969: signal is true;
	signal WX970: std_logic; attribute dont_touch of WX970: signal is true;
	signal WX971: std_logic; attribute dont_touch of WX971: signal is true;
	signal WX972: std_logic; attribute dont_touch of WX972: signal is true;
	signal WX973: std_logic; attribute dont_touch of WX973: signal is true;
	signal WX974: std_logic; attribute dont_touch of WX974: signal is true;
	signal WX975: std_logic; attribute dont_touch of WX975: signal is true;
	signal WX976: std_logic; attribute dont_touch of WX976: signal is true;
	signal WX977: std_logic; attribute dont_touch of WX977: signal is true;
	signal WX978: std_logic; attribute dont_touch of WX978: signal is true;
	signal WX979: std_logic; attribute dont_touch of WX979: signal is true;
	signal WX980: std_logic; attribute dont_touch of WX980: signal is true;
	signal WX981: std_logic; attribute dont_touch of WX981: signal is true;
	signal WX982: std_logic; attribute dont_touch of WX982: signal is true;
	signal WX983: std_logic; attribute dont_touch of WX983: signal is true;
	signal WX984: std_logic; attribute dont_touch of WX984: signal is true;
	signal WX985: std_logic; attribute dont_touch of WX985: signal is true;
	signal WX986: std_logic; attribute dont_touch of WX986: signal is true;
	signal WX987: std_logic; attribute dont_touch of WX987: signal is true;
	signal WX988: std_logic; attribute dont_touch of WX988: signal is true;
	signal WX989: std_logic; attribute dont_touch of WX989: signal is true;
	signal WX990: std_logic; attribute dont_touch of WX990: signal is true;
	signal WX991: std_logic; attribute dont_touch of WX991: signal is true;
	signal WX992: std_logic; attribute dont_touch of WX992: signal is true;
	signal WX993: std_logic; attribute dont_touch of WX993: signal is true;
	signal WX994: std_logic; attribute dont_touch of WX994: signal is true;
	signal WX995: std_logic; attribute dont_touch of WX995: signal is true;
	signal WX996: std_logic; attribute dont_touch of WX996: signal is true;
	signal WX997: std_logic; attribute dont_touch of WX997: signal is true;
	signal WX998: std_logic; attribute dont_touch of WX998: signal is true;
	signal WX999: std_logic; attribute dont_touch of WX999: signal is true;
	signal WX1000: std_logic; attribute dont_touch of WX1000: signal is true;
	signal WX1001: std_logic; attribute dont_touch of WX1001: signal is true;
	signal WX1002: std_logic; attribute dont_touch of WX1002: signal is true;
	signal WX1003: std_logic; attribute dont_touch of WX1003: signal is true;
	signal WX1004: std_logic; attribute dont_touch of WX1004: signal is true;
	signal WX1005: std_logic; attribute dont_touch of WX1005: signal is true;
	signal WX1006: std_logic; attribute dont_touch of WX1006: signal is true;
	signal WX1007: std_logic; attribute dont_touch of WX1007: signal is true;
	signal WX1008: std_logic; attribute dont_touch of WX1008: signal is true;
	signal WX1009: std_logic; attribute dont_touch of WX1009: signal is true;
	signal WX1010: std_logic; attribute dont_touch of WX1010: signal is true;
	signal WX1011: std_logic; attribute dont_touch of WX1011: signal is true;
	signal WX1013: std_logic; attribute dont_touch of WX1013: signal is true;
	signal WX1014: std_logic; attribute dont_touch of WX1014: signal is true;
	signal WX1015: std_logic; attribute dont_touch of WX1015: signal is true;
	signal WX1016: std_logic; attribute dont_touch of WX1016: signal is true;
	signal WX1017: std_logic; attribute dont_touch of WX1017: signal is true;
	signal WX1018: std_logic; attribute dont_touch of WX1018: signal is true;
	signal WX1020: std_logic; attribute dont_touch of WX1020: signal is true;
	signal WX1021: std_logic; attribute dont_touch of WX1021: signal is true;
	signal WX1022: std_logic; attribute dont_touch of WX1022: signal is true;
	signal WX1023: std_logic; attribute dont_touch of WX1023: signal is true;
	signal WX1024: std_logic; attribute dont_touch of WX1024: signal is true;
	signal WX1025: std_logic; attribute dont_touch of WX1025: signal is true;
	signal WX1027: std_logic; attribute dont_touch of WX1027: signal is true;
	signal WX1028: std_logic; attribute dont_touch of WX1028: signal is true;
	signal WX1029: std_logic; attribute dont_touch of WX1029: signal is true;
	signal WX1030: std_logic; attribute dont_touch of WX1030: signal is true;
	signal WX1031: std_logic; attribute dont_touch of WX1031: signal is true;
	signal WX1032: std_logic; attribute dont_touch of WX1032: signal is true;
	signal WX1034: std_logic; attribute dont_touch of WX1034: signal is true;
	signal WX1035: std_logic; attribute dont_touch of WX1035: signal is true;
	signal WX1036: std_logic; attribute dont_touch of WX1036: signal is true;
	signal WX1037: std_logic; attribute dont_touch of WX1037: signal is true;
	signal WX1038: std_logic; attribute dont_touch of WX1038: signal is true;
	signal WX1039: std_logic; attribute dont_touch of WX1039: signal is true;
	signal WX1041: std_logic; attribute dont_touch of WX1041: signal is true;
	signal WX1042: std_logic; attribute dont_touch of WX1042: signal is true;
	signal WX1043: std_logic; attribute dont_touch of WX1043: signal is true;
	signal WX1044: std_logic; attribute dont_touch of WX1044: signal is true;
	signal WX1045: std_logic; attribute dont_touch of WX1045: signal is true;
	signal WX1046: std_logic; attribute dont_touch of WX1046: signal is true;
	signal WX1048: std_logic; attribute dont_touch of WX1048: signal is true;
	signal WX1049: std_logic; attribute dont_touch of WX1049: signal is true;
	signal WX1050: std_logic; attribute dont_touch of WX1050: signal is true;
	signal WX1051: std_logic; attribute dont_touch of WX1051: signal is true;
	signal WX1052: std_logic; attribute dont_touch of WX1052: signal is true;
	signal WX1053: std_logic; attribute dont_touch of WX1053: signal is true;
	signal WX1055: std_logic; attribute dont_touch of WX1055: signal is true;
	signal WX1056: std_logic; attribute dont_touch of WX1056: signal is true;
	signal WX1057: std_logic; attribute dont_touch of WX1057: signal is true;
	signal WX1058: std_logic; attribute dont_touch of WX1058: signal is true;
	signal WX1059: std_logic; attribute dont_touch of WX1059: signal is true;
	signal WX1060: std_logic; attribute dont_touch of WX1060: signal is true;
	signal WX1062: std_logic; attribute dont_touch of WX1062: signal is true;
	signal WX1063: std_logic; attribute dont_touch of WX1063: signal is true;
	signal WX1064: std_logic; attribute dont_touch of WX1064: signal is true;
	signal WX1065: std_logic; attribute dont_touch of WX1065: signal is true;
	signal WX1066: std_logic; attribute dont_touch of WX1066: signal is true;
	signal WX1067: std_logic; attribute dont_touch of WX1067: signal is true;
	signal WX1069: std_logic; attribute dont_touch of WX1069: signal is true;
	signal WX1070: std_logic; attribute dont_touch of WX1070: signal is true;
	signal WX1071: std_logic; attribute dont_touch of WX1071: signal is true;
	signal WX1072: std_logic; attribute dont_touch of WX1072: signal is true;
	signal WX1073: std_logic; attribute dont_touch of WX1073: signal is true;
	signal WX1074: std_logic; attribute dont_touch of WX1074: signal is true;
	signal WX1076: std_logic; attribute dont_touch of WX1076: signal is true;
	signal WX1077: std_logic; attribute dont_touch of WX1077: signal is true;
	signal WX1078: std_logic; attribute dont_touch of WX1078: signal is true;
	signal WX1079: std_logic; attribute dont_touch of WX1079: signal is true;
	signal WX1080: std_logic; attribute dont_touch of WX1080: signal is true;
	signal WX1081: std_logic; attribute dont_touch of WX1081: signal is true;
	signal WX1083: std_logic; attribute dont_touch of WX1083: signal is true;
	signal WX1084: std_logic; attribute dont_touch of WX1084: signal is true;
	signal WX1085: std_logic; attribute dont_touch of WX1085: signal is true;
	signal WX1086: std_logic; attribute dont_touch of WX1086: signal is true;
	signal WX1087: std_logic; attribute dont_touch of WX1087: signal is true;
	signal WX1088: std_logic; attribute dont_touch of WX1088: signal is true;
	signal WX1090: std_logic; attribute dont_touch of WX1090: signal is true;
	signal WX1091: std_logic; attribute dont_touch of WX1091: signal is true;
	signal WX1092: std_logic; attribute dont_touch of WX1092: signal is true;
	signal WX1093: std_logic; attribute dont_touch of WX1093: signal is true;
	signal WX1094: std_logic; attribute dont_touch of WX1094: signal is true;
	signal WX1095: std_logic; attribute dont_touch of WX1095: signal is true;
	signal WX1097: std_logic; attribute dont_touch of WX1097: signal is true;
	signal WX1098: std_logic; attribute dont_touch of WX1098: signal is true;
	signal WX1099: std_logic; attribute dont_touch of WX1099: signal is true;
	signal WX1100: std_logic; attribute dont_touch of WX1100: signal is true;
	signal WX1101: std_logic; attribute dont_touch of WX1101: signal is true;
	signal WX1102: std_logic; attribute dont_touch of WX1102: signal is true;
	signal WX1104: std_logic; attribute dont_touch of WX1104: signal is true;
	signal WX1105: std_logic; attribute dont_touch of WX1105: signal is true;
	signal WX1106: std_logic; attribute dont_touch of WX1106: signal is true;
	signal WX1107: std_logic; attribute dont_touch of WX1107: signal is true;
	signal WX1108: std_logic; attribute dont_touch of WX1108: signal is true;
	signal WX1109: std_logic; attribute dont_touch of WX1109: signal is true;
	signal WX1111: std_logic; attribute dont_touch of WX1111: signal is true;
	signal WX1112: std_logic; attribute dont_touch of WX1112: signal is true;
	signal WX1113: std_logic; attribute dont_touch of WX1113: signal is true;
	signal WX1114: std_logic; attribute dont_touch of WX1114: signal is true;
	signal WX1115: std_logic; attribute dont_touch of WX1115: signal is true;
	signal WX1116: std_logic; attribute dont_touch of WX1116: signal is true;
	signal WX1118: std_logic; attribute dont_touch of WX1118: signal is true;
	signal WX1119: std_logic; attribute dont_touch of WX1119: signal is true;
	signal WX1120: std_logic; attribute dont_touch of WX1120: signal is true;
	signal WX1121: std_logic; attribute dont_touch of WX1121: signal is true;
	signal WX1122: std_logic; attribute dont_touch of WX1122: signal is true;
	signal WX1123: std_logic; attribute dont_touch of WX1123: signal is true;
	signal WX1125: std_logic; attribute dont_touch of WX1125: signal is true;
	signal WX1126: std_logic; attribute dont_touch of WX1126: signal is true;
	signal WX1127: std_logic; attribute dont_touch of WX1127: signal is true;
	signal WX1128: std_logic; attribute dont_touch of WX1128: signal is true;
	signal WX1129: std_logic; attribute dont_touch of WX1129: signal is true;
	signal WX1130: std_logic; attribute dont_touch of WX1130: signal is true;
	signal WX1132: std_logic; attribute dont_touch of WX1132: signal is true;
	signal WX1133: std_logic; attribute dont_touch of WX1133: signal is true;
	signal WX1134: std_logic; attribute dont_touch of WX1134: signal is true;
	signal WX1135: std_logic; attribute dont_touch of WX1135: signal is true;
	signal WX1136: std_logic; attribute dont_touch of WX1136: signal is true;
	signal WX1137: std_logic; attribute dont_touch of WX1137: signal is true;
	signal WX1139: std_logic; attribute dont_touch of WX1139: signal is true;
	signal WX1140: std_logic; attribute dont_touch of WX1140: signal is true;
	signal WX1141: std_logic; attribute dont_touch of WX1141: signal is true;
	signal WX1142: std_logic; attribute dont_touch of WX1142: signal is true;
	signal WX1143: std_logic; attribute dont_touch of WX1143: signal is true;
	signal WX1144: std_logic; attribute dont_touch of WX1144: signal is true;
	signal WX1146: std_logic; attribute dont_touch of WX1146: signal is true;
	signal WX1147: std_logic; attribute dont_touch of WX1147: signal is true;
	signal WX1148: std_logic; attribute dont_touch of WX1148: signal is true;
	signal WX1149: std_logic; attribute dont_touch of WX1149: signal is true;
	signal WX1150: std_logic; attribute dont_touch of WX1150: signal is true;
	signal WX1151: std_logic; attribute dont_touch of WX1151: signal is true;
	signal WX1153: std_logic; attribute dont_touch of WX1153: signal is true;
	signal WX1154: std_logic; attribute dont_touch of WX1154: signal is true;
	signal WX1155: std_logic; attribute dont_touch of WX1155: signal is true;
	signal WX1156: std_logic; attribute dont_touch of WX1156: signal is true;
	signal WX1157: std_logic; attribute dont_touch of WX1157: signal is true;
	signal WX1158: std_logic; attribute dont_touch of WX1158: signal is true;
	signal WX1160: std_logic; attribute dont_touch of WX1160: signal is true;
	signal WX1161: std_logic; attribute dont_touch of WX1161: signal is true;
	signal WX1162: std_logic; attribute dont_touch of WX1162: signal is true;
	signal WX1163: std_logic; attribute dont_touch of WX1163: signal is true;
	signal WX1164: std_logic; attribute dont_touch of WX1164: signal is true;
	signal WX1165: std_logic; attribute dont_touch of WX1165: signal is true;
	signal WX1167: std_logic; attribute dont_touch of WX1167: signal is true;
	signal WX1168: std_logic; attribute dont_touch of WX1168: signal is true;
	signal WX1169: std_logic; attribute dont_touch of WX1169: signal is true;
	signal WX1170: std_logic; attribute dont_touch of WX1170: signal is true;
	signal WX1171: std_logic; attribute dont_touch of WX1171: signal is true;
	signal WX1172: std_logic; attribute dont_touch of WX1172: signal is true;
	signal WX1174: std_logic; attribute dont_touch of WX1174: signal is true;
	signal WX1175: std_logic; attribute dont_touch of WX1175: signal is true;
	signal WX1176: std_logic; attribute dont_touch of WX1176: signal is true;
	signal WX1177: std_logic; attribute dont_touch of WX1177: signal is true;
	signal WX1178: std_logic; attribute dont_touch of WX1178: signal is true;
	signal WX1179: std_logic; attribute dont_touch of WX1179: signal is true;
	signal WX1181: std_logic; attribute dont_touch of WX1181: signal is true;
	signal WX1182: std_logic; attribute dont_touch of WX1182: signal is true;
	signal WX1183: std_logic; attribute dont_touch of WX1183: signal is true;
	signal WX1184: std_logic; attribute dont_touch of WX1184: signal is true;
	signal WX1185: std_logic; attribute dont_touch of WX1185: signal is true;
	signal WX1186: std_logic; attribute dont_touch of WX1186: signal is true;
	signal WX1188: std_logic; attribute dont_touch of WX1188: signal is true;
	signal WX1189: std_logic; attribute dont_touch of WX1189: signal is true;
	signal WX1190: std_logic; attribute dont_touch of WX1190: signal is true;
	signal WX1191: std_logic; attribute dont_touch of WX1191: signal is true;
	signal WX1192: std_logic; attribute dont_touch of WX1192: signal is true;
	signal WX1193: std_logic; attribute dont_touch of WX1193: signal is true;
	signal WX1195: std_logic; attribute dont_touch of WX1195: signal is true;
	signal WX1196: std_logic; attribute dont_touch of WX1196: signal is true;
	signal WX1197: std_logic; attribute dont_touch of WX1197: signal is true;
	signal WX1198: std_logic; attribute dont_touch of WX1198: signal is true;
	signal WX1199: std_logic; attribute dont_touch of WX1199: signal is true;
	signal WX1200: std_logic; attribute dont_touch of WX1200: signal is true;
	signal WX1202: std_logic; attribute dont_touch of WX1202: signal is true;
	signal WX1203: std_logic; attribute dont_touch of WX1203: signal is true;
	signal WX1204: std_logic; attribute dont_touch of WX1204: signal is true;
	signal WX1205: std_logic; attribute dont_touch of WX1205: signal is true;
	signal WX1206: std_logic; attribute dont_touch of WX1206: signal is true;
	signal WX1207: std_logic; attribute dont_touch of WX1207: signal is true;
	signal WX1209: std_logic; attribute dont_touch of WX1209: signal is true;
	signal WX1210: std_logic; attribute dont_touch of WX1210: signal is true;
	signal WX1211: std_logic; attribute dont_touch of WX1211: signal is true;
	signal WX1212: std_logic; attribute dont_touch of WX1212: signal is true;
	signal WX1213: std_logic; attribute dont_touch of WX1213: signal is true;
	signal WX1214: std_logic; attribute dont_touch of WX1214: signal is true;
	signal WX1216: std_logic; attribute dont_touch of WX1216: signal is true;
	signal WX1217: std_logic; attribute dont_touch of WX1217: signal is true;
	signal WX1218: std_logic; attribute dont_touch of WX1218: signal is true;
	signal WX1219: std_logic; attribute dont_touch of WX1219: signal is true;
	signal WX1220: std_logic; attribute dont_touch of WX1220: signal is true;
	signal WX1221: std_logic; attribute dont_touch of WX1221: signal is true;
	signal WX1223: std_logic; attribute dont_touch of WX1223: signal is true;
	signal WX1224: std_logic; attribute dont_touch of WX1224: signal is true;
	signal WX1225: std_logic; attribute dont_touch of WX1225: signal is true;
	signal WX1226: std_logic; attribute dont_touch of WX1226: signal is true;
	signal WX1227: std_logic; attribute dont_touch of WX1227: signal is true;
	signal WX1228: std_logic; attribute dont_touch of WX1228: signal is true;
	signal WX1230: std_logic; attribute dont_touch of WX1230: signal is true;
	signal WX1231: std_logic; attribute dont_touch of WX1231: signal is true;
	signal WX1232: std_logic; attribute dont_touch of WX1232: signal is true;
	signal WX1233: std_logic; attribute dont_touch of WX1233: signal is true;
	signal WX1234: std_logic; attribute dont_touch of WX1234: signal is true;
	signal WX1235: std_logic; attribute dont_touch of WX1235: signal is true;
	signal WX1236: std_logic; attribute dont_touch of WX1236: signal is true;
	signal WX1237: std_logic; attribute dont_touch of WX1237: signal is true;
	signal WX1238: std_logic; attribute dont_touch of WX1238: signal is true;
	signal WX1239: std_logic; attribute dont_touch of WX1239: signal is true;
	signal WX1240: std_logic; attribute dont_touch of WX1240: signal is true;
	signal WX1241: std_logic; attribute dont_touch of WX1241: signal is true;
	signal WX1242: std_logic; attribute dont_touch of WX1242: signal is true;
	signal WX1243: std_logic; attribute dont_touch of WX1243: signal is true;
	signal WX1244: std_logic; attribute dont_touch of WX1244: signal is true;
	signal WX1245: std_logic; attribute dont_touch of WX1245: signal is true;
	signal WX1246: std_logic; attribute dont_touch of WX1246: signal is true;
	signal WX1247: std_logic; attribute dont_touch of WX1247: signal is true;
	signal WX1248: std_logic; attribute dont_touch of WX1248: signal is true;
	signal WX1249: std_logic; attribute dont_touch of WX1249: signal is true;
	signal WX1250: std_logic; attribute dont_touch of WX1250: signal is true;
	signal WX1251: std_logic; attribute dont_touch of WX1251: signal is true;
	signal WX1252: std_logic; attribute dont_touch of WX1252: signal is true;
	signal WX1253: std_logic; attribute dont_touch of WX1253: signal is true;
	signal WX1254: std_logic; attribute dont_touch of WX1254: signal is true;
	signal WX1255: std_logic; attribute dont_touch of WX1255: signal is true;
	signal WX1256: std_logic; attribute dont_touch of WX1256: signal is true;
	signal WX1257: std_logic; attribute dont_touch of WX1257: signal is true;
	signal WX1258: std_logic; attribute dont_touch of WX1258: signal is true;
	signal WX1259: std_logic; attribute dont_touch of WX1259: signal is true;
	signal WX1260: std_logic; attribute dont_touch of WX1260: signal is true;
	signal WX1261: std_logic; attribute dont_touch of WX1261: signal is true;
	signal WX1262: std_logic; attribute dont_touch of WX1262: signal is true;
	signal WX1263: std_logic; attribute dont_touch of WX1263: signal is true;
	signal WX1264: std_logic; attribute dont_touch of WX1264: signal is true;
	signal WX1266: std_logic; attribute dont_touch of WX1266: signal is true;
	signal WX1268: std_logic; attribute dont_touch of WX1268: signal is true;
	signal WX1270: std_logic; attribute dont_touch of WX1270: signal is true;
	signal WX1272: std_logic; attribute dont_touch of WX1272: signal is true;
	signal WX1274: std_logic; attribute dont_touch of WX1274: signal is true;
	signal WX1276: std_logic; attribute dont_touch of WX1276: signal is true;
	signal WX1278: std_logic; attribute dont_touch of WX1278: signal is true;
	signal WX1280: std_logic; attribute dont_touch of WX1280: signal is true;
	signal WX1282: std_logic; attribute dont_touch of WX1282: signal is true;
	signal WX1284: std_logic; attribute dont_touch of WX1284: signal is true;
	signal WX1286: std_logic; attribute dont_touch of WX1286: signal is true;
	signal WX1288: std_logic; attribute dont_touch of WX1288: signal is true;
	signal WX1290: std_logic; attribute dont_touch of WX1290: signal is true;
	signal WX1292: std_logic; attribute dont_touch of WX1292: signal is true;
	signal WX1294: std_logic; attribute dont_touch of WX1294: signal is true;
	signal WX1296: std_logic; attribute dont_touch of WX1296: signal is true;
	signal WX1298: std_logic; attribute dont_touch of WX1298: signal is true;
	signal WX1300: std_logic; attribute dont_touch of WX1300: signal is true;
	signal WX1302: std_logic; attribute dont_touch of WX1302: signal is true;
	signal WX1304: std_logic; attribute dont_touch of WX1304: signal is true;
	signal WX1306: std_logic; attribute dont_touch of WX1306: signal is true;
	signal WX1308: std_logic; attribute dont_touch of WX1308: signal is true;
	signal WX1310: std_logic; attribute dont_touch of WX1310: signal is true;
	signal WX1312: std_logic; attribute dont_touch of WX1312: signal is true;
	signal WX1314: std_logic; attribute dont_touch of WX1314: signal is true;
	signal WX1316: std_logic; attribute dont_touch of WX1316: signal is true;
	signal WX1318: std_logic; attribute dont_touch of WX1318: signal is true;
	signal WX1320: std_logic; attribute dont_touch of WX1320: signal is true;
	signal WX1322: std_logic; attribute dont_touch of WX1322: signal is true;
	signal WX1324: std_logic; attribute dont_touch of WX1324: signal is true;
	signal WX1326: std_logic; attribute dont_touch of WX1326: signal is true;
	signal WX1328: std_logic; attribute dont_touch of WX1328: signal is true;
	signal WX1329: std_logic; attribute dont_touch of WX1329: signal is true;
	signal WX1330: std_logic; attribute dont_touch of WX1330: signal is true;
	signal WX1331: std_logic; attribute dont_touch of WX1331: signal is true;
	signal WX1332: std_logic; attribute dont_touch of WX1332: signal is true;
	signal WX1333: std_logic; attribute dont_touch of WX1333: signal is true;
	signal WX1334: std_logic; attribute dont_touch of WX1334: signal is true;
	signal WX1335: std_logic; attribute dont_touch of WX1335: signal is true;
	signal WX1336: std_logic; attribute dont_touch of WX1336: signal is true;
	signal WX1337: std_logic; attribute dont_touch of WX1337: signal is true;
	signal WX1338: std_logic; attribute dont_touch of WX1338: signal is true;
	signal WX1339: std_logic; attribute dont_touch of WX1339: signal is true;
	signal WX1340: std_logic; attribute dont_touch of WX1340: signal is true;
	signal WX1341: std_logic; attribute dont_touch of WX1341: signal is true;
	signal WX1342: std_logic; attribute dont_touch of WX1342: signal is true;
	signal WX1343: std_logic; attribute dont_touch of WX1343: signal is true;
	signal WX1344: std_logic; attribute dont_touch of WX1344: signal is true;
	signal WX1345: std_logic; attribute dont_touch of WX1345: signal is true;
	signal WX1346: std_logic; attribute dont_touch of WX1346: signal is true;
	signal WX1347: std_logic; attribute dont_touch of WX1347: signal is true;
	signal WX1348: std_logic; attribute dont_touch of WX1348: signal is true;
	signal WX1349: std_logic; attribute dont_touch of WX1349: signal is true;
	signal WX1350: std_logic; attribute dont_touch of WX1350: signal is true;
	signal WX1351: std_logic; attribute dont_touch of WX1351: signal is true;
	signal WX1352: std_logic; attribute dont_touch of WX1352: signal is true;
	signal WX1353: std_logic; attribute dont_touch of WX1353: signal is true;
	signal WX1354: std_logic; attribute dont_touch of WX1354: signal is true;
	signal WX1355: std_logic; attribute dont_touch of WX1355: signal is true;
	signal WX1356: std_logic; attribute dont_touch of WX1356: signal is true;
	signal WX1357: std_logic; attribute dont_touch of WX1357: signal is true;
	signal WX1358: std_logic; attribute dont_touch of WX1358: signal is true;
	signal WX1359: std_logic; attribute dont_touch of WX1359: signal is true;
	signal WX1360: std_logic; attribute dont_touch of WX1360: signal is true;
	signal WX1361: std_logic; attribute dont_touch of WX1361: signal is true;
	signal WX1362: std_logic; attribute dont_touch of WX1362: signal is true;
	signal WX1363: std_logic; attribute dont_touch of WX1363: signal is true;
	signal WX1364: std_logic; attribute dont_touch of WX1364: signal is true;
	signal WX1365: std_logic; attribute dont_touch of WX1365: signal is true;
	signal WX1366: std_logic; attribute dont_touch of WX1366: signal is true;
	signal WX1367: std_logic; attribute dont_touch of WX1367: signal is true;
	signal WX1368: std_logic; attribute dont_touch of WX1368: signal is true;
	signal WX1369: std_logic; attribute dont_touch of WX1369: signal is true;
	signal WX1370: std_logic; attribute dont_touch of WX1370: signal is true;
	signal WX1371: std_logic; attribute dont_touch of WX1371: signal is true;
	signal WX1372: std_logic; attribute dont_touch of WX1372: signal is true;
	signal WX1373: std_logic; attribute dont_touch of WX1373: signal is true;
	signal WX1374: std_logic; attribute dont_touch of WX1374: signal is true;
	signal WX1375: std_logic; attribute dont_touch of WX1375: signal is true;
	signal WX1376: std_logic; attribute dont_touch of WX1376: signal is true;
	signal WX1377: std_logic; attribute dont_touch of WX1377: signal is true;
	signal WX1378: std_logic; attribute dont_touch of WX1378: signal is true;
	signal WX1379: std_logic; attribute dont_touch of WX1379: signal is true;
	signal WX1380: std_logic; attribute dont_touch of WX1380: signal is true;
	signal WX1381: std_logic; attribute dont_touch of WX1381: signal is true;
	signal WX1382: std_logic; attribute dont_touch of WX1382: signal is true;
	signal WX1383: std_logic; attribute dont_touch of WX1383: signal is true;
	signal WX1384: std_logic; attribute dont_touch of WX1384: signal is true;
	signal WX1385: std_logic; attribute dont_touch of WX1385: signal is true;
	signal WX1386: std_logic; attribute dont_touch of WX1386: signal is true;
	signal WX1387: std_logic; attribute dont_touch of WX1387: signal is true;
	signal WX1388: std_logic; attribute dont_touch of WX1388: signal is true;
	signal WX1389: std_logic; attribute dont_touch of WX1389: signal is true;
	signal WX1390: std_logic; attribute dont_touch of WX1390: signal is true;
	signal WX1391: std_logic; attribute dont_touch of WX1391: signal is true;
	signal WX1392: std_logic; attribute dont_touch of WX1392: signal is true;
	signal WX1393: std_logic; attribute dont_touch of WX1393: signal is true;
	signal WX1394: std_logic; attribute dont_touch of WX1394: signal is true;
	signal WX1395: std_logic; attribute dont_touch of WX1395: signal is true;
	signal WX1396: std_logic; attribute dont_touch of WX1396: signal is true;
	signal WX1397: std_logic; attribute dont_touch of WX1397: signal is true;
	signal WX1398: std_logic; attribute dont_touch of WX1398: signal is true;
	signal WX1399: std_logic; attribute dont_touch of WX1399: signal is true;
	signal WX1400: std_logic; attribute dont_touch of WX1400: signal is true;
	signal WX1401: std_logic; attribute dont_touch of WX1401: signal is true;
	signal WX1402: std_logic; attribute dont_touch of WX1402: signal is true;
	signal WX1403: std_logic; attribute dont_touch of WX1403: signal is true;
	signal WX1404: std_logic; attribute dont_touch of WX1404: signal is true;
	signal WX1405: std_logic; attribute dont_touch of WX1405: signal is true;
	signal WX1406: std_logic; attribute dont_touch of WX1406: signal is true;
	signal WX1407: std_logic; attribute dont_touch of WX1407: signal is true;
	signal WX1408: std_logic; attribute dont_touch of WX1408: signal is true;
	signal WX1409: std_logic; attribute dont_touch of WX1409: signal is true;
	signal WX1410: std_logic; attribute dont_touch of WX1410: signal is true;
	signal WX1411: std_logic; attribute dont_touch of WX1411: signal is true;
	signal WX1412: std_logic; attribute dont_touch of WX1412: signal is true;
	signal WX1413: std_logic; attribute dont_touch of WX1413: signal is true;
	signal WX1414: std_logic; attribute dont_touch of WX1414: signal is true;
	signal WX1415: std_logic; attribute dont_touch of WX1415: signal is true;
	signal WX1416: std_logic; attribute dont_touch of WX1416: signal is true;
	signal WX1417: std_logic; attribute dont_touch of WX1417: signal is true;
	signal WX1418: std_logic; attribute dont_touch of WX1418: signal is true;
	signal WX1419: std_logic; attribute dont_touch of WX1419: signal is true;
	signal WX1420: std_logic; attribute dont_touch of WX1420: signal is true;
	signal WX1421: std_logic; attribute dont_touch of WX1421: signal is true;
	signal WX1422: std_logic; attribute dont_touch of WX1422: signal is true;
	signal WX1423: std_logic; attribute dont_touch of WX1423: signal is true;
	signal WX1424: std_logic; attribute dont_touch of WX1424: signal is true;
	signal WX1425: std_logic; attribute dont_touch of WX1425: signal is true;
	signal WX1426: std_logic; attribute dont_touch of WX1426: signal is true;
	signal WX1427: std_logic; attribute dont_touch of WX1427: signal is true;
	signal WX1428: std_logic; attribute dont_touch of WX1428: signal is true;
	signal WX1429: std_logic; attribute dont_touch of WX1429: signal is true;
	signal WX1430: std_logic; attribute dont_touch of WX1430: signal is true;
	signal WX1431: std_logic; attribute dont_touch of WX1431: signal is true;
	signal WX1432: std_logic; attribute dont_touch of WX1432: signal is true;
	signal WX1433: std_logic; attribute dont_touch of WX1433: signal is true;
	signal WX1434: std_logic; attribute dont_touch of WX1434: signal is true;
	signal WX1435: std_logic; attribute dont_touch of WX1435: signal is true;
	signal WX1436: std_logic; attribute dont_touch of WX1436: signal is true;
	signal WX1437: std_logic; attribute dont_touch of WX1437: signal is true;
	signal WX1438: std_logic; attribute dont_touch of WX1438: signal is true;
	signal WX1439: std_logic; attribute dont_touch of WX1439: signal is true;
	signal WX1440: std_logic; attribute dont_touch of WX1440: signal is true;
	signal WX1441: std_logic; attribute dont_touch of WX1441: signal is true;
	signal WX1442: std_logic; attribute dont_touch of WX1442: signal is true;
	signal WX1443: std_logic; attribute dont_touch of WX1443: signal is true;
	signal WX1444: std_logic; attribute dont_touch of WX1444: signal is true;
	signal WX1445: std_logic; attribute dont_touch of WX1445: signal is true;
	signal WX1446: std_logic; attribute dont_touch of WX1446: signal is true;
	signal WX1447: std_logic; attribute dont_touch of WX1447: signal is true;
	signal WX1448: std_logic; attribute dont_touch of WX1448: signal is true;
	signal WX1449: std_logic; attribute dont_touch of WX1449: signal is true;
	signal WX1450: std_logic; attribute dont_touch of WX1450: signal is true;
	signal WX1451: std_logic; attribute dont_touch of WX1451: signal is true;
	signal WX1452: std_logic; attribute dont_touch of WX1452: signal is true;
	signal WX1453: std_logic; attribute dont_touch of WX1453: signal is true;
	signal WX1454: std_logic; attribute dont_touch of WX1454: signal is true;
	signal WX1455: std_logic; attribute dont_touch of WX1455: signal is true;
	signal WX1456: std_logic; attribute dont_touch of WX1456: signal is true;
	signal WX1457: std_logic; attribute dont_touch of WX1457: signal is true;
	signal WX1458: std_logic; attribute dont_touch of WX1458: signal is true;
	signal WX1459: std_logic; attribute dont_touch of WX1459: signal is true;
	signal WX1460: std_logic; attribute dont_touch of WX1460: signal is true;
	signal WX1461: std_logic; attribute dont_touch of WX1461: signal is true;
	signal WX1462: std_logic; attribute dont_touch of WX1462: signal is true;
	signal WX1463: std_logic; attribute dont_touch of WX1463: signal is true;
	signal WX1464: std_logic; attribute dont_touch of WX1464: signal is true;
	signal WX1465: std_logic; attribute dont_touch of WX1465: signal is true;
	signal WX1466: std_logic; attribute dont_touch of WX1466: signal is true;
	signal WX1467: std_logic; attribute dont_touch of WX1467: signal is true;
	signal WX1468: std_logic; attribute dont_touch of WX1468: signal is true;
	signal WX1469: std_logic; attribute dont_touch of WX1469: signal is true;
	signal WX1470: std_logic; attribute dont_touch of WX1470: signal is true;
	signal WX1471: std_logic; attribute dont_touch of WX1471: signal is true;
	signal WX1472: std_logic; attribute dont_touch of WX1472: signal is true;
	signal WX1473: std_logic; attribute dont_touch of WX1473: signal is true;
	signal WX1474: std_logic; attribute dont_touch of WX1474: signal is true;
	signal WX1475: std_logic; attribute dont_touch of WX1475: signal is true;
	signal WX1476: std_logic; attribute dont_touch of WX1476: signal is true;
	signal WX1477: std_logic; attribute dont_touch of WX1477: signal is true;
	signal WX1478: std_logic; attribute dont_touch of WX1478: signal is true;
	signal WX1479: std_logic; attribute dont_touch of WX1479: signal is true;
	signal WX1480: std_logic; attribute dont_touch of WX1480: signal is true;
	signal WX1481: std_logic; attribute dont_touch of WX1481: signal is true;
	signal WX1482: std_logic; attribute dont_touch of WX1482: signal is true;
	signal WX1483: std_logic; attribute dont_touch of WX1483: signal is true;
	signal WX1484: std_logic; attribute dont_touch of WX1484: signal is true;
	signal WX1485: std_logic; attribute dont_touch of WX1485: signal is true;
	signal WX1486: std_logic; attribute dont_touch of WX1486: signal is true;
	signal WX1487: std_logic; attribute dont_touch of WX1487: signal is true;
	signal WX1488: std_logic; attribute dont_touch of WX1488: signal is true;
	signal WX1489: std_logic; attribute dont_touch of WX1489: signal is true;
	signal WX1490: std_logic; attribute dont_touch of WX1490: signal is true;
	signal WX1491: std_logic; attribute dont_touch of WX1491: signal is true;
	signal WX1492: std_logic; attribute dont_touch of WX1492: signal is true;
	signal WX1493: std_logic; attribute dont_touch of WX1493: signal is true;
	signal WX1494: std_logic; attribute dont_touch of WX1494: signal is true;
	signal WX1495: std_logic; attribute dont_touch of WX1495: signal is true;
	signal WX1496: std_logic; attribute dont_touch of WX1496: signal is true;
	signal WX1497: std_logic; attribute dont_touch of WX1497: signal is true;
	signal WX1498: std_logic; attribute dont_touch of WX1498: signal is true;
	signal WX1499: std_logic; attribute dont_touch of WX1499: signal is true;
	signal WX1500: std_logic; attribute dont_touch of WX1500: signal is true;
	signal WX1501: std_logic; attribute dont_touch of WX1501: signal is true;
	signal WX1502: std_logic; attribute dont_touch of WX1502: signal is true;
	signal WX1503: std_logic; attribute dont_touch of WX1503: signal is true;
	signal WX1504: std_logic; attribute dont_touch of WX1504: signal is true;
	signal WX1505: std_logic; attribute dont_touch of WX1505: signal is true;
	signal WX1506: std_logic; attribute dont_touch of WX1506: signal is true;
	signal WX1507: std_logic; attribute dont_touch of WX1507: signal is true;
	signal WX1508: std_logic; attribute dont_touch of WX1508: signal is true;
	signal WX1509: std_logic; attribute dont_touch of WX1509: signal is true;
	signal WX1510: std_logic; attribute dont_touch of WX1510: signal is true;
	signal WX1511: std_logic; attribute dont_touch of WX1511: signal is true;
	signal WX1512: std_logic; attribute dont_touch of WX1512: signal is true;
	signal WX1513: std_logic; attribute dont_touch of WX1513: signal is true;
	signal WX1514: std_logic; attribute dont_touch of WX1514: signal is true;
	signal WX1515: std_logic; attribute dont_touch of WX1515: signal is true;
	signal WX1516: std_logic; attribute dont_touch of WX1516: signal is true;
	signal WX1517: std_logic; attribute dont_touch of WX1517: signal is true;
	signal WX1518: std_logic; attribute dont_touch of WX1518: signal is true;
	signal WX1519: std_logic; attribute dont_touch of WX1519: signal is true;
	signal WX1520: std_logic; attribute dont_touch of WX1520: signal is true;
	signal WX1521: std_logic; attribute dont_touch of WX1521: signal is true;
	signal WX1522: std_logic; attribute dont_touch of WX1522: signal is true;
	signal WX1523: std_logic; attribute dont_touch of WX1523: signal is true;
	signal WX1524: std_logic; attribute dont_touch of WX1524: signal is true;
	signal WX1525: std_logic; attribute dont_touch of WX1525: signal is true;
	signal WX1526: std_logic; attribute dont_touch of WX1526: signal is true;
	signal WX1527: std_logic; attribute dont_touch of WX1527: signal is true;
	signal WX1528: std_logic; attribute dont_touch of WX1528: signal is true;
	signal WX1529: std_logic; attribute dont_touch of WX1529: signal is true;
	signal WX1530: std_logic; attribute dont_touch of WX1530: signal is true;
	signal WX1531: std_logic; attribute dont_touch of WX1531: signal is true;
	signal WX1532: std_logic; attribute dont_touch of WX1532: signal is true;
	signal WX1533: std_logic; attribute dont_touch of WX1533: signal is true;
	signal WX1534: std_logic; attribute dont_touch of WX1534: signal is true;
	signal WX1535: std_logic; attribute dont_touch of WX1535: signal is true;
	signal WX1536: std_logic; attribute dont_touch of WX1536: signal is true;
	signal WX1537: std_logic; attribute dont_touch of WX1537: signal is true;
	signal WX1538: std_logic; attribute dont_touch of WX1538: signal is true;
	signal WX1539: std_logic; attribute dont_touch of WX1539: signal is true;
	signal WX1540: std_logic; attribute dont_touch of WX1540: signal is true;
	signal WX1541: std_logic; attribute dont_touch of WX1541: signal is true;
	signal WX1542: std_logic; attribute dont_touch of WX1542: signal is true;
	signal WX1543: std_logic; attribute dont_touch of WX1543: signal is true;
	signal WX1544: std_logic; attribute dont_touch of WX1544: signal is true;
	signal WX1545: std_logic; attribute dont_touch of WX1545: signal is true;
	signal WX1546: std_logic; attribute dont_touch of WX1546: signal is true;
	signal WX1547: std_logic; attribute dont_touch of WX1547: signal is true;
	signal WX1548: std_logic; attribute dont_touch of WX1548: signal is true;
	signal WX1549: std_logic; attribute dont_touch of WX1549: signal is true;
	signal WX1550: std_logic; attribute dont_touch of WX1550: signal is true;
	signal WX1551: std_logic; attribute dont_touch of WX1551: signal is true;
	signal WX1552: std_logic; attribute dont_touch of WX1552: signal is true;
	signal WX1553: std_logic; attribute dont_touch of WX1553: signal is true;
	signal WX1554: std_logic; attribute dont_touch of WX1554: signal is true;
	signal WX1555: std_logic; attribute dont_touch of WX1555: signal is true;
	signal WX1556: std_logic; attribute dont_touch of WX1556: signal is true;
	signal WX1557: std_logic; attribute dont_touch of WX1557: signal is true;
	signal WX1558: std_logic; attribute dont_touch of WX1558: signal is true;
	signal WX1559: std_logic; attribute dont_touch of WX1559: signal is true;
	signal WX1560: std_logic; attribute dont_touch of WX1560: signal is true;
	signal WX1561: std_logic; attribute dont_touch of WX1561: signal is true;
	signal WX1562: std_logic; attribute dont_touch of WX1562: signal is true;
	signal WX1563: std_logic; attribute dont_touch of WX1563: signal is true;
	signal WX1564: std_logic; attribute dont_touch of WX1564: signal is true;
	signal WX1565: std_logic; attribute dont_touch of WX1565: signal is true;
	signal WX1566: std_logic; attribute dont_touch of WX1566: signal is true;
	signal WX1567: std_logic; attribute dont_touch of WX1567: signal is true;
	signal WX1568: std_logic; attribute dont_touch of WX1568: signal is true;
	signal WX1569: std_logic; attribute dont_touch of WX1569: signal is true;
	signal WX1570: std_logic; attribute dont_touch of WX1570: signal is true;
	signal WX1571: std_logic; attribute dont_touch of WX1571: signal is true;
	signal WX1572: std_logic; attribute dont_touch of WX1572: signal is true;
	signal WX1573: std_logic; attribute dont_touch of WX1573: signal is true;
	signal WX1574: std_logic; attribute dont_touch of WX1574: signal is true;
	signal WX1575: std_logic; attribute dont_touch of WX1575: signal is true;
	signal WX1576: std_logic; attribute dont_touch of WX1576: signal is true;
	signal WX1577: std_logic; attribute dont_touch of WX1577: signal is true;
	signal WX1578: std_logic; attribute dont_touch of WX1578: signal is true;
	signal WX1579: std_logic; attribute dont_touch of WX1579: signal is true;
	signal WX1580: std_logic; attribute dont_touch of WX1580: signal is true;
	signal WX1581: std_logic; attribute dont_touch of WX1581: signal is true;
	signal WX1582: std_logic; attribute dont_touch of WX1582: signal is true;
	signal WX1583: std_logic; attribute dont_touch of WX1583: signal is true;
	signal WX1584: std_logic; attribute dont_touch of WX1584: signal is true;
	signal WX1585: std_logic; attribute dont_touch of WX1585: signal is true;
	signal WX1586: std_logic; attribute dont_touch of WX1586: signal is true;
	signal WX1587: std_logic; attribute dont_touch of WX1587: signal is true;
	signal WX1588: std_logic; attribute dont_touch of WX1588: signal is true;
	signal WX1589: std_logic; attribute dont_touch of WX1589: signal is true;
	signal WX1590: std_logic; attribute dont_touch of WX1590: signal is true;
	signal WX1591: std_logic; attribute dont_touch of WX1591: signal is true;
	signal WX1592: std_logic; attribute dont_touch of WX1592: signal is true;
	signal WX1593: std_logic; attribute dont_touch of WX1593: signal is true;
	signal WX1594: std_logic; attribute dont_touch of WX1594: signal is true;
	signal WX1595: std_logic; attribute dont_touch of WX1595: signal is true;
	signal WX1596: std_logic; attribute dont_touch of WX1596: signal is true;
	signal WX1597: std_logic; attribute dont_touch of WX1597: signal is true;
	signal WX1598: std_logic; attribute dont_touch of WX1598: signal is true;
	signal WX1599: std_logic; attribute dont_touch of WX1599: signal is true;
	signal WX1600: std_logic; attribute dont_touch of WX1600: signal is true;
	signal WX1601: std_logic; attribute dont_touch of WX1601: signal is true;
	signal WX1602: std_logic; attribute dont_touch of WX1602: signal is true;
	signal WX1603: std_logic; attribute dont_touch of WX1603: signal is true;
	signal WX1604: std_logic; attribute dont_touch of WX1604: signal is true;
	signal WX1605: std_logic; attribute dont_touch of WX1605: signal is true;
	signal WX1606: std_logic; attribute dont_touch of WX1606: signal is true;
	signal WX1607: std_logic; attribute dont_touch of WX1607: signal is true;
	signal WX1608: std_logic; attribute dont_touch of WX1608: signal is true;
	signal WX1609: std_logic; attribute dont_touch of WX1609: signal is true;
	signal WX1610: std_logic; attribute dont_touch of WX1610: signal is true;
	signal WX1611: std_logic; attribute dont_touch of WX1611: signal is true;
	signal WX1612: std_logic; attribute dont_touch of WX1612: signal is true;
	signal WX1613: std_logic; attribute dont_touch of WX1613: signal is true;
	signal WX1614: std_logic; attribute dont_touch of WX1614: signal is true;
	signal WX1615: std_logic; attribute dont_touch of WX1615: signal is true;
	signal WX1616: std_logic; attribute dont_touch of WX1616: signal is true;
	signal WX1617: std_logic; attribute dont_touch of WX1617: signal is true;
	signal WX1618: std_logic; attribute dont_touch of WX1618: signal is true;
	signal WX1619: std_logic; attribute dont_touch of WX1619: signal is true;
	signal WX1620: std_logic; attribute dont_touch of WX1620: signal is true;
	signal WX1621: std_logic; attribute dont_touch of WX1621: signal is true;
	signal WX1622: std_logic; attribute dont_touch of WX1622: signal is true;
	signal WX1623: std_logic; attribute dont_touch of WX1623: signal is true;
	signal WX1624: std_logic; attribute dont_touch of WX1624: signal is true;
	signal WX1625: std_logic; attribute dont_touch of WX1625: signal is true;
	signal WX1626: std_logic; attribute dont_touch of WX1626: signal is true;
	signal WX1627: std_logic; attribute dont_touch of WX1627: signal is true;
	signal WX1628: std_logic; attribute dont_touch of WX1628: signal is true;
	signal WX1629: std_logic; attribute dont_touch of WX1629: signal is true;
	signal WX1630: std_logic; attribute dont_touch of WX1630: signal is true;
	signal WX1631: std_logic; attribute dont_touch of WX1631: signal is true;
	signal WX1632: std_logic; attribute dont_touch of WX1632: signal is true;
	signal WX1633: std_logic; attribute dont_touch of WX1633: signal is true;
	signal WX1634: std_logic; attribute dont_touch of WX1634: signal is true;
	signal WX1635: std_logic; attribute dont_touch of WX1635: signal is true;
	signal WX1636: std_logic; attribute dont_touch of WX1636: signal is true;
	signal WX1637: std_logic; attribute dont_touch of WX1637: signal is true;
	signal WX1638: std_logic; attribute dont_touch of WX1638: signal is true;
	signal WX1639: std_logic; attribute dont_touch of WX1639: signal is true;
	signal WX1640: std_logic; attribute dont_touch of WX1640: signal is true;
	signal WX1641: std_logic; attribute dont_touch of WX1641: signal is true;
	signal WX1642: std_logic; attribute dont_touch of WX1642: signal is true;
	signal WX1643: std_logic; attribute dont_touch of WX1643: signal is true;
	signal WX1644: std_logic; attribute dont_touch of WX1644: signal is true;
	signal WX1645: std_logic; attribute dont_touch of WX1645: signal is true;
	signal WX1646: std_logic; attribute dont_touch of WX1646: signal is true;
	signal WX1647: std_logic; attribute dont_touch of WX1647: signal is true;
	signal WX1648: std_logic; attribute dont_touch of WX1648: signal is true;
	signal WX1649: std_logic; attribute dont_touch of WX1649: signal is true;
	signal WX1650: std_logic; attribute dont_touch of WX1650: signal is true;
	signal WX1651: std_logic; attribute dont_touch of WX1651: signal is true;
	signal WX1652: std_logic; attribute dont_touch of WX1652: signal is true;
	signal WX1653: std_logic; attribute dont_touch of WX1653: signal is true;
	signal WX1654: std_logic; attribute dont_touch of WX1654: signal is true;
	signal WX1655: std_logic; attribute dont_touch of WX1655: signal is true;
	signal WX1656: std_logic; attribute dont_touch of WX1656: signal is true;
	signal WX1657: std_logic; attribute dont_touch of WX1657: signal is true;
	signal WX1658: std_logic; attribute dont_touch of WX1658: signal is true;
	signal WX1659: std_logic; attribute dont_touch of WX1659: signal is true;
	signal WX1660: std_logic; attribute dont_touch of WX1660: signal is true;
	signal WX1661: std_logic; attribute dont_touch of WX1661: signal is true;
	signal WX1662: std_logic; attribute dont_touch of WX1662: signal is true;
	signal WX1663: std_logic; attribute dont_touch of WX1663: signal is true;
	signal WX1664: std_logic; attribute dont_touch of WX1664: signal is true;
	signal WX1665: std_logic; attribute dont_touch of WX1665: signal is true;
	signal WX1666: std_logic; attribute dont_touch of WX1666: signal is true;
	signal WX1667: std_logic; attribute dont_touch of WX1667: signal is true;
	signal WX1668: std_logic; attribute dont_touch of WX1668: signal is true;
	signal WX1669: std_logic; attribute dont_touch of WX1669: signal is true;
	signal WX1670: std_logic; attribute dont_touch of WX1670: signal is true;
	signal WX1671: std_logic; attribute dont_touch of WX1671: signal is true;
	signal WX1672: std_logic; attribute dont_touch of WX1672: signal is true;
	signal WX1673: std_logic; attribute dont_touch of WX1673: signal is true;
	signal WX1674: std_logic; attribute dont_touch of WX1674: signal is true;
	signal WX1675: std_logic; attribute dont_touch of WX1675: signal is true;
	signal WX1676: std_logic; attribute dont_touch of WX1676: signal is true;
	signal WX1677: std_logic; attribute dont_touch of WX1677: signal is true;
	signal WX1678: std_logic; attribute dont_touch of WX1678: signal is true;
	signal WX1679: std_logic; attribute dont_touch of WX1679: signal is true;
	signal WX1680: std_logic; attribute dont_touch of WX1680: signal is true;
	signal WX1681: std_logic; attribute dont_touch of WX1681: signal is true;
	signal WX1682: std_logic; attribute dont_touch of WX1682: signal is true;
	signal WX1683: std_logic; attribute dont_touch of WX1683: signal is true;
	signal WX1684: std_logic; attribute dont_touch of WX1684: signal is true;
	signal WX1685: std_logic; attribute dont_touch of WX1685: signal is true;
	signal WX1686: std_logic; attribute dont_touch of WX1686: signal is true;
	signal WX1687: std_logic; attribute dont_touch of WX1687: signal is true;
	signal WX1688: std_logic; attribute dont_touch of WX1688: signal is true;
	signal WX1689: std_logic; attribute dont_touch of WX1689: signal is true;
	signal WX1690: std_logic; attribute dont_touch of WX1690: signal is true;
	signal WX1691: std_logic; attribute dont_touch of WX1691: signal is true;
	signal WX1692: std_logic; attribute dont_touch of WX1692: signal is true;
	signal WX1693: std_logic; attribute dont_touch of WX1693: signal is true;
	signal WX1694: std_logic; attribute dont_touch of WX1694: signal is true;
	signal WX1695: std_logic; attribute dont_touch of WX1695: signal is true;
	signal WX1696: std_logic; attribute dont_touch of WX1696: signal is true;
	signal WX1697: std_logic; attribute dont_touch of WX1697: signal is true;
	signal WX1698: std_logic; attribute dont_touch of WX1698: signal is true;
	signal WX1699: std_logic; attribute dont_touch of WX1699: signal is true;
	signal WX1700: std_logic; attribute dont_touch of WX1700: signal is true;
	signal WX1701: std_logic; attribute dont_touch of WX1701: signal is true;
	signal WX1702: std_logic; attribute dont_touch of WX1702: signal is true;
	signal WX1703: std_logic; attribute dont_touch of WX1703: signal is true;
	signal WX1704: std_logic; attribute dont_touch of WX1704: signal is true;
	signal WX1705: std_logic; attribute dont_touch of WX1705: signal is true;
	signal WX1706: std_logic; attribute dont_touch of WX1706: signal is true;
	signal WX1707: std_logic; attribute dont_touch of WX1707: signal is true;
	signal WX1708: std_logic; attribute dont_touch of WX1708: signal is true;
	signal WX1709: std_logic; attribute dont_touch of WX1709: signal is true;
	signal WX1710: std_logic; attribute dont_touch of WX1710: signal is true;
	signal WX1711: std_logic; attribute dont_touch of WX1711: signal is true;
	signal WX1712: std_logic; attribute dont_touch of WX1712: signal is true;
	signal WX1713: std_logic; attribute dont_touch of WX1713: signal is true;
	signal WX1714: std_logic; attribute dont_touch of WX1714: signal is true;
	signal WX1715: std_logic; attribute dont_touch of WX1715: signal is true;
	signal WX1716: std_logic; attribute dont_touch of WX1716: signal is true;
	signal WX1717: std_logic; attribute dont_touch of WX1717: signal is true;
	signal WX1718: std_logic; attribute dont_touch of WX1718: signal is true;
	signal WX1719: std_logic; attribute dont_touch of WX1719: signal is true;
	signal WX1720: std_logic; attribute dont_touch of WX1720: signal is true;
	signal WX1721: std_logic; attribute dont_touch of WX1721: signal is true;
	signal WX1722: std_logic; attribute dont_touch of WX1722: signal is true;
	signal WX1723: std_logic; attribute dont_touch of WX1723: signal is true;
	signal WX1724: std_logic; attribute dont_touch of WX1724: signal is true;
	signal WX1725: std_logic; attribute dont_touch of WX1725: signal is true;
	signal WX1726: std_logic; attribute dont_touch of WX1726: signal is true;
	signal WX1727: std_logic; attribute dont_touch of WX1727: signal is true;
	signal WX1728: std_logic; attribute dont_touch of WX1728: signal is true;
	signal WX1729: std_logic; attribute dont_touch of WX1729: signal is true;
	signal WX1730: std_logic; attribute dont_touch of WX1730: signal is true;
	signal WX1731: std_logic; attribute dont_touch of WX1731: signal is true;
	signal WX1732: std_logic; attribute dont_touch of WX1732: signal is true;
	signal WX1733: std_logic; attribute dont_touch of WX1733: signal is true;
	signal WX1734: std_logic; attribute dont_touch of WX1734: signal is true;
	signal WX1735: std_logic; attribute dont_touch of WX1735: signal is true;
	signal WX1736: std_logic; attribute dont_touch of WX1736: signal is true;
	signal WX1737: std_logic; attribute dont_touch of WX1737: signal is true;
	signal WX1738: std_logic; attribute dont_touch of WX1738: signal is true;
	signal WX1739: std_logic; attribute dont_touch of WX1739: signal is true;
	signal WX1740: std_logic; attribute dont_touch of WX1740: signal is true;
	signal WX1741: std_logic; attribute dont_touch of WX1741: signal is true;
	signal WX1742: std_logic; attribute dont_touch of WX1742: signal is true;
	signal WX1743: std_logic; attribute dont_touch of WX1743: signal is true;
	signal WX1744: std_logic; attribute dont_touch of WX1744: signal is true;
	signal WX1745: std_logic; attribute dont_touch of WX1745: signal is true;
	signal WX1746: std_logic; attribute dont_touch of WX1746: signal is true;
	signal WX1747: std_logic; attribute dont_touch of WX1747: signal is true;
	signal WX1748: std_logic; attribute dont_touch of WX1748: signal is true;
	signal WX1749: std_logic; attribute dont_touch of WX1749: signal is true;
	signal WX1750: std_logic; attribute dont_touch of WX1750: signal is true;
	signal WX1751: std_logic; attribute dont_touch of WX1751: signal is true;
	signal WX1752: std_logic; attribute dont_touch of WX1752: signal is true;
	signal WX1753: std_logic; attribute dont_touch of WX1753: signal is true;
	signal WX1754: std_logic; attribute dont_touch of WX1754: signal is true;
	signal WX1755: std_logic; attribute dont_touch of WX1755: signal is true;
	signal WX1756: std_logic; attribute dont_touch of WX1756: signal is true;
	signal WX1757: std_logic; attribute dont_touch of WX1757: signal is true;
	signal WX1758: std_logic; attribute dont_touch of WX1758: signal is true;
	signal WX1759: std_logic; attribute dont_touch of WX1759: signal is true;
	signal WX1760: std_logic; attribute dont_touch of WX1760: signal is true;
	signal WX1761: std_logic; attribute dont_touch of WX1761: signal is true;
	signal WX1762: std_logic; attribute dont_touch of WX1762: signal is true;
	signal WX1763: std_logic; attribute dont_touch of WX1763: signal is true;
	signal WX1764: std_logic; attribute dont_touch of WX1764: signal is true;
	signal WX1765: std_logic; attribute dont_touch of WX1765: signal is true;
	signal WX1766: std_logic; attribute dont_touch of WX1766: signal is true;
	signal WX1767: std_logic; attribute dont_touch of WX1767: signal is true;
	signal WX1768: std_logic; attribute dont_touch of WX1768: signal is true;
	signal WX1769: std_logic; attribute dont_touch of WX1769: signal is true;
	signal WX1770: std_logic; attribute dont_touch of WX1770: signal is true;
	signal WX1771: std_logic; attribute dont_touch of WX1771: signal is true;
	signal WX1772: std_logic; attribute dont_touch of WX1772: signal is true;
	signal WX1773: std_logic; attribute dont_touch of WX1773: signal is true;
	signal WX1774: std_logic; attribute dont_touch of WX1774: signal is true;
	signal WX1775: std_logic; attribute dont_touch of WX1775: signal is true;
	signal WX1776: std_logic; attribute dont_touch of WX1776: signal is true;
	signal WX1777: std_logic; attribute dont_touch of WX1777: signal is true;
	signal WX1778: std_logic; attribute dont_touch of WX1778: signal is true;
	signal WX1779: std_logic; attribute dont_touch of WX1779: signal is true;
	signal WX1780: std_logic; attribute dont_touch of WX1780: signal is true;
	signal WX1781: std_logic; attribute dont_touch of WX1781: signal is true;
	signal WX1782: std_logic; attribute dont_touch of WX1782: signal is true;
	signal WX1783: std_logic; attribute dont_touch of WX1783: signal is true;
	signal WX1784: std_logic; attribute dont_touch of WX1784: signal is true;
	signal WX1785: std_logic; attribute dont_touch of WX1785: signal is true;
	signal WX1786: std_logic; attribute dont_touch of WX1786: signal is true;
	signal WX1787: std_logic; attribute dont_touch of WX1787: signal is true;
	signal WX1788: std_logic; attribute dont_touch of WX1788: signal is true;
	signal WX1789: std_logic; attribute dont_touch of WX1789: signal is true;
	signal WX1790: std_logic; attribute dont_touch of WX1790: signal is true;
	signal WX1791: std_logic; attribute dont_touch of WX1791: signal is true;
	signal WX1792: std_logic; attribute dont_touch of WX1792: signal is true;
	signal WX1793: std_logic; attribute dont_touch of WX1793: signal is true;
	signal WX1794: std_logic; attribute dont_touch of WX1794: signal is true;
	signal WX1795: std_logic; attribute dont_touch of WX1795: signal is true;
	signal WX1796: std_logic; attribute dont_touch of WX1796: signal is true;
	signal WX1797: std_logic; attribute dont_touch of WX1797: signal is true;
	signal WX1798: std_logic; attribute dont_touch of WX1798: signal is true;
	signal WX1799: std_logic; attribute dont_touch of WX1799: signal is true;
	signal WX1800: std_logic; attribute dont_touch of WX1800: signal is true;
	signal WX1801: std_logic; attribute dont_touch of WX1801: signal is true;
	signal WX1802: std_logic; attribute dont_touch of WX1802: signal is true;
	signal WX1803: std_logic; attribute dont_touch of WX1803: signal is true;
	signal WX1804: std_logic; attribute dont_touch of WX1804: signal is true;
	signal WX1805: std_logic; attribute dont_touch of WX1805: signal is true;
	signal WX1806: std_logic; attribute dont_touch of WX1806: signal is true;
	signal WX1807: std_logic; attribute dont_touch of WX1807: signal is true;
	signal WX1808: std_logic; attribute dont_touch of WX1808: signal is true;
	signal WX1809: std_logic; attribute dont_touch of WX1809: signal is true;
	signal WX1810: std_logic; attribute dont_touch of WX1810: signal is true;
	signal WX1811: std_logic; attribute dont_touch of WX1811: signal is true;
	signal WX1812: std_logic; attribute dont_touch of WX1812: signal is true;
	signal WX1813: std_logic; attribute dont_touch of WX1813: signal is true;
	signal WX1814: std_logic; attribute dont_touch of WX1814: signal is true;
	signal WX1815: std_logic; attribute dont_touch of WX1815: signal is true;
	signal WX1816: std_logic; attribute dont_touch of WX1816: signal is true;
	signal WX1817: std_logic; attribute dont_touch of WX1817: signal is true;
	signal WX1818: std_logic; attribute dont_touch of WX1818: signal is true;
	signal WX1819: std_logic; attribute dont_touch of WX1819: signal is true;
	signal WX1820: std_logic; attribute dont_touch of WX1820: signal is true;
	signal WX1821: std_logic; attribute dont_touch of WX1821: signal is true;
	signal WX1822: std_logic; attribute dont_touch of WX1822: signal is true;
	signal WX1823: std_logic; attribute dont_touch of WX1823: signal is true;
	signal WX1824: std_logic; attribute dont_touch of WX1824: signal is true;
	signal WX1825: std_logic; attribute dont_touch of WX1825: signal is true;
	signal WX1826: std_logic; attribute dont_touch of WX1826: signal is true;
	signal WX1827: std_logic; attribute dont_touch of WX1827: signal is true;
	signal WX1828: std_logic; attribute dont_touch of WX1828: signal is true;
	signal WX1829: std_logic; attribute dont_touch of WX1829: signal is true;
	signal WX1830: std_logic; attribute dont_touch of WX1830: signal is true;
	signal WX1831: std_logic; attribute dont_touch of WX1831: signal is true;
	signal WX1832: std_logic; attribute dont_touch of WX1832: signal is true;
	signal WX1833: std_logic; attribute dont_touch of WX1833: signal is true;
	signal WX1834: std_logic; attribute dont_touch of WX1834: signal is true;
	signal WX1835: std_logic; attribute dont_touch of WX1835: signal is true;
	signal WX1836: std_logic; attribute dont_touch of WX1836: signal is true;
	signal WX1837: std_logic; attribute dont_touch of WX1837: signal is true;
	signal WX1838: std_logic; attribute dont_touch of WX1838: signal is true;
	signal WX1839: std_logic; attribute dont_touch of WX1839: signal is true;
	signal WX1840: std_logic; attribute dont_touch of WX1840: signal is true;
	signal WX1841: std_logic; attribute dont_touch of WX1841: signal is true;
	signal WX1842: std_logic; attribute dont_touch of WX1842: signal is true;
	signal WX1843: std_logic; attribute dont_touch of WX1843: signal is true;
	signal WX1844: std_logic; attribute dont_touch of WX1844: signal is true;
	signal WX1845: std_logic; attribute dont_touch of WX1845: signal is true;
	signal WX1846: std_logic; attribute dont_touch of WX1846: signal is true;
	signal WX1847: std_logic; attribute dont_touch of WX1847: signal is true;
	signal WX1848: std_logic; attribute dont_touch of WX1848: signal is true;
	signal WX1849: std_logic; attribute dont_touch of WX1849: signal is true;
	signal WX1850: std_logic; attribute dont_touch of WX1850: signal is true;
	signal WX1851: std_logic; attribute dont_touch of WX1851: signal is true;
	signal WX1852: std_logic; attribute dont_touch of WX1852: signal is true;
	signal WX1853: std_logic; attribute dont_touch of WX1853: signal is true;
	signal WX1854: std_logic; attribute dont_touch of WX1854: signal is true;
	signal WX1855: std_logic; attribute dont_touch of WX1855: signal is true;
	signal WX1856: std_logic; attribute dont_touch of WX1856: signal is true;
	signal WX1857: std_logic; attribute dont_touch of WX1857: signal is true;
	signal WX1858: std_logic; attribute dont_touch of WX1858: signal is true;
	signal WX1859: std_logic; attribute dont_touch of WX1859: signal is true;
	signal WX1860: std_logic; attribute dont_touch of WX1860: signal is true;
	signal WX1861: std_logic; attribute dont_touch of WX1861: signal is true;
	signal WX1862: std_logic; attribute dont_touch of WX1862: signal is true;
	signal WX1863: std_logic; attribute dont_touch of WX1863: signal is true;
	signal WX1864: std_logic; attribute dont_touch of WX1864: signal is true;
	signal WX1865: std_logic; attribute dont_touch of WX1865: signal is true;
	signal WX1866: std_logic; attribute dont_touch of WX1866: signal is true;
	signal WX1867: std_logic; attribute dont_touch of WX1867: signal is true;
	signal WX1868: std_logic; attribute dont_touch of WX1868: signal is true;
	signal WX1869: std_logic; attribute dont_touch of WX1869: signal is true;
	signal WX1870: std_logic; attribute dont_touch of WX1870: signal is true;
	signal WX1871: std_logic; attribute dont_touch of WX1871: signal is true;
	signal WX1872: std_logic; attribute dont_touch of WX1872: signal is true;
	signal WX1873: std_logic; attribute dont_touch of WX1873: signal is true;
	signal WX1874: std_logic; attribute dont_touch of WX1874: signal is true;
	signal WX1875: std_logic; attribute dont_touch of WX1875: signal is true;
	signal WX1876: std_logic; attribute dont_touch of WX1876: signal is true;
	signal WX1877: std_logic; attribute dont_touch of WX1877: signal is true;
	signal WX1878: std_logic; attribute dont_touch of WX1878: signal is true;
	signal WX1879: std_logic; attribute dont_touch of WX1879: signal is true;
	signal WX1880: std_logic; attribute dont_touch of WX1880: signal is true;
	signal WX1881: std_logic; attribute dont_touch of WX1881: signal is true;
	signal WX1882: std_logic; attribute dont_touch of WX1882: signal is true;
	signal WX1883: std_logic; attribute dont_touch of WX1883: signal is true;
	signal WX1884: std_logic; attribute dont_touch of WX1884: signal is true;
	signal WX1885: std_logic; attribute dont_touch of WX1885: signal is true;
	signal WX1886: std_logic; attribute dont_touch of WX1886: signal is true;
	signal WX1887: std_logic; attribute dont_touch of WX1887: signal is true;
	signal WX1888: std_logic; attribute dont_touch of WX1888: signal is true;
	signal WX1889: std_logic; attribute dont_touch of WX1889: signal is true;
	signal WX1890: std_logic; attribute dont_touch of WX1890: signal is true;
	signal WX1891: std_logic; attribute dont_touch of WX1891: signal is true;
	signal WX1892: std_logic; attribute dont_touch of WX1892: signal is true;
	signal WX1893: std_logic; attribute dont_touch of WX1893: signal is true;
	signal WX1894: std_logic; attribute dont_touch of WX1894: signal is true;
	signal WX1895: std_logic; attribute dont_touch of WX1895: signal is true;
	signal WX1896: std_logic; attribute dont_touch of WX1896: signal is true;
	signal WX1897: std_logic; attribute dont_touch of WX1897: signal is true;
	signal WX1898: std_logic; attribute dont_touch of WX1898: signal is true;
	signal WX1899: std_logic; attribute dont_touch of WX1899: signal is true;
	signal WX1900: std_logic; attribute dont_touch of WX1900: signal is true;
	signal WX1901: std_logic; attribute dont_touch of WX1901: signal is true;
	signal WX1902: std_logic; attribute dont_touch of WX1902: signal is true;
	signal WX1903: std_logic; attribute dont_touch of WX1903: signal is true;
	signal WX1904: std_logic; attribute dont_touch of WX1904: signal is true;
	signal WX1905: std_logic; attribute dont_touch of WX1905: signal is true;
	signal WX1906: std_logic; attribute dont_touch of WX1906: signal is true;
	signal WX1907: std_logic; attribute dont_touch of WX1907: signal is true;
	signal WX1908: std_logic; attribute dont_touch of WX1908: signal is true;
	signal WX1909: std_logic; attribute dont_touch of WX1909: signal is true;
	signal WX1910: std_logic; attribute dont_touch of WX1910: signal is true;
	signal WX1911: std_logic; attribute dont_touch of WX1911: signal is true;
	signal WX1912: std_logic; attribute dont_touch of WX1912: signal is true;
	signal WX1913: std_logic; attribute dont_touch of WX1913: signal is true;
	signal WX1914: std_logic; attribute dont_touch of WX1914: signal is true;
	signal WX1915: std_logic; attribute dont_touch of WX1915: signal is true;
	signal WX1916: std_logic; attribute dont_touch of WX1916: signal is true;
	signal WX1917: std_logic; attribute dont_touch of WX1917: signal is true;
	signal WX1918: std_logic; attribute dont_touch of WX1918: signal is true;
	signal WX1919: std_logic; attribute dont_touch of WX1919: signal is true;
	signal WX1920: std_logic; attribute dont_touch of WX1920: signal is true;
	signal WX1921: std_logic; attribute dont_touch of WX1921: signal is true;
	signal WX1922: std_logic; attribute dont_touch of WX1922: signal is true;
	signal WX1923: std_logic; attribute dont_touch of WX1923: signal is true;
	signal WX1924: std_logic; attribute dont_touch of WX1924: signal is true;
	signal WX1925: std_logic; attribute dont_touch of WX1925: signal is true;
	signal WX1926: std_logic; attribute dont_touch of WX1926: signal is true;
	signal WX1927: std_logic; attribute dont_touch of WX1927: signal is true;
	signal WX1928: std_logic; attribute dont_touch of WX1928: signal is true;
	signal WX1929: std_logic; attribute dont_touch of WX1929: signal is true;
	signal WX1930: std_logic; attribute dont_touch of WX1930: signal is true;
	signal WX1931: std_logic; attribute dont_touch of WX1931: signal is true;
	signal WX1932: std_logic; attribute dont_touch of WX1932: signal is true;
	signal WX1933: std_logic; attribute dont_touch of WX1933: signal is true;
	signal WX1934: std_logic; attribute dont_touch of WX1934: signal is true;
	signal WX1935: std_logic; attribute dont_touch of WX1935: signal is true;
	signal WX1936: std_logic; attribute dont_touch of WX1936: signal is true;
	signal WX1937: std_logic; attribute dont_touch of WX1937: signal is true;
	signal WX1938: std_logic; attribute dont_touch of WX1938: signal is true;
	signal WX1939: std_logic; attribute dont_touch of WX1939: signal is true;
	signal WX1940: std_logic; attribute dont_touch of WX1940: signal is true;
	signal WX1941: std_logic; attribute dont_touch of WX1941: signal is true;
	signal WX1942: std_logic; attribute dont_touch of WX1942: signal is true;
	signal WX1943: std_logic; attribute dont_touch of WX1943: signal is true;
	signal WX1944: std_logic; attribute dont_touch of WX1944: signal is true;
	signal WX1945: std_logic; attribute dont_touch of WX1945: signal is true;
	signal WX1946: std_logic; attribute dont_touch of WX1946: signal is true;
	signal WX1947: std_logic; attribute dont_touch of WX1947: signal is true;
	signal WX1948: std_logic; attribute dont_touch of WX1948: signal is true;
	signal WX1949: std_logic; attribute dont_touch of WX1949: signal is true;
	signal WX1950: std_logic; attribute dont_touch of WX1950: signal is true;
	signal WX1951: std_logic; attribute dont_touch of WX1951: signal is true;
	signal WX1952: std_logic; attribute dont_touch of WX1952: signal is true;
	signal WX1953: std_logic; attribute dont_touch of WX1953: signal is true;
	signal WX1954: std_logic; attribute dont_touch of WX1954: signal is true;
	signal WX1955: std_logic; attribute dont_touch of WX1955: signal is true;
	signal WX1956: std_logic; attribute dont_touch of WX1956: signal is true;
	signal WX1957: std_logic; attribute dont_touch of WX1957: signal is true;
	signal WX1958: std_logic; attribute dont_touch of WX1958: signal is true;
	signal WX1959: std_logic; attribute dont_touch of WX1959: signal is true;
	signal WX1960: std_logic; attribute dont_touch of WX1960: signal is true;
	signal WX1961: std_logic; attribute dont_touch of WX1961: signal is true;
	signal WX1962: std_logic; attribute dont_touch of WX1962: signal is true;
	signal WX1963: std_logic; attribute dont_touch of WX1963: signal is true;
	signal WX1964: std_logic; attribute dont_touch of WX1964: signal is true;
	signal WX1965: std_logic; attribute dont_touch of WX1965: signal is true;
	signal WX1966: std_logic; attribute dont_touch of WX1966: signal is true;
	signal WX1967: std_logic; attribute dont_touch of WX1967: signal is true;
	signal WX1968: std_logic; attribute dont_touch of WX1968: signal is true;
	signal WX1969: std_logic; attribute dont_touch of WX1969: signal is true;
	signal WX1970: std_logic; attribute dont_touch of WX1970: signal is true;
	signal WX1971: std_logic; attribute dont_touch of WX1971: signal is true;
	signal WX1972: std_logic; attribute dont_touch of WX1972: signal is true;
	signal WX1973: std_logic; attribute dont_touch of WX1973: signal is true;
	signal WX1974: std_logic; attribute dont_touch of WX1974: signal is true;
	signal WX1975: std_logic; attribute dont_touch of WX1975: signal is true;
	signal WX1976: std_logic; attribute dont_touch of WX1976: signal is true;
	signal WX1977: std_logic; attribute dont_touch of WX1977: signal is true;
	signal WX1978: std_logic; attribute dont_touch of WX1978: signal is true;
	signal WX1979: std_logic; attribute dont_touch of WX1979: signal is true;
	signal WX1980: std_logic; attribute dont_touch of WX1980: signal is true;
	signal WX1981: std_logic; attribute dont_touch of WX1981: signal is true;
	signal WX1982: std_logic; attribute dont_touch of WX1982: signal is true;
	signal WX1983: std_logic; attribute dont_touch of WX1983: signal is true;
	signal WX1984: std_logic; attribute dont_touch of WX1984: signal is true;
	signal WX1985: std_logic; attribute dont_touch of WX1985: signal is true;
	signal WX1986: std_logic; attribute dont_touch of WX1986: signal is true;
	signal WX1987: std_logic; attribute dont_touch of WX1987: signal is true;
	signal WX1988: std_logic; attribute dont_touch of WX1988: signal is true;
	signal WX1989: std_logic; attribute dont_touch of WX1989: signal is true;
	signal WX1990: std_logic; attribute dont_touch of WX1990: signal is true;
	signal WX1991: std_logic; attribute dont_touch of WX1991: signal is true;
	signal WX1992: std_logic; attribute dont_touch of WX1992: signal is true;
	signal WX1993: std_logic; attribute dont_touch of WX1993: signal is true;
	signal WX1994: std_logic; attribute dont_touch of WX1994: signal is true;
	signal WX1995: std_logic; attribute dont_touch of WX1995: signal is true;
	signal WX1996: std_logic; attribute dont_touch of WX1996: signal is true;
	signal WX1997: std_logic; attribute dont_touch of WX1997: signal is true;
	signal WX1998: std_logic; attribute dont_touch of WX1998: signal is true;
	signal WX1999: std_logic; attribute dont_touch of WX1999: signal is true;
	signal WX2000: std_logic; attribute dont_touch of WX2000: signal is true;
	signal WX2001: std_logic; attribute dont_touch of WX2001: signal is true;
	signal WX2002: std_logic; attribute dont_touch of WX2002: signal is true;
	signal WX2003: std_logic; attribute dont_touch of WX2003: signal is true;
	signal WX2004: std_logic; attribute dont_touch of WX2004: signal is true;
	signal WX2005: std_logic; attribute dont_touch of WX2005: signal is true;
	signal WX2006: std_logic; attribute dont_touch of WX2006: signal is true;
	signal WX2007: std_logic; attribute dont_touch of WX2007: signal is true;
	signal WX2008: std_logic; attribute dont_touch of WX2008: signal is true;
	signal WX2009: std_logic; attribute dont_touch of WX2009: signal is true;
	signal WX2010: std_logic; attribute dont_touch of WX2010: signal is true;
	signal WX2011: std_logic; attribute dont_touch of WX2011: signal is true;
	signal WX2012: std_logic; attribute dont_touch of WX2012: signal is true;
	signal WX2013: std_logic; attribute dont_touch of WX2013: signal is true;
	signal WX2014: std_logic; attribute dont_touch of WX2014: signal is true;
	signal WX2015: std_logic; attribute dont_touch of WX2015: signal is true;
	signal WX2016: std_logic; attribute dont_touch of WX2016: signal is true;
	signal WX2017: std_logic; attribute dont_touch of WX2017: signal is true;
	signal WX2018: std_logic; attribute dont_touch of WX2018: signal is true;
	signal WX2019: std_logic; attribute dont_touch of WX2019: signal is true;
	signal WX2020: std_logic; attribute dont_touch of WX2020: signal is true;
	signal WX2021: std_logic; attribute dont_touch of WX2021: signal is true;
	signal WX2022: std_logic; attribute dont_touch of WX2022: signal is true;
	signal WX2023: std_logic; attribute dont_touch of WX2023: signal is true;
	signal WX2024: std_logic; attribute dont_touch of WX2024: signal is true;
	signal WX2025: std_logic; attribute dont_touch of WX2025: signal is true;
	signal WX2026: std_logic; attribute dont_touch of WX2026: signal is true;
	signal WX2027: std_logic; attribute dont_touch of WX2027: signal is true;
	signal WX2028: std_logic; attribute dont_touch of WX2028: signal is true;
	signal WX2029: std_logic; attribute dont_touch of WX2029: signal is true;
	signal WX2030: std_logic; attribute dont_touch of WX2030: signal is true;
	signal WX2031: std_logic; attribute dont_touch of WX2031: signal is true;
	signal WX2032: std_logic; attribute dont_touch of WX2032: signal is true;
	signal WX2033: std_logic; attribute dont_touch of WX2033: signal is true;
	signal WX2034: std_logic; attribute dont_touch of WX2034: signal is true;
	signal WX2035: std_logic; attribute dont_touch of WX2035: signal is true;
	signal WX2036: std_logic; attribute dont_touch of WX2036: signal is true;
	signal WX2037: std_logic; attribute dont_touch of WX2037: signal is true;
	signal WX2038: std_logic; attribute dont_touch of WX2038: signal is true;
	signal WX2039: std_logic; attribute dont_touch of WX2039: signal is true;
	signal WX2040: std_logic; attribute dont_touch of WX2040: signal is true;
	signal WX2041: std_logic; attribute dont_touch of WX2041: signal is true;
	signal WX2042: std_logic; attribute dont_touch of WX2042: signal is true;
	signal WX2043: std_logic; attribute dont_touch of WX2043: signal is true;
	signal WX2044: std_logic; attribute dont_touch of WX2044: signal is true;
	signal WX2045: std_logic; attribute dont_touch of WX2045: signal is true;
	signal WX2046: std_logic; attribute dont_touch of WX2046: signal is true;
	signal WX2047: std_logic; attribute dont_touch of WX2047: signal is true;
	signal WX2048: std_logic; attribute dont_touch of WX2048: signal is true;
	signal WX2049: std_logic; attribute dont_touch of WX2049: signal is true;
	signal WX2050: std_logic; attribute dont_touch of WX2050: signal is true;
	signal WX2051: std_logic; attribute dont_touch of WX2051: signal is true;
	signal WX2052: std_logic; attribute dont_touch of WX2052: signal is true;
	signal WX2053: std_logic; attribute dont_touch of WX2053: signal is true;
	signal WX2054: std_logic; attribute dont_touch of WX2054: signal is true;
	signal WX2055: std_logic; attribute dont_touch of WX2055: signal is true;
	signal WX2056: std_logic; attribute dont_touch of WX2056: signal is true;
	signal WX2057: std_logic; attribute dont_touch of WX2057: signal is true;
	signal WX2058: std_logic; attribute dont_touch of WX2058: signal is true;
	signal WX2059: std_logic; attribute dont_touch of WX2059: signal is true;
	signal WX2060: std_logic; attribute dont_touch of WX2060: signal is true;
	signal WX2061: std_logic; attribute dont_touch of WX2061: signal is true;
	signal WX2062: std_logic; attribute dont_touch of WX2062: signal is true;
	signal WX2063: std_logic; attribute dont_touch of WX2063: signal is true;
	signal WX2064: std_logic; attribute dont_touch of WX2064: signal is true;
	signal WX2065: std_logic; attribute dont_touch of WX2065: signal is true;
	signal WX2066: std_logic; attribute dont_touch of WX2066: signal is true;
	signal WX2067: std_logic; attribute dont_touch of WX2067: signal is true;
	signal WX2068: std_logic; attribute dont_touch of WX2068: signal is true;
	signal WX2069: std_logic; attribute dont_touch of WX2069: signal is true;
	signal WX2070: std_logic; attribute dont_touch of WX2070: signal is true;
	signal WX2071: std_logic; attribute dont_touch of WX2071: signal is true;
	signal WX2072: std_logic; attribute dont_touch of WX2072: signal is true;
	signal WX2073: std_logic; attribute dont_touch of WX2073: signal is true;
	signal WX2074: std_logic; attribute dont_touch of WX2074: signal is true;
	signal WX2075: std_logic; attribute dont_touch of WX2075: signal is true;
	signal WX2076: std_logic; attribute dont_touch of WX2076: signal is true;
	signal WX2077: std_logic; attribute dont_touch of WX2077: signal is true;
	signal WX2078: std_logic; attribute dont_touch of WX2078: signal is true;
	signal WX2079: std_logic; attribute dont_touch of WX2079: signal is true;
	signal WX2080: std_logic; attribute dont_touch of WX2080: signal is true;
	signal WX2081: std_logic; attribute dont_touch of WX2081: signal is true;
	signal WX2082: std_logic; attribute dont_touch of WX2082: signal is true;
	signal WX2083: std_logic; attribute dont_touch of WX2083: signal is true;
	signal WX2084: std_logic; attribute dont_touch of WX2084: signal is true;
	signal WX2085: std_logic; attribute dont_touch of WX2085: signal is true;
	signal WX2086: std_logic; attribute dont_touch of WX2086: signal is true;
	signal WX2087: std_logic; attribute dont_touch of WX2087: signal is true;
	signal WX2088: std_logic; attribute dont_touch of WX2088: signal is true;
	signal WX2089: std_logic; attribute dont_touch of WX2089: signal is true;
	signal WX2090: std_logic; attribute dont_touch of WX2090: signal is true;
	signal WX2091: std_logic; attribute dont_touch of WX2091: signal is true;
	signal WX2092: std_logic; attribute dont_touch of WX2092: signal is true;
	signal WX2093: std_logic; attribute dont_touch of WX2093: signal is true;
	signal WX2094: std_logic; attribute dont_touch of WX2094: signal is true;
	signal WX2095: std_logic; attribute dont_touch of WX2095: signal is true;
	signal WX2096: std_logic; attribute dont_touch of WX2096: signal is true;
	signal WX2097: std_logic; attribute dont_touch of WX2097: signal is true;
	signal WX2098: std_logic; attribute dont_touch of WX2098: signal is true;
	signal WX2099: std_logic; attribute dont_touch of WX2099: signal is true;
	signal WX2100: std_logic; attribute dont_touch of WX2100: signal is true;
	signal WX2101: std_logic; attribute dont_touch of WX2101: signal is true;
	signal WX2102: std_logic; attribute dont_touch of WX2102: signal is true;
	signal WX2103: std_logic; attribute dont_touch of WX2103: signal is true;
	signal WX2104: std_logic; attribute dont_touch of WX2104: signal is true;
	signal WX2105: std_logic; attribute dont_touch of WX2105: signal is true;
	signal WX2106: std_logic; attribute dont_touch of WX2106: signal is true;
	signal WX2107: std_logic; attribute dont_touch of WX2107: signal is true;
	signal WX2108: std_logic; attribute dont_touch of WX2108: signal is true;
	signal WX2109: std_logic; attribute dont_touch of WX2109: signal is true;
	signal WX2110: std_logic; attribute dont_touch of WX2110: signal is true;
	signal WX2111: std_logic; attribute dont_touch of WX2111: signal is true;
	signal WX2112: std_logic; attribute dont_touch of WX2112: signal is true;
	signal WX2113: std_logic; attribute dont_touch of WX2113: signal is true;
	signal WX2114: std_logic; attribute dont_touch of WX2114: signal is true;
	signal WX2115: std_logic; attribute dont_touch of WX2115: signal is true;
	signal WX2116: std_logic; attribute dont_touch of WX2116: signal is true;
	signal WX2117: std_logic; attribute dont_touch of WX2117: signal is true;
	signal WX2118: std_logic; attribute dont_touch of WX2118: signal is true;
	signal WX2119: std_logic; attribute dont_touch of WX2119: signal is true;
	signal WX2120: std_logic; attribute dont_touch of WX2120: signal is true;
	signal WX2121: std_logic; attribute dont_touch of WX2121: signal is true;
	signal WX2122: std_logic; attribute dont_touch of WX2122: signal is true;
	signal WX2123: std_logic; attribute dont_touch of WX2123: signal is true;
	signal WX2124: std_logic; attribute dont_touch of WX2124: signal is true;
	signal WX2125: std_logic; attribute dont_touch of WX2125: signal is true;
	signal WX2126: std_logic; attribute dont_touch of WX2126: signal is true;
	signal WX2127: std_logic; attribute dont_touch of WX2127: signal is true;
	signal WX2128: std_logic; attribute dont_touch of WX2128: signal is true;
	signal WX2129: std_logic; attribute dont_touch of WX2129: signal is true;
	signal WX2130: std_logic; attribute dont_touch of WX2130: signal is true;
	signal WX2131: std_logic; attribute dont_touch of WX2131: signal is true;
	signal WX2132: std_logic; attribute dont_touch of WX2132: signal is true;
	signal WX2133: std_logic; attribute dont_touch of WX2133: signal is true;
	signal WX2134: std_logic; attribute dont_touch of WX2134: signal is true;
	signal WX2135: std_logic; attribute dont_touch of WX2135: signal is true;
	signal WX2136: std_logic; attribute dont_touch of WX2136: signal is true;
	signal WX2137: std_logic; attribute dont_touch of WX2137: signal is true;
	signal WX2138: std_logic; attribute dont_touch of WX2138: signal is true;
	signal WX2139: std_logic; attribute dont_touch of WX2139: signal is true;
	signal WX2140: std_logic; attribute dont_touch of WX2140: signal is true;
	signal WX2141: std_logic; attribute dont_touch of WX2141: signal is true;
	signal WX2142: std_logic; attribute dont_touch of WX2142: signal is true;
	signal WX2143: std_logic; attribute dont_touch of WX2143: signal is true;
	signal WX2144: std_logic; attribute dont_touch of WX2144: signal is true;
	signal WX2145: std_logic; attribute dont_touch of WX2145: signal is true;
	signal WX2146: std_logic; attribute dont_touch of WX2146: signal is true;
	signal WX2147: std_logic; attribute dont_touch of WX2147: signal is true;
	signal WX2148: std_logic; attribute dont_touch of WX2148: signal is true;
	signal WX2149: std_logic; attribute dont_touch of WX2149: signal is true;
	signal WX2150: std_logic; attribute dont_touch of WX2150: signal is true;
	signal WX2151: std_logic; attribute dont_touch of WX2151: signal is true;
	signal WX2152: std_logic; attribute dont_touch of WX2152: signal is true;
	signal WX2153: std_logic; attribute dont_touch of WX2153: signal is true;
	signal WX2154: std_logic; attribute dont_touch of WX2154: signal is true;
	signal WX2155: std_logic; attribute dont_touch of WX2155: signal is true;
	signal WX2156: std_logic; attribute dont_touch of WX2156: signal is true;
	signal WX2157: std_logic; attribute dont_touch of WX2157: signal is true;
	signal WX2158: std_logic; attribute dont_touch of WX2158: signal is true;
	signal WX2159: std_logic; attribute dont_touch of WX2159: signal is true;
	signal WX2160: std_logic; attribute dont_touch of WX2160: signal is true;
	signal WX2161: std_logic; attribute dont_touch of WX2161: signal is true;
	signal WX2162: std_logic; attribute dont_touch of WX2162: signal is true;
	signal WX2163: std_logic; attribute dont_touch of WX2163: signal is true;
	signal WX2164: std_logic; attribute dont_touch of WX2164: signal is true;
	signal WX2165: std_logic; attribute dont_touch of WX2165: signal is true;
	signal WX2166: std_logic; attribute dont_touch of WX2166: signal is true;
	signal WX2167: std_logic; attribute dont_touch of WX2167: signal is true;
	signal WX2168: std_logic; attribute dont_touch of WX2168: signal is true;
	signal WX2169: std_logic; attribute dont_touch of WX2169: signal is true;
	signal WX2170: std_logic; attribute dont_touch of WX2170: signal is true;
	signal WX2171: std_logic; attribute dont_touch of WX2171: signal is true;
	signal WX2172: std_logic; attribute dont_touch of WX2172: signal is true;
	signal WX2173: std_logic; attribute dont_touch of WX2173: signal is true;
	signal WX2174: std_logic; attribute dont_touch of WX2174: signal is true;
	signal WX2175: std_logic; attribute dont_touch of WX2175: signal is true;
	signal WX2176: std_logic; attribute dont_touch of WX2176: signal is true;
	signal WX2177: std_logic; attribute dont_touch of WX2177: signal is true;
	signal WX2178: std_logic; attribute dont_touch of WX2178: signal is true;
	signal WX2179: std_logic; attribute dont_touch of WX2179: signal is true;
	signal WX2180: std_logic; attribute dont_touch of WX2180: signal is true;
	signal WX2181: std_logic; attribute dont_touch of WX2181: signal is true;
	signal WX2182: std_logic; attribute dont_touch of WX2182: signal is true;
	signal WX2183: std_logic; attribute dont_touch of WX2183: signal is true;
	signal WX2184: std_logic; attribute dont_touch of WX2184: signal is true;
	signal WX2185: std_logic; attribute dont_touch of WX2185: signal is true;
	signal WX2186: std_logic; attribute dont_touch of WX2186: signal is true;
	signal WX2187: std_logic; attribute dont_touch of WX2187: signal is true;
	signal WX2188: std_logic; attribute dont_touch of WX2188: signal is true;
	signal WX2189: std_logic; attribute dont_touch of WX2189: signal is true;
	signal WX2190: std_logic; attribute dont_touch of WX2190: signal is true;
	signal WX2191: std_logic; attribute dont_touch of WX2191: signal is true;
	signal WX2192: std_logic; attribute dont_touch of WX2192: signal is true;
	signal WX2193: std_logic; attribute dont_touch of WX2193: signal is true;
	signal WX2194: std_logic; attribute dont_touch of WX2194: signal is true;
	signal WX2195: std_logic; attribute dont_touch of WX2195: signal is true;
	signal WX2196: std_logic; attribute dont_touch of WX2196: signal is true;
	signal WX2197: std_logic; attribute dont_touch of WX2197: signal is true;
	signal WX2198: std_logic; attribute dont_touch of WX2198: signal is true;
	signal WX2199: std_logic; attribute dont_touch of WX2199: signal is true;
	signal WX2200: std_logic; attribute dont_touch of WX2200: signal is true;
	signal WX2201: std_logic; attribute dont_touch of WX2201: signal is true;
	signal WX2202: std_logic; attribute dont_touch of WX2202: signal is true;
	signal WX2203: std_logic; attribute dont_touch of WX2203: signal is true;
	signal WX2204: std_logic; attribute dont_touch of WX2204: signal is true;
	signal WX2205: std_logic; attribute dont_touch of WX2205: signal is true;
	signal WX2206: std_logic; attribute dont_touch of WX2206: signal is true;
	signal WX2207: std_logic; attribute dont_touch of WX2207: signal is true;
	signal WX2208: std_logic; attribute dont_touch of WX2208: signal is true;
	signal WX2209: std_logic; attribute dont_touch of WX2209: signal is true;
	signal WX2210: std_logic; attribute dont_touch of WX2210: signal is true;
	signal WX2211: std_logic; attribute dont_touch of WX2211: signal is true;
	signal WX2212: std_logic; attribute dont_touch of WX2212: signal is true;
	signal WX2213: std_logic; attribute dont_touch of WX2213: signal is true;
	signal WX2214: std_logic; attribute dont_touch of WX2214: signal is true;
	signal WX2215: std_logic; attribute dont_touch of WX2215: signal is true;
	signal WX2216: std_logic; attribute dont_touch of WX2216: signal is true;
	signal WX2217: std_logic; attribute dont_touch of WX2217: signal is true;
	signal WX2218: std_logic; attribute dont_touch of WX2218: signal is true;
	signal WX2219: std_logic; attribute dont_touch of WX2219: signal is true;
	signal WX2220: std_logic; attribute dont_touch of WX2220: signal is true;
	signal WX2221: std_logic; attribute dont_touch of WX2221: signal is true;
	signal WX2222: std_logic; attribute dont_touch of WX2222: signal is true;
	signal WX2223: std_logic; attribute dont_touch of WX2223: signal is true;
	signal WX2224: std_logic; attribute dont_touch of WX2224: signal is true;
	signal WX2225: std_logic; attribute dont_touch of WX2225: signal is true;
	signal WX2226: std_logic; attribute dont_touch of WX2226: signal is true;
	signal WX2227: std_logic; attribute dont_touch of WX2227: signal is true;
	signal WX2228: std_logic; attribute dont_touch of WX2228: signal is true;
	signal WX2229: std_logic; attribute dont_touch of WX2229: signal is true;
	signal WX2230: std_logic; attribute dont_touch of WX2230: signal is true;
	signal WX2231: std_logic; attribute dont_touch of WX2231: signal is true;
	signal WX2232: std_logic; attribute dont_touch of WX2232: signal is true;
	signal WX2233: std_logic; attribute dont_touch of WX2233: signal is true;
	signal WX2234: std_logic; attribute dont_touch of WX2234: signal is true;
	signal WX2235: std_logic; attribute dont_touch of WX2235: signal is true;
	signal WX2236: std_logic; attribute dont_touch of WX2236: signal is true;
	signal WX2237: std_logic; attribute dont_touch of WX2237: signal is true;
	signal WX2238: std_logic; attribute dont_touch of WX2238: signal is true;
	signal WX2239: std_logic; attribute dont_touch of WX2239: signal is true;
	signal WX2240: std_logic; attribute dont_touch of WX2240: signal is true;
	signal WX2241: std_logic; attribute dont_touch of WX2241: signal is true;
	signal WX2242: std_logic; attribute dont_touch of WX2242: signal is true;
	signal WX2243: std_logic; attribute dont_touch of WX2243: signal is true;
	signal WX2244: std_logic; attribute dont_touch of WX2244: signal is true;
	signal WX2245: std_logic; attribute dont_touch of WX2245: signal is true;
	signal WX2246: std_logic; attribute dont_touch of WX2246: signal is true;
	signal WX2247: std_logic; attribute dont_touch of WX2247: signal is true;
	signal WX2248: std_logic; attribute dont_touch of WX2248: signal is true;
	signal WX2249: std_logic; attribute dont_touch of WX2249: signal is true;
	signal WX2250: std_logic; attribute dont_touch of WX2250: signal is true;
	signal WX2251: std_logic; attribute dont_touch of WX2251: signal is true;
	signal WX2252: std_logic; attribute dont_touch of WX2252: signal is true;
	signal WX2253: std_logic; attribute dont_touch of WX2253: signal is true;
	signal WX2254: std_logic; attribute dont_touch of WX2254: signal is true;
	signal WX2255: std_logic; attribute dont_touch of WX2255: signal is true;
	signal WX2256: std_logic; attribute dont_touch of WX2256: signal is true;
	signal WX2257: std_logic; attribute dont_touch of WX2257: signal is true;
	signal WX2258: std_logic; attribute dont_touch of WX2258: signal is true;
	signal WX2259: std_logic; attribute dont_touch of WX2259: signal is true;
	signal WX2260: std_logic; attribute dont_touch of WX2260: signal is true;
	signal WX2261: std_logic; attribute dont_touch of WX2261: signal is true;
	signal WX2262: std_logic; attribute dont_touch of WX2262: signal is true;
	signal WX2263: std_logic; attribute dont_touch of WX2263: signal is true;
	signal WX2264: std_logic; attribute dont_touch of WX2264: signal is true;
	signal WX2265: std_logic; attribute dont_touch of WX2265: signal is true;
	signal WX2266: std_logic; attribute dont_touch of WX2266: signal is true;
	signal WX2267: std_logic; attribute dont_touch of WX2267: signal is true;
	signal WX2268: std_logic; attribute dont_touch of WX2268: signal is true;
	signal WX2269: std_logic; attribute dont_touch of WX2269: signal is true;
	signal WX2270: std_logic; attribute dont_touch of WX2270: signal is true;
	signal WX2271: std_logic; attribute dont_touch of WX2271: signal is true;
	signal WX2272: std_logic; attribute dont_touch of WX2272: signal is true;
	signal WX2273: std_logic; attribute dont_touch of WX2273: signal is true;
	signal WX2274: std_logic; attribute dont_touch of WX2274: signal is true;
	signal WX2275: std_logic; attribute dont_touch of WX2275: signal is true;
	signal WX2276: std_logic; attribute dont_touch of WX2276: signal is true;
	signal WX2277: std_logic; attribute dont_touch of WX2277: signal is true;
	signal WX2278: std_logic; attribute dont_touch of WX2278: signal is true;
	signal WX2279: std_logic; attribute dont_touch of WX2279: signal is true;
	signal WX2280: std_logic; attribute dont_touch of WX2280: signal is true;
	signal WX2281: std_logic; attribute dont_touch of WX2281: signal is true;
	signal WX2282: std_logic; attribute dont_touch of WX2282: signal is true;
	signal WX2283: std_logic; attribute dont_touch of WX2283: signal is true;
	signal WX2284: std_logic; attribute dont_touch of WX2284: signal is true;
	signal WX2285: std_logic; attribute dont_touch of WX2285: signal is true;
	signal WX2286: std_logic; attribute dont_touch of WX2286: signal is true;
	signal WX2287: std_logic; attribute dont_touch of WX2287: signal is true;
	signal WX2288: std_logic; attribute dont_touch of WX2288: signal is true;
	signal WX2289: std_logic; attribute dont_touch of WX2289: signal is true;
	signal WX2290: std_logic; attribute dont_touch of WX2290: signal is true;
	signal WX2291: std_logic; attribute dont_touch of WX2291: signal is true;
	signal WX2292: std_logic; attribute dont_touch of WX2292: signal is true;
	signal WX2293: std_logic; attribute dont_touch of WX2293: signal is true;
	signal WX2294: std_logic; attribute dont_touch of WX2294: signal is true;
	signal WX2295: std_logic; attribute dont_touch of WX2295: signal is true;
	signal WX2296: std_logic; attribute dont_touch of WX2296: signal is true;
	signal WX2297: std_logic; attribute dont_touch of WX2297: signal is true;
	signal WX2298: std_logic; attribute dont_touch of WX2298: signal is true;
	signal WX2299: std_logic; attribute dont_touch of WX2299: signal is true;
	signal WX2300: std_logic; attribute dont_touch of WX2300: signal is true;
	signal WX2301: std_logic; attribute dont_touch of WX2301: signal is true;
	signal WX2302: std_logic; attribute dont_touch of WX2302: signal is true;
	signal WX2303: std_logic; attribute dont_touch of WX2303: signal is true;
	signal WX2304: std_logic; attribute dont_touch of WX2304: signal is true;
	signal WX2305: std_logic; attribute dont_touch of WX2305: signal is true;
	signal WX2306: std_logic; attribute dont_touch of WX2306: signal is true;
	signal WX2307: std_logic; attribute dont_touch of WX2307: signal is true;
	signal WX2308: std_logic; attribute dont_touch of WX2308: signal is true;
	signal WX2309: std_logic; attribute dont_touch of WX2309: signal is true;
	signal WX2310: std_logic; attribute dont_touch of WX2310: signal is true;
	signal WX2311: std_logic; attribute dont_touch of WX2311: signal is true;
	signal WX2312: std_logic; attribute dont_touch of WX2312: signal is true;
	signal WX2313: std_logic; attribute dont_touch of WX2313: signal is true;
	signal WX2314: std_logic; attribute dont_touch of WX2314: signal is true;
	signal WX2315: std_logic; attribute dont_touch of WX2315: signal is true;
	signal WX2316: std_logic; attribute dont_touch of WX2316: signal is true;
	signal WX2317: std_logic; attribute dont_touch of WX2317: signal is true;
	signal WX2318: std_logic; attribute dont_touch of WX2318: signal is true;
	signal WX2319: std_logic; attribute dont_touch of WX2319: signal is true;
	signal WX2320: std_logic; attribute dont_touch of WX2320: signal is true;
	signal WX2321: std_logic; attribute dont_touch of WX2321: signal is true;
	signal WX2322: std_logic; attribute dont_touch of WX2322: signal is true;
	signal WX2323: std_logic; attribute dont_touch of WX2323: signal is true;
	signal WX2324: std_logic; attribute dont_touch of WX2324: signal is true;
	signal WX2325: std_logic; attribute dont_touch of WX2325: signal is true;
	signal WX2326: std_logic; attribute dont_touch of WX2326: signal is true;
	signal WX2327: std_logic; attribute dont_touch of WX2327: signal is true;
	signal WX2328: std_logic; attribute dont_touch of WX2328: signal is true;
	signal WX2329: std_logic; attribute dont_touch of WX2329: signal is true;
	signal WX2330: std_logic; attribute dont_touch of WX2330: signal is true;
	signal WX2331: std_logic; attribute dont_touch of WX2331: signal is true;
	signal WX2332: std_logic; attribute dont_touch of WX2332: signal is true;
	signal WX2333: std_logic; attribute dont_touch of WX2333: signal is true;
	signal WX2334: std_logic; attribute dont_touch of WX2334: signal is true;
	signal WX2335: std_logic; attribute dont_touch of WX2335: signal is true;
	signal WX2336: std_logic; attribute dont_touch of WX2336: signal is true;
	signal WX2337: std_logic; attribute dont_touch of WX2337: signal is true;
	signal WX2338: std_logic; attribute dont_touch of WX2338: signal is true;
	signal WX2339: std_logic; attribute dont_touch of WX2339: signal is true;
	signal WX2340: std_logic; attribute dont_touch of WX2340: signal is true;
	signal WX2341: std_logic; attribute dont_touch of WX2341: signal is true;
	signal WX2342: std_logic; attribute dont_touch of WX2342: signal is true;
	signal WX2343: std_logic; attribute dont_touch of WX2343: signal is true;
	signal WX2344: std_logic; attribute dont_touch of WX2344: signal is true;
	signal WX2345: std_logic; attribute dont_touch of WX2345: signal is true;
	signal WX2346: std_logic; attribute dont_touch of WX2346: signal is true;
	signal WX2347: std_logic; attribute dont_touch of WX2347: signal is true;
	signal WX2348: std_logic; attribute dont_touch of WX2348: signal is true;
	signal WX2349: std_logic; attribute dont_touch of WX2349: signal is true;
	signal WX2350: std_logic; attribute dont_touch of WX2350: signal is true;
	signal WX2351: std_logic; attribute dont_touch of WX2351: signal is true;
	signal WX2352: std_logic; attribute dont_touch of WX2352: signal is true;
	signal WX2353: std_logic; attribute dont_touch of WX2353: signal is true;
	signal WX2354: std_logic; attribute dont_touch of WX2354: signal is true;
	signal WX2355: std_logic; attribute dont_touch of WX2355: signal is true;
	signal WX2356: std_logic; attribute dont_touch of WX2356: signal is true;
	signal WX2357: std_logic; attribute dont_touch of WX2357: signal is true;
	signal WX2358: std_logic; attribute dont_touch of WX2358: signal is true;
	signal WX2359: std_logic; attribute dont_touch of WX2359: signal is true;
	signal WX2360: std_logic; attribute dont_touch of WX2360: signal is true;
	signal WX2361: std_logic; attribute dont_touch of WX2361: signal is true;
	signal WX2362: std_logic; attribute dont_touch of WX2362: signal is true;
	signal WX2363: std_logic; attribute dont_touch of WX2363: signal is true;
	signal WX2364: std_logic; attribute dont_touch of WX2364: signal is true;
	signal WX2365: std_logic; attribute dont_touch of WX2365: signal is true;
	signal WX2366: std_logic; attribute dont_touch of WX2366: signal is true;
	signal WX2367: std_logic; attribute dont_touch of WX2367: signal is true;
	signal WX2368: std_logic; attribute dont_touch of WX2368: signal is true;
	signal WX2369: std_logic; attribute dont_touch of WX2369: signal is true;
	signal WX2370: std_logic; attribute dont_touch of WX2370: signal is true;
	signal WX2371: std_logic; attribute dont_touch of WX2371: signal is true;
	signal WX2372: std_logic; attribute dont_touch of WX2372: signal is true;
	signal WX2373: std_logic; attribute dont_touch of WX2373: signal is true;
	signal WX2374: std_logic; attribute dont_touch of WX2374: signal is true;
	signal WX2375: std_logic; attribute dont_touch of WX2375: signal is true;
	signal WX2376: std_logic; attribute dont_touch of WX2376: signal is true;
	signal WX2377: std_logic; attribute dont_touch of WX2377: signal is true;
	signal WX2378: std_logic; attribute dont_touch of WX2378: signal is true;
	signal WX2379: std_logic; attribute dont_touch of WX2379: signal is true;
	signal WX2380: std_logic; attribute dont_touch of WX2380: signal is true;
	signal WX2381: std_logic; attribute dont_touch of WX2381: signal is true;
	signal WX2382: std_logic; attribute dont_touch of WX2382: signal is true;
	signal WX2383: std_logic; attribute dont_touch of WX2383: signal is true;
	signal WX2384: std_logic; attribute dont_touch of WX2384: signal is true;
	signal WX2385: std_logic; attribute dont_touch of WX2385: signal is true;
	signal WX2386: std_logic; attribute dont_touch of WX2386: signal is true;
	signal WX2387: std_logic; attribute dont_touch of WX2387: signal is true;
	signal WX2388: std_logic; attribute dont_touch of WX2388: signal is true;
	signal WX2389: std_logic; attribute dont_touch of WX2389: signal is true;
	signal WX2390: std_logic; attribute dont_touch of WX2390: signal is true;
	signal WX2391: std_logic; attribute dont_touch of WX2391: signal is true;
	signal WX2392: std_logic; attribute dont_touch of WX2392: signal is true;
	signal WX2393: std_logic; attribute dont_touch of WX2393: signal is true;
	signal WX2394: std_logic; attribute dont_touch of WX2394: signal is true;
	signal WX2395: std_logic; attribute dont_touch of WX2395: signal is true;
	signal WX2396: std_logic; attribute dont_touch of WX2396: signal is true;
	signal WX2397: std_logic; attribute dont_touch of WX2397: signal is true;
	signal WX2398: std_logic; attribute dont_touch of WX2398: signal is true;
	signal WX2399: std_logic; attribute dont_touch of WX2399: signal is true;
	signal WX2400: std_logic; attribute dont_touch of WX2400: signal is true;
	signal WX2401: std_logic; attribute dont_touch of WX2401: signal is true;
	signal WX2402: std_logic; attribute dont_touch of WX2402: signal is true;
	signal WX2403: std_logic; attribute dont_touch of WX2403: signal is true;
	signal WX2404: std_logic; attribute dont_touch of WX2404: signal is true;
	signal WX2405: std_logic; attribute dont_touch of WX2405: signal is true;
	signal WX2406: std_logic; attribute dont_touch of WX2406: signal is true;
	signal WX2407: std_logic; attribute dont_touch of WX2407: signal is true;
	signal WX2408: std_logic; attribute dont_touch of WX2408: signal is true;
	signal WX2409: std_logic; attribute dont_touch of WX2409: signal is true;
	signal WX2410: std_logic; attribute dont_touch of WX2410: signal is true;
	signal WX2411: std_logic; attribute dont_touch of WX2411: signal is true;
	signal WX2412: std_logic; attribute dont_touch of WX2412: signal is true;
	signal WX2413: std_logic; attribute dont_touch of WX2413: signal is true;
	signal WX2414: std_logic; attribute dont_touch of WX2414: signal is true;
	signal WX2415: std_logic; attribute dont_touch of WX2415: signal is true;
	signal WX2416: std_logic; attribute dont_touch of WX2416: signal is true;
	signal WX2417: std_logic; attribute dont_touch of WX2417: signal is true;
	signal WX2418: std_logic; attribute dont_touch of WX2418: signal is true;
	signal WX2419: std_logic; attribute dont_touch of WX2419: signal is true;
	signal WX2420: std_logic; attribute dont_touch of WX2420: signal is true;
	signal WX2421: std_logic; attribute dont_touch of WX2421: signal is true;
	signal WX2422: std_logic; attribute dont_touch of WX2422: signal is true;
	signal WX2423: std_logic; attribute dont_touch of WX2423: signal is true;
	signal WX2424: std_logic; attribute dont_touch of WX2424: signal is true;
	signal WX2425: std_logic; attribute dont_touch of WX2425: signal is true;
	signal WX2426: std_logic; attribute dont_touch of WX2426: signal is true;
	signal WX2427: std_logic; attribute dont_touch of WX2427: signal is true;
	signal WX2428: std_logic; attribute dont_touch of WX2428: signal is true;
	signal WX2429: std_logic; attribute dont_touch of WX2429: signal is true;
	signal WX2430: std_logic; attribute dont_touch of WX2430: signal is true;
	signal WX2431: std_logic; attribute dont_touch of WX2431: signal is true;
	signal WX2432: std_logic; attribute dont_touch of WX2432: signal is true;
	signal WX2433: std_logic; attribute dont_touch of WX2433: signal is true;
	signal WX2434: std_logic; attribute dont_touch of WX2434: signal is true;
	signal WX2435: std_logic; attribute dont_touch of WX2435: signal is true;
	signal WX2436: std_logic; attribute dont_touch of WX2436: signal is true;
	signal WX2437: std_logic; attribute dont_touch of WX2437: signal is true;
	signal WX2438: std_logic; attribute dont_touch of WX2438: signal is true;
	signal WX2439: std_logic; attribute dont_touch of WX2439: signal is true;
	signal WX2440: std_logic; attribute dont_touch of WX2440: signal is true;
	signal WX2441: std_logic; attribute dont_touch of WX2441: signal is true;
	signal WX2442: std_logic; attribute dont_touch of WX2442: signal is true;
	signal WX2443: std_logic; attribute dont_touch of WX2443: signal is true;
	signal WX2444: std_logic; attribute dont_touch of WX2444: signal is true;
	signal WX2445: std_logic; attribute dont_touch of WX2445: signal is true;
	signal WX2446: std_logic; attribute dont_touch of WX2446: signal is true;
	signal WX2447: std_logic; attribute dont_touch of WX2447: signal is true;
	signal WX2448: std_logic; attribute dont_touch of WX2448: signal is true;
	signal WX2449: std_logic; attribute dont_touch of WX2449: signal is true;
	signal WX2450: std_logic; attribute dont_touch of WX2450: signal is true;
	signal WX2451: std_logic; attribute dont_touch of WX2451: signal is true;
	signal WX2452: std_logic; attribute dont_touch of WX2452: signal is true;
	signal WX2453: std_logic; attribute dont_touch of WX2453: signal is true;
	signal WX2454: std_logic; attribute dont_touch of WX2454: signal is true;
	signal WX2455: std_logic; attribute dont_touch of WX2455: signal is true;
	signal WX2456: std_logic; attribute dont_touch of WX2456: signal is true;
	signal WX2457: std_logic; attribute dont_touch of WX2457: signal is true;
	signal WX2458: std_logic; attribute dont_touch of WX2458: signal is true;
	signal WX2459: std_logic; attribute dont_touch of WX2459: signal is true;
	signal WX2460: std_logic; attribute dont_touch of WX2460: signal is true;
	signal WX2461: std_logic; attribute dont_touch of WX2461: signal is true;
	signal WX2462: std_logic; attribute dont_touch of WX2462: signal is true;
	signal WX2463: std_logic; attribute dont_touch of WX2463: signal is true;
	signal WX2464: std_logic; attribute dont_touch of WX2464: signal is true;
	signal WX2465: std_logic; attribute dont_touch of WX2465: signal is true;
	signal WX2466: std_logic; attribute dont_touch of WX2466: signal is true;
	signal WX2467: std_logic; attribute dont_touch of WX2467: signal is true;
	signal WX2468: std_logic; attribute dont_touch of WX2468: signal is true;
	signal WX2469: std_logic; attribute dont_touch of WX2469: signal is true;
	signal WX2470: std_logic; attribute dont_touch of WX2470: signal is true;
	signal WX2471: std_logic; attribute dont_touch of WX2471: signal is true;
	signal WX2472: std_logic; attribute dont_touch of WX2472: signal is true;
	signal WX2473: std_logic; attribute dont_touch of WX2473: signal is true;
	signal WX2474: std_logic; attribute dont_touch of WX2474: signal is true;
	signal WX2475: std_logic; attribute dont_touch of WX2475: signal is true;
	signal WX2476: std_logic; attribute dont_touch of WX2476: signal is true;
	signal WX2477: std_logic; attribute dont_touch of WX2477: signal is true;
	signal WX2478: std_logic; attribute dont_touch of WX2478: signal is true;
	signal WX2479: std_logic; attribute dont_touch of WX2479: signal is true;
	signal WX2480: std_logic; attribute dont_touch of WX2480: signal is true;
	signal WX2481: std_logic; attribute dont_touch of WX2481: signal is true;
	signal WX2482: std_logic; attribute dont_touch of WX2482: signal is true;
	signal WX2483: std_logic; attribute dont_touch of WX2483: signal is true;
	signal WX2484: std_logic; attribute dont_touch of WX2484: signal is true;
	signal WX2485: std_logic; attribute dont_touch of WX2485: signal is true;
	signal WX2486: std_logic; attribute dont_touch of WX2486: signal is true;
	signal WX2487: std_logic; attribute dont_touch of WX2487: signal is true;
	signal WX2488: std_logic; attribute dont_touch of WX2488: signal is true;
	signal WX2489: std_logic; attribute dont_touch of WX2489: signal is true;
	signal WX2490: std_logic; attribute dont_touch of WX2490: signal is true;
	signal WX2491: std_logic; attribute dont_touch of WX2491: signal is true;
	signal WX2492: std_logic; attribute dont_touch of WX2492: signal is true;
	signal WX2493: std_logic; attribute dont_touch of WX2493: signal is true;
	signal WX2494: std_logic; attribute dont_touch of WX2494: signal is true;
	signal WX2495: std_logic; attribute dont_touch of WX2495: signal is true;
	signal WX2496: std_logic; attribute dont_touch of WX2496: signal is true;
	signal WX2497: std_logic; attribute dont_touch of WX2497: signal is true;
	signal WX2498: std_logic; attribute dont_touch of WX2498: signal is true;
	signal WX2499: std_logic; attribute dont_touch of WX2499: signal is true;
	signal WX2500: std_logic; attribute dont_touch of WX2500: signal is true;
	signal WX2501: std_logic; attribute dont_touch of WX2501: signal is true;
	signal WX2502: std_logic; attribute dont_touch of WX2502: signal is true;
	signal WX2503: std_logic; attribute dont_touch of WX2503: signal is true;
	signal WX2504: std_logic; attribute dont_touch of WX2504: signal is true;
	signal WX2505: std_logic; attribute dont_touch of WX2505: signal is true;
	signal WX2506: std_logic; attribute dont_touch of WX2506: signal is true;
	signal WX2507: std_logic; attribute dont_touch of WX2507: signal is true;
	signal WX2508: std_logic; attribute dont_touch of WX2508: signal is true;
	signal WX2509: std_logic; attribute dont_touch of WX2509: signal is true;
	signal WX2510: std_logic; attribute dont_touch of WX2510: signal is true;
	signal WX2511: std_logic; attribute dont_touch of WX2511: signal is true;
	signal WX2512: std_logic; attribute dont_touch of WX2512: signal is true;
	signal WX2513: std_logic; attribute dont_touch of WX2513: signal is true;
	signal WX2514: std_logic; attribute dont_touch of WX2514: signal is true;
	signal WX2515: std_logic; attribute dont_touch of WX2515: signal is true;
	signal WX2516: std_logic; attribute dont_touch of WX2516: signal is true;
	signal WX2517: std_logic; attribute dont_touch of WX2517: signal is true;
	signal WX2518: std_logic; attribute dont_touch of WX2518: signal is true;
	signal WX2519: std_logic; attribute dont_touch of WX2519: signal is true;
	signal WX2520: std_logic; attribute dont_touch of WX2520: signal is true;
	signal WX2521: std_logic; attribute dont_touch of WX2521: signal is true;
	signal WX2522: std_logic; attribute dont_touch of WX2522: signal is true;
	signal WX2523: std_logic; attribute dont_touch of WX2523: signal is true;
	signal WX2524: std_logic; attribute dont_touch of WX2524: signal is true;
	signal WX2525: std_logic; attribute dont_touch of WX2525: signal is true;
	signal WX2526: std_logic; attribute dont_touch of WX2526: signal is true;
	signal WX2527: std_logic; attribute dont_touch of WX2527: signal is true;
	signal WX2528: std_logic; attribute dont_touch of WX2528: signal is true;
	signal WX2529: std_logic; attribute dont_touch of WX2529: signal is true;
	signal WX2530: std_logic; attribute dont_touch of WX2530: signal is true;
	signal WX2531: std_logic; attribute dont_touch of WX2531: signal is true;
	signal WX2532: std_logic; attribute dont_touch of WX2532: signal is true;
	signal WX2533: std_logic; attribute dont_touch of WX2533: signal is true;
	signal WX2534: std_logic; attribute dont_touch of WX2534: signal is true;
	signal WX2535: std_logic; attribute dont_touch of WX2535: signal is true;
	signal WX2536: std_logic; attribute dont_touch of WX2536: signal is true;
	signal WX2537: std_logic; attribute dont_touch of WX2537: signal is true;
	signal WX2538: std_logic; attribute dont_touch of WX2538: signal is true;
	signal WX2539: std_logic; attribute dont_touch of WX2539: signal is true;
	signal WX2540: std_logic; attribute dont_touch of WX2540: signal is true;
	signal WX2541: std_logic; attribute dont_touch of WX2541: signal is true;
	signal WX2542: std_logic; attribute dont_touch of WX2542: signal is true;
	signal WX2543: std_logic; attribute dont_touch of WX2543: signal is true;
	signal WX2544: std_logic; attribute dont_touch of WX2544: signal is true;
	signal WX2545: std_logic; attribute dont_touch of WX2545: signal is true;
	signal WX2546: std_logic; attribute dont_touch of WX2546: signal is true;
	signal WX2547: std_logic; attribute dont_touch of WX2547: signal is true;
	signal WX2548: std_logic; attribute dont_touch of WX2548: signal is true;
	signal WX2549: std_logic; attribute dont_touch of WX2549: signal is true;
	signal WX2550: std_logic; attribute dont_touch of WX2550: signal is true;
	signal WX2551: std_logic; attribute dont_touch of WX2551: signal is true;
	signal WX2552: std_logic; attribute dont_touch of WX2552: signal is true;
	signal WX2553: std_logic; attribute dont_touch of WX2553: signal is true;
	signal WX2554: std_logic; attribute dont_touch of WX2554: signal is true;
	signal WX2555: std_logic; attribute dont_touch of WX2555: signal is true;
	signal WX2556: std_logic; attribute dont_touch of WX2556: signal is true;
	signal WX2557: std_logic; attribute dont_touch of WX2557: signal is true;
	signal WX2559: std_logic; attribute dont_touch of WX2559: signal is true;
	signal WX2561: std_logic; attribute dont_touch of WX2561: signal is true;
	signal WX2563: std_logic; attribute dont_touch of WX2563: signal is true;
	signal WX2565: std_logic; attribute dont_touch of WX2565: signal is true;
	signal WX2567: std_logic; attribute dont_touch of WX2567: signal is true;
	signal WX2569: std_logic; attribute dont_touch of WX2569: signal is true;
	signal WX2571: std_logic; attribute dont_touch of WX2571: signal is true;
	signal WX2573: std_logic; attribute dont_touch of WX2573: signal is true;
	signal WX2575: std_logic; attribute dont_touch of WX2575: signal is true;
	signal WX2577: std_logic; attribute dont_touch of WX2577: signal is true;
	signal WX2579: std_logic; attribute dont_touch of WX2579: signal is true;
	signal WX2581: std_logic; attribute dont_touch of WX2581: signal is true;
	signal WX2583: std_logic; attribute dont_touch of WX2583: signal is true;
	signal WX2585: std_logic; attribute dont_touch of WX2585: signal is true;
	signal WX2587: std_logic; attribute dont_touch of WX2587: signal is true;
	signal WX2589: std_logic; attribute dont_touch of WX2589: signal is true;
	signal WX2591: std_logic; attribute dont_touch of WX2591: signal is true;
	signal WX2593: std_logic; attribute dont_touch of WX2593: signal is true;
	signal WX2595: std_logic; attribute dont_touch of WX2595: signal is true;
	signal WX2597: std_logic; attribute dont_touch of WX2597: signal is true;
	signal WX2599: std_logic; attribute dont_touch of WX2599: signal is true;
	signal WX2601: std_logic; attribute dont_touch of WX2601: signal is true;
	signal WX2603: std_logic; attribute dont_touch of WX2603: signal is true;
	signal WX2605: std_logic; attribute dont_touch of WX2605: signal is true;
	signal WX2607: std_logic; attribute dont_touch of WX2607: signal is true;
	signal WX2609: std_logic; attribute dont_touch of WX2609: signal is true;
	signal WX2611: std_logic; attribute dont_touch of WX2611: signal is true;
	signal WX2613: std_logic; attribute dont_touch of WX2613: signal is true;
	signal WX2615: std_logic; attribute dont_touch of WX2615: signal is true;
	signal WX2617: std_logic; attribute dont_touch of WX2617: signal is true;
	signal WX2619: std_logic; attribute dont_touch of WX2619: signal is true;
	signal WX2621: std_logic; attribute dont_touch of WX2621: signal is true;
	signal WX2622: std_logic; attribute dont_touch of WX2622: signal is true;
	signal WX2623: std_logic; attribute dont_touch of WX2623: signal is true;
	signal WX2624: std_logic; attribute dont_touch of WX2624: signal is true;
	signal WX2625: std_logic; attribute dont_touch of WX2625: signal is true;
	signal WX2626: std_logic; attribute dont_touch of WX2626: signal is true;
	signal WX2627: std_logic; attribute dont_touch of WX2627: signal is true;
	signal WX2628: std_logic; attribute dont_touch of WX2628: signal is true;
	signal WX2629: std_logic; attribute dont_touch of WX2629: signal is true;
	signal WX2630: std_logic; attribute dont_touch of WX2630: signal is true;
	signal WX2631: std_logic; attribute dont_touch of WX2631: signal is true;
	signal WX2632: std_logic; attribute dont_touch of WX2632: signal is true;
	signal WX2633: std_logic; attribute dont_touch of WX2633: signal is true;
	signal WX2634: std_logic; attribute dont_touch of WX2634: signal is true;
	signal WX2635: std_logic; attribute dont_touch of WX2635: signal is true;
	signal WX2636: std_logic; attribute dont_touch of WX2636: signal is true;
	signal WX2637: std_logic; attribute dont_touch of WX2637: signal is true;
	signal WX2638: std_logic; attribute dont_touch of WX2638: signal is true;
	signal WX2639: std_logic; attribute dont_touch of WX2639: signal is true;
	signal WX2640: std_logic; attribute dont_touch of WX2640: signal is true;
	signal WX2641: std_logic; attribute dont_touch of WX2641: signal is true;
	signal WX2642: std_logic; attribute dont_touch of WX2642: signal is true;
	signal WX2643: std_logic; attribute dont_touch of WX2643: signal is true;
	signal WX2644: std_logic; attribute dont_touch of WX2644: signal is true;
	signal WX2645: std_logic; attribute dont_touch of WX2645: signal is true;
	signal WX2646: std_logic; attribute dont_touch of WX2646: signal is true;
	signal WX2647: std_logic; attribute dont_touch of WX2647: signal is true;
	signal WX2648: std_logic; attribute dont_touch of WX2648: signal is true;
	signal WX2649: std_logic; attribute dont_touch of WX2649: signal is true;
	signal WX2650: std_logic; attribute dont_touch of WX2650: signal is true;
	signal WX2651: std_logic; attribute dont_touch of WX2651: signal is true;
	signal WX2652: std_logic; attribute dont_touch of WX2652: signal is true;
	signal WX2653: std_logic; attribute dont_touch of WX2653: signal is true;
	signal WX2654: std_logic; attribute dont_touch of WX2654: signal is true;
	signal WX2655: std_logic; attribute dont_touch of WX2655: signal is true;
	signal WX2656: std_logic; attribute dont_touch of WX2656: signal is true;
	signal WX2657: std_logic; attribute dont_touch of WX2657: signal is true;
	signal WX2658: std_logic; attribute dont_touch of WX2658: signal is true;
	signal WX2659: std_logic; attribute dont_touch of WX2659: signal is true;
	signal WX2660: std_logic; attribute dont_touch of WX2660: signal is true;
	signal WX2661: std_logic; attribute dont_touch of WX2661: signal is true;
	signal WX2662: std_logic; attribute dont_touch of WX2662: signal is true;
	signal WX2663: std_logic; attribute dont_touch of WX2663: signal is true;
	signal WX2664: std_logic; attribute dont_touch of WX2664: signal is true;
	signal WX2665: std_logic; attribute dont_touch of WX2665: signal is true;
	signal WX2666: std_logic; attribute dont_touch of WX2666: signal is true;
	signal WX2667: std_logic; attribute dont_touch of WX2667: signal is true;
	signal WX2668: std_logic; attribute dont_touch of WX2668: signal is true;
	signal WX2669: std_logic; attribute dont_touch of WX2669: signal is true;
	signal WX2670: std_logic; attribute dont_touch of WX2670: signal is true;
	signal WX2671: std_logic; attribute dont_touch of WX2671: signal is true;
	signal WX2672: std_logic; attribute dont_touch of WX2672: signal is true;
	signal WX2673: std_logic; attribute dont_touch of WX2673: signal is true;
	signal WX2674: std_logic; attribute dont_touch of WX2674: signal is true;
	signal WX2675: std_logic; attribute dont_touch of WX2675: signal is true;
	signal WX2676: std_logic; attribute dont_touch of WX2676: signal is true;
	signal WX2677: std_logic; attribute dont_touch of WX2677: signal is true;
	signal WX2678: std_logic; attribute dont_touch of WX2678: signal is true;
	signal WX2679: std_logic; attribute dont_touch of WX2679: signal is true;
	signal WX2680: std_logic; attribute dont_touch of WX2680: signal is true;
	signal WX2681: std_logic; attribute dont_touch of WX2681: signal is true;
	signal WX2682: std_logic; attribute dont_touch of WX2682: signal is true;
	signal WX2683: std_logic; attribute dont_touch of WX2683: signal is true;
	signal WX2684: std_logic; attribute dont_touch of WX2684: signal is true;
	signal WX2685: std_logic; attribute dont_touch of WX2685: signal is true;
	signal WX2686: std_logic; attribute dont_touch of WX2686: signal is true;
	signal WX2687: std_logic; attribute dont_touch of WX2687: signal is true;
	signal WX2688: std_logic; attribute dont_touch of WX2688: signal is true;
	signal WX2689: std_logic; attribute dont_touch of WX2689: signal is true;
	signal WX2690: std_logic; attribute dont_touch of WX2690: signal is true;
	signal WX2691: std_logic; attribute dont_touch of WX2691: signal is true;
	signal WX2692: std_logic; attribute dont_touch of WX2692: signal is true;
	signal WX2693: std_logic; attribute dont_touch of WX2693: signal is true;
	signal WX2694: std_logic; attribute dont_touch of WX2694: signal is true;
	signal WX2695: std_logic; attribute dont_touch of WX2695: signal is true;
	signal WX2696: std_logic; attribute dont_touch of WX2696: signal is true;
	signal WX2697: std_logic; attribute dont_touch of WX2697: signal is true;
	signal WX2698: std_logic; attribute dont_touch of WX2698: signal is true;
	signal WX2699: std_logic; attribute dont_touch of WX2699: signal is true;
	signal WX2700: std_logic; attribute dont_touch of WX2700: signal is true;
	signal WX2701: std_logic; attribute dont_touch of WX2701: signal is true;
	signal WX2702: std_logic; attribute dont_touch of WX2702: signal is true;
	signal WX2703: std_logic; attribute dont_touch of WX2703: signal is true;
	signal WX2704: std_logic; attribute dont_touch of WX2704: signal is true;
	signal WX2705: std_logic; attribute dont_touch of WX2705: signal is true;
	signal WX2706: std_logic; attribute dont_touch of WX2706: signal is true;
	signal WX2707: std_logic; attribute dont_touch of WX2707: signal is true;
	signal WX2708: std_logic; attribute dont_touch of WX2708: signal is true;
	signal WX2709: std_logic; attribute dont_touch of WX2709: signal is true;
	signal WX2710: std_logic; attribute dont_touch of WX2710: signal is true;
	signal WX2711: std_logic; attribute dont_touch of WX2711: signal is true;
	signal WX2712: std_logic; attribute dont_touch of WX2712: signal is true;
	signal WX2713: std_logic; attribute dont_touch of WX2713: signal is true;
	signal WX2714: std_logic; attribute dont_touch of WX2714: signal is true;
	signal WX2715: std_logic; attribute dont_touch of WX2715: signal is true;
	signal WX2716: std_logic; attribute dont_touch of WX2716: signal is true;
	signal WX2717: std_logic; attribute dont_touch of WX2717: signal is true;
	signal WX2718: std_logic; attribute dont_touch of WX2718: signal is true;
	signal WX2719: std_logic; attribute dont_touch of WX2719: signal is true;
	signal WX2720: std_logic; attribute dont_touch of WX2720: signal is true;
	signal WX2721: std_logic; attribute dont_touch of WX2721: signal is true;
	signal WX2722: std_logic; attribute dont_touch of WX2722: signal is true;
	signal WX2723: std_logic; attribute dont_touch of WX2723: signal is true;
	signal WX2724: std_logic; attribute dont_touch of WX2724: signal is true;
	signal WX2725: std_logic; attribute dont_touch of WX2725: signal is true;
	signal WX2726: std_logic; attribute dont_touch of WX2726: signal is true;
	signal WX2727: std_logic; attribute dont_touch of WX2727: signal is true;
	signal WX2728: std_logic; attribute dont_touch of WX2728: signal is true;
	signal WX2729: std_logic; attribute dont_touch of WX2729: signal is true;
	signal WX2730: std_logic; attribute dont_touch of WX2730: signal is true;
	signal WX2731: std_logic; attribute dont_touch of WX2731: signal is true;
	signal WX2732: std_logic; attribute dont_touch of WX2732: signal is true;
	signal WX2733: std_logic; attribute dont_touch of WX2733: signal is true;
	signal WX2734: std_logic; attribute dont_touch of WX2734: signal is true;
	signal WX2735: std_logic; attribute dont_touch of WX2735: signal is true;
	signal WX2736: std_logic; attribute dont_touch of WX2736: signal is true;
	signal WX2737: std_logic; attribute dont_touch of WX2737: signal is true;
	signal WX2738: std_logic; attribute dont_touch of WX2738: signal is true;
	signal WX2739: std_logic; attribute dont_touch of WX2739: signal is true;
	signal WX2740: std_logic; attribute dont_touch of WX2740: signal is true;
	signal WX2741: std_logic; attribute dont_touch of WX2741: signal is true;
	signal WX2742: std_logic; attribute dont_touch of WX2742: signal is true;
	signal WX2743: std_logic; attribute dont_touch of WX2743: signal is true;
	signal WX2744: std_logic; attribute dont_touch of WX2744: signal is true;
	signal WX2745: std_logic; attribute dont_touch of WX2745: signal is true;
	signal WX2746: std_logic; attribute dont_touch of WX2746: signal is true;
	signal WX2747: std_logic; attribute dont_touch of WX2747: signal is true;
	signal WX2748: std_logic; attribute dont_touch of WX2748: signal is true;
	signal WX2749: std_logic; attribute dont_touch of WX2749: signal is true;
	signal WX2750: std_logic; attribute dont_touch of WX2750: signal is true;
	signal WX2751: std_logic; attribute dont_touch of WX2751: signal is true;
	signal WX2752: std_logic; attribute dont_touch of WX2752: signal is true;
	signal WX2753: std_logic; attribute dont_touch of WX2753: signal is true;
	signal WX2754: std_logic; attribute dont_touch of WX2754: signal is true;
	signal WX2755: std_logic; attribute dont_touch of WX2755: signal is true;
	signal WX2756: std_logic; attribute dont_touch of WX2756: signal is true;
	signal WX2757: std_logic; attribute dont_touch of WX2757: signal is true;
	signal WX2758: std_logic; attribute dont_touch of WX2758: signal is true;
	signal WX2759: std_logic; attribute dont_touch of WX2759: signal is true;
	signal WX2760: std_logic; attribute dont_touch of WX2760: signal is true;
	signal WX2761: std_logic; attribute dont_touch of WX2761: signal is true;
	signal WX2762: std_logic; attribute dont_touch of WX2762: signal is true;
	signal WX2763: std_logic; attribute dont_touch of WX2763: signal is true;
	signal WX2764: std_logic; attribute dont_touch of WX2764: signal is true;
	signal WX2765: std_logic; attribute dont_touch of WX2765: signal is true;
	signal WX2766: std_logic; attribute dont_touch of WX2766: signal is true;
	signal WX2767: std_logic; attribute dont_touch of WX2767: signal is true;
	signal WX2768: std_logic; attribute dont_touch of WX2768: signal is true;
	signal WX2769: std_logic; attribute dont_touch of WX2769: signal is true;
	signal WX2770: std_logic; attribute dont_touch of WX2770: signal is true;
	signal WX2771: std_logic; attribute dont_touch of WX2771: signal is true;
	signal WX2772: std_logic; attribute dont_touch of WX2772: signal is true;
	signal WX2773: std_logic; attribute dont_touch of WX2773: signal is true;
	signal WX2774: std_logic; attribute dont_touch of WX2774: signal is true;
	signal WX2775: std_logic; attribute dont_touch of WX2775: signal is true;
	signal WX2776: std_logic; attribute dont_touch of WX2776: signal is true;
	signal WX2777: std_logic; attribute dont_touch of WX2777: signal is true;
	signal WX2778: std_logic; attribute dont_touch of WX2778: signal is true;
	signal WX2779: std_logic; attribute dont_touch of WX2779: signal is true;
	signal WX2780: std_logic; attribute dont_touch of WX2780: signal is true;
	signal WX2781: std_logic; attribute dont_touch of WX2781: signal is true;
	signal WX2782: std_logic; attribute dont_touch of WX2782: signal is true;
	signal WX2783: std_logic; attribute dont_touch of WX2783: signal is true;
	signal WX2784: std_logic; attribute dont_touch of WX2784: signal is true;
	signal WX2785: std_logic; attribute dont_touch of WX2785: signal is true;
	signal WX2786: std_logic; attribute dont_touch of WX2786: signal is true;
	signal WX2787: std_logic; attribute dont_touch of WX2787: signal is true;
	signal WX2788: std_logic; attribute dont_touch of WX2788: signal is true;
	signal WX2789: std_logic; attribute dont_touch of WX2789: signal is true;
	signal WX2790: std_logic; attribute dont_touch of WX2790: signal is true;
	signal WX2791: std_logic; attribute dont_touch of WX2791: signal is true;
	signal WX2792: std_logic; attribute dont_touch of WX2792: signal is true;
	signal WX2793: std_logic; attribute dont_touch of WX2793: signal is true;
	signal WX2794: std_logic; attribute dont_touch of WX2794: signal is true;
	signal WX2795: std_logic; attribute dont_touch of WX2795: signal is true;
	signal WX2796: std_logic; attribute dont_touch of WX2796: signal is true;
	signal WX2797: std_logic; attribute dont_touch of WX2797: signal is true;
	signal WX2798: std_logic; attribute dont_touch of WX2798: signal is true;
	signal WX2799: std_logic; attribute dont_touch of WX2799: signal is true;
	signal WX2800: std_logic; attribute dont_touch of WX2800: signal is true;
	signal WX2801: std_logic; attribute dont_touch of WX2801: signal is true;
	signal WX2802: std_logic; attribute dont_touch of WX2802: signal is true;
	signal WX2803: std_logic; attribute dont_touch of WX2803: signal is true;
	signal WX2804: std_logic; attribute dont_touch of WX2804: signal is true;
	signal WX2805: std_logic; attribute dont_touch of WX2805: signal is true;
	signal WX2806: std_logic; attribute dont_touch of WX2806: signal is true;
	signal WX2807: std_logic; attribute dont_touch of WX2807: signal is true;
	signal WX2808: std_logic; attribute dont_touch of WX2808: signal is true;
	signal WX2809: std_logic; attribute dont_touch of WX2809: signal is true;
	signal WX2810: std_logic; attribute dont_touch of WX2810: signal is true;
	signal WX2811: std_logic; attribute dont_touch of WX2811: signal is true;
	signal WX2812: std_logic; attribute dont_touch of WX2812: signal is true;
	signal WX2813: std_logic; attribute dont_touch of WX2813: signal is true;
	signal WX2814: std_logic; attribute dont_touch of WX2814: signal is true;
	signal WX2815: std_logic; attribute dont_touch of WX2815: signal is true;
	signal WX2816: std_logic; attribute dont_touch of WX2816: signal is true;
	signal WX2817: std_logic; attribute dont_touch of WX2817: signal is true;
	signal WX2818: std_logic; attribute dont_touch of WX2818: signal is true;
	signal WX2819: std_logic; attribute dont_touch of WX2819: signal is true;
	signal WX2820: std_logic; attribute dont_touch of WX2820: signal is true;
	signal WX2821: std_logic; attribute dont_touch of WX2821: signal is true;
	signal WX2822: std_logic; attribute dont_touch of WX2822: signal is true;
	signal WX2823: std_logic; attribute dont_touch of WX2823: signal is true;
	signal WX2824: std_logic; attribute dont_touch of WX2824: signal is true;
	signal WX2825: std_logic; attribute dont_touch of WX2825: signal is true;
	signal WX2826: std_logic; attribute dont_touch of WX2826: signal is true;
	signal WX2827: std_logic; attribute dont_touch of WX2827: signal is true;
	signal WX2828: std_logic; attribute dont_touch of WX2828: signal is true;
	signal WX2829: std_logic; attribute dont_touch of WX2829: signal is true;
	signal WX2830: std_logic; attribute dont_touch of WX2830: signal is true;
	signal WX2831: std_logic; attribute dont_touch of WX2831: signal is true;
	signal WX2832: std_logic; attribute dont_touch of WX2832: signal is true;
	signal WX2833: std_logic; attribute dont_touch of WX2833: signal is true;
	signal WX2834: std_logic; attribute dont_touch of WX2834: signal is true;
	signal WX2835: std_logic; attribute dont_touch of WX2835: signal is true;
	signal WX2836: std_logic; attribute dont_touch of WX2836: signal is true;
	signal WX2837: std_logic; attribute dont_touch of WX2837: signal is true;
	signal WX2838: std_logic; attribute dont_touch of WX2838: signal is true;
	signal WX2839: std_logic; attribute dont_touch of WX2839: signal is true;
	signal WX2840: std_logic; attribute dont_touch of WX2840: signal is true;
	signal WX2841: std_logic; attribute dont_touch of WX2841: signal is true;
	signal WX2842: std_logic; attribute dont_touch of WX2842: signal is true;
	signal WX2843: std_logic; attribute dont_touch of WX2843: signal is true;
	signal WX2844: std_logic; attribute dont_touch of WX2844: signal is true;
	signal WX2845: std_logic; attribute dont_touch of WX2845: signal is true;
	signal WX2846: std_logic; attribute dont_touch of WX2846: signal is true;
	signal WX2847: std_logic; attribute dont_touch of WX2847: signal is true;
	signal WX2848: std_logic; attribute dont_touch of WX2848: signal is true;
	signal WX2849: std_logic; attribute dont_touch of WX2849: signal is true;
	signal WX2850: std_logic; attribute dont_touch of WX2850: signal is true;
	signal WX2851: std_logic; attribute dont_touch of WX2851: signal is true;
	signal WX2852: std_logic; attribute dont_touch of WX2852: signal is true;
	signal WX2853: std_logic; attribute dont_touch of WX2853: signal is true;
	signal WX2854: std_logic; attribute dont_touch of WX2854: signal is true;
	signal WX2855: std_logic; attribute dont_touch of WX2855: signal is true;
	signal WX2856: std_logic; attribute dont_touch of WX2856: signal is true;
	signal WX2857: std_logic; attribute dont_touch of WX2857: signal is true;
	signal WX2858: std_logic; attribute dont_touch of WX2858: signal is true;
	signal WX2859: std_logic; attribute dont_touch of WX2859: signal is true;
	signal WX2860: std_logic; attribute dont_touch of WX2860: signal is true;
	signal WX2861: std_logic; attribute dont_touch of WX2861: signal is true;
	signal WX2862: std_logic; attribute dont_touch of WX2862: signal is true;
	signal WX2863: std_logic; attribute dont_touch of WX2863: signal is true;
	signal WX2864: std_logic; attribute dont_touch of WX2864: signal is true;
	signal WX2865: std_logic; attribute dont_touch of WX2865: signal is true;
	signal WX2866: std_logic; attribute dont_touch of WX2866: signal is true;
	signal WX2867: std_logic; attribute dont_touch of WX2867: signal is true;
	signal WX2868: std_logic; attribute dont_touch of WX2868: signal is true;
	signal WX2869: std_logic; attribute dont_touch of WX2869: signal is true;
	signal WX2870: std_logic; attribute dont_touch of WX2870: signal is true;
	signal WX2871: std_logic; attribute dont_touch of WX2871: signal is true;
	signal WX2872: std_logic; attribute dont_touch of WX2872: signal is true;
	signal WX2873: std_logic; attribute dont_touch of WX2873: signal is true;
	signal WX2874: std_logic; attribute dont_touch of WX2874: signal is true;
	signal WX2875: std_logic; attribute dont_touch of WX2875: signal is true;
	signal WX2876: std_logic; attribute dont_touch of WX2876: signal is true;
	signal WX2877: std_logic; attribute dont_touch of WX2877: signal is true;
	signal WX2878: std_logic; attribute dont_touch of WX2878: signal is true;
	signal WX2879: std_logic; attribute dont_touch of WX2879: signal is true;
	signal WX2880: std_logic; attribute dont_touch of WX2880: signal is true;
	signal WX2881: std_logic; attribute dont_touch of WX2881: signal is true;
	signal WX2882: std_logic; attribute dont_touch of WX2882: signal is true;
	signal WX2883: std_logic; attribute dont_touch of WX2883: signal is true;
	signal WX2884: std_logic; attribute dont_touch of WX2884: signal is true;
	signal WX2885: std_logic; attribute dont_touch of WX2885: signal is true;
	signal WX2886: std_logic; attribute dont_touch of WX2886: signal is true;
	signal WX2887: std_logic; attribute dont_touch of WX2887: signal is true;
	signal WX2888: std_logic; attribute dont_touch of WX2888: signal is true;
	signal WX2889: std_logic; attribute dont_touch of WX2889: signal is true;
	signal WX2890: std_logic; attribute dont_touch of WX2890: signal is true;
	signal WX2891: std_logic; attribute dont_touch of WX2891: signal is true;
	signal WX2892: std_logic; attribute dont_touch of WX2892: signal is true;
	signal WX2893: std_logic; attribute dont_touch of WX2893: signal is true;
	signal WX2894: std_logic; attribute dont_touch of WX2894: signal is true;
	signal WX2895: std_logic; attribute dont_touch of WX2895: signal is true;
	signal WX2896: std_logic; attribute dont_touch of WX2896: signal is true;
	signal WX2897: std_logic; attribute dont_touch of WX2897: signal is true;
	signal WX2898: std_logic; attribute dont_touch of WX2898: signal is true;
	signal WX2899: std_logic; attribute dont_touch of WX2899: signal is true;
	signal WX2900: std_logic; attribute dont_touch of WX2900: signal is true;
	signal WX2901: std_logic; attribute dont_touch of WX2901: signal is true;
	signal WX2902: std_logic; attribute dont_touch of WX2902: signal is true;
	signal WX2903: std_logic; attribute dont_touch of WX2903: signal is true;
	signal WX2904: std_logic; attribute dont_touch of WX2904: signal is true;
	signal WX2905: std_logic; attribute dont_touch of WX2905: signal is true;
	signal WX2906: std_logic; attribute dont_touch of WX2906: signal is true;
	signal WX2907: std_logic; attribute dont_touch of WX2907: signal is true;
	signal WX2908: std_logic; attribute dont_touch of WX2908: signal is true;
	signal WX2909: std_logic; attribute dont_touch of WX2909: signal is true;
	signal WX2910: std_logic; attribute dont_touch of WX2910: signal is true;
	signal WX2911: std_logic; attribute dont_touch of WX2911: signal is true;
	signal WX2912: std_logic; attribute dont_touch of WX2912: signal is true;
	signal WX2913: std_logic; attribute dont_touch of WX2913: signal is true;
	signal WX2914: std_logic; attribute dont_touch of WX2914: signal is true;
	signal WX2915: std_logic; attribute dont_touch of WX2915: signal is true;
	signal WX2916: std_logic; attribute dont_touch of WX2916: signal is true;
	signal WX2917: std_logic; attribute dont_touch of WX2917: signal is true;
	signal WX2918: std_logic; attribute dont_touch of WX2918: signal is true;
	signal WX2919: std_logic; attribute dont_touch of WX2919: signal is true;
	signal WX2920: std_logic; attribute dont_touch of WX2920: signal is true;
	signal WX2921: std_logic; attribute dont_touch of WX2921: signal is true;
	signal WX2922: std_logic; attribute dont_touch of WX2922: signal is true;
	signal WX2923: std_logic; attribute dont_touch of WX2923: signal is true;
	signal WX2924: std_logic; attribute dont_touch of WX2924: signal is true;
	signal WX2925: std_logic; attribute dont_touch of WX2925: signal is true;
	signal WX2926: std_logic; attribute dont_touch of WX2926: signal is true;
	signal WX2927: std_logic; attribute dont_touch of WX2927: signal is true;
	signal WX2928: std_logic; attribute dont_touch of WX2928: signal is true;
	signal WX2929: std_logic; attribute dont_touch of WX2929: signal is true;
	signal WX2930: std_logic; attribute dont_touch of WX2930: signal is true;
	signal WX2931: std_logic; attribute dont_touch of WX2931: signal is true;
	signal WX2932: std_logic; attribute dont_touch of WX2932: signal is true;
	signal WX2933: std_logic; attribute dont_touch of WX2933: signal is true;
	signal WX2934: std_logic; attribute dont_touch of WX2934: signal is true;
	signal WX2935: std_logic; attribute dont_touch of WX2935: signal is true;
	signal WX2936: std_logic; attribute dont_touch of WX2936: signal is true;
	signal WX2937: std_logic; attribute dont_touch of WX2937: signal is true;
	signal WX2938: std_logic; attribute dont_touch of WX2938: signal is true;
	signal WX2939: std_logic; attribute dont_touch of WX2939: signal is true;
	signal WX2940: std_logic; attribute dont_touch of WX2940: signal is true;
	signal WX2941: std_logic; attribute dont_touch of WX2941: signal is true;
	signal WX2942: std_logic; attribute dont_touch of WX2942: signal is true;
	signal WX2943: std_logic; attribute dont_touch of WX2943: signal is true;
	signal WX2944: std_logic; attribute dont_touch of WX2944: signal is true;
	signal WX2945: std_logic; attribute dont_touch of WX2945: signal is true;
	signal WX2946: std_logic; attribute dont_touch of WX2946: signal is true;
	signal WX2947: std_logic; attribute dont_touch of WX2947: signal is true;
	signal WX2948: std_logic; attribute dont_touch of WX2948: signal is true;
	signal WX2949: std_logic; attribute dont_touch of WX2949: signal is true;
	signal WX2950: std_logic; attribute dont_touch of WX2950: signal is true;
	signal WX2951: std_logic; attribute dont_touch of WX2951: signal is true;
	signal WX2952: std_logic; attribute dont_touch of WX2952: signal is true;
	signal WX2953: std_logic; attribute dont_touch of WX2953: signal is true;
	signal WX2954: std_logic; attribute dont_touch of WX2954: signal is true;
	signal WX2955: std_logic; attribute dont_touch of WX2955: signal is true;
	signal WX2956: std_logic; attribute dont_touch of WX2956: signal is true;
	signal WX2957: std_logic; attribute dont_touch of WX2957: signal is true;
	signal WX2958: std_logic; attribute dont_touch of WX2958: signal is true;
	signal WX2959: std_logic; attribute dont_touch of WX2959: signal is true;
	signal WX2960: std_logic; attribute dont_touch of WX2960: signal is true;
	signal WX2961: std_logic; attribute dont_touch of WX2961: signal is true;
	signal WX2962: std_logic; attribute dont_touch of WX2962: signal is true;
	signal WX2963: std_logic; attribute dont_touch of WX2963: signal is true;
	signal WX2964: std_logic; attribute dont_touch of WX2964: signal is true;
	signal WX2965: std_logic; attribute dont_touch of WX2965: signal is true;
	signal WX2966: std_logic; attribute dont_touch of WX2966: signal is true;
	signal WX2967: std_logic; attribute dont_touch of WX2967: signal is true;
	signal WX2968: std_logic; attribute dont_touch of WX2968: signal is true;
	signal WX2969: std_logic; attribute dont_touch of WX2969: signal is true;
	signal WX2970: std_logic; attribute dont_touch of WX2970: signal is true;
	signal WX2971: std_logic; attribute dont_touch of WX2971: signal is true;
	signal WX2972: std_logic; attribute dont_touch of WX2972: signal is true;
	signal WX2973: std_logic; attribute dont_touch of WX2973: signal is true;
	signal WX2974: std_logic; attribute dont_touch of WX2974: signal is true;
	signal WX2975: std_logic; attribute dont_touch of WX2975: signal is true;
	signal WX2976: std_logic; attribute dont_touch of WX2976: signal is true;
	signal WX2977: std_logic; attribute dont_touch of WX2977: signal is true;
	signal WX2978: std_logic; attribute dont_touch of WX2978: signal is true;
	signal WX2979: std_logic; attribute dont_touch of WX2979: signal is true;
	signal WX2980: std_logic; attribute dont_touch of WX2980: signal is true;
	signal WX2981: std_logic; attribute dont_touch of WX2981: signal is true;
	signal WX2982: std_logic; attribute dont_touch of WX2982: signal is true;
	signal WX2983: std_logic; attribute dont_touch of WX2983: signal is true;
	signal WX2984: std_logic; attribute dont_touch of WX2984: signal is true;
	signal WX2985: std_logic; attribute dont_touch of WX2985: signal is true;
	signal WX2986: std_logic; attribute dont_touch of WX2986: signal is true;
	signal WX2987: std_logic; attribute dont_touch of WX2987: signal is true;
	signal WX2988: std_logic; attribute dont_touch of WX2988: signal is true;
	signal WX2989: std_logic; attribute dont_touch of WX2989: signal is true;
	signal WX2990: std_logic; attribute dont_touch of WX2990: signal is true;
	signal WX2991: std_logic; attribute dont_touch of WX2991: signal is true;
	signal WX2992: std_logic; attribute dont_touch of WX2992: signal is true;
	signal WX2993: std_logic; attribute dont_touch of WX2993: signal is true;
	signal WX2994: std_logic; attribute dont_touch of WX2994: signal is true;
	signal WX2995: std_logic; attribute dont_touch of WX2995: signal is true;
	signal WX2996: std_logic; attribute dont_touch of WX2996: signal is true;
	signal WX2997: std_logic; attribute dont_touch of WX2997: signal is true;
	signal WX2998: std_logic; attribute dont_touch of WX2998: signal is true;
	signal WX2999: std_logic; attribute dont_touch of WX2999: signal is true;
	signal WX3000: std_logic; attribute dont_touch of WX3000: signal is true;
	signal WX3001: std_logic; attribute dont_touch of WX3001: signal is true;
	signal WX3002: std_logic; attribute dont_touch of WX3002: signal is true;
	signal WX3003: std_logic; attribute dont_touch of WX3003: signal is true;
	signal WX3004: std_logic; attribute dont_touch of WX3004: signal is true;
	signal WX3005: std_logic; attribute dont_touch of WX3005: signal is true;
	signal WX3006: std_logic; attribute dont_touch of WX3006: signal is true;
	signal WX3007: std_logic; attribute dont_touch of WX3007: signal is true;
	signal WX3008: std_logic; attribute dont_touch of WX3008: signal is true;
	signal WX3009: std_logic; attribute dont_touch of WX3009: signal is true;
	signal WX3010: std_logic; attribute dont_touch of WX3010: signal is true;
	signal WX3011: std_logic; attribute dont_touch of WX3011: signal is true;
	signal WX3012: std_logic; attribute dont_touch of WX3012: signal is true;
	signal WX3013: std_logic; attribute dont_touch of WX3013: signal is true;
	signal WX3014: std_logic; attribute dont_touch of WX3014: signal is true;
	signal WX3015: std_logic; attribute dont_touch of WX3015: signal is true;
	signal WX3016: std_logic; attribute dont_touch of WX3016: signal is true;
	signal WX3017: std_logic; attribute dont_touch of WX3017: signal is true;
	signal WX3018: std_logic; attribute dont_touch of WX3018: signal is true;
	signal WX3019: std_logic; attribute dont_touch of WX3019: signal is true;
	signal WX3020: std_logic; attribute dont_touch of WX3020: signal is true;
	signal WX3021: std_logic; attribute dont_touch of WX3021: signal is true;
	signal WX3022: std_logic; attribute dont_touch of WX3022: signal is true;
	signal WX3023: std_logic; attribute dont_touch of WX3023: signal is true;
	signal WX3024: std_logic; attribute dont_touch of WX3024: signal is true;
	signal WX3025: std_logic; attribute dont_touch of WX3025: signal is true;
	signal WX3026: std_logic; attribute dont_touch of WX3026: signal is true;
	signal WX3027: std_logic; attribute dont_touch of WX3027: signal is true;
	signal WX3028: std_logic; attribute dont_touch of WX3028: signal is true;
	signal WX3029: std_logic; attribute dont_touch of WX3029: signal is true;
	signal WX3030: std_logic; attribute dont_touch of WX3030: signal is true;
	signal WX3031: std_logic; attribute dont_touch of WX3031: signal is true;
	signal WX3032: std_logic; attribute dont_touch of WX3032: signal is true;
	signal WX3033: std_logic; attribute dont_touch of WX3033: signal is true;
	signal WX3034: std_logic; attribute dont_touch of WX3034: signal is true;
	signal WX3035: std_logic; attribute dont_touch of WX3035: signal is true;
	signal WX3036: std_logic; attribute dont_touch of WX3036: signal is true;
	signal WX3037: std_logic; attribute dont_touch of WX3037: signal is true;
	signal WX3038: std_logic; attribute dont_touch of WX3038: signal is true;
	signal WX3039: std_logic; attribute dont_touch of WX3039: signal is true;
	signal WX3040: std_logic; attribute dont_touch of WX3040: signal is true;
	signal WX3041: std_logic; attribute dont_touch of WX3041: signal is true;
	signal WX3042: std_logic; attribute dont_touch of WX3042: signal is true;
	signal WX3043: std_logic; attribute dont_touch of WX3043: signal is true;
	signal WX3044: std_logic; attribute dont_touch of WX3044: signal is true;
	signal WX3045: std_logic; attribute dont_touch of WX3045: signal is true;
	signal WX3046: std_logic; attribute dont_touch of WX3046: signal is true;
	signal WX3047: std_logic; attribute dont_touch of WX3047: signal is true;
	signal WX3048: std_logic; attribute dont_touch of WX3048: signal is true;
	signal WX3049: std_logic; attribute dont_touch of WX3049: signal is true;
	signal WX3050: std_logic; attribute dont_touch of WX3050: signal is true;
	signal WX3051: std_logic; attribute dont_touch of WX3051: signal is true;
	signal WX3052: std_logic; attribute dont_touch of WX3052: signal is true;
	signal WX3053: std_logic; attribute dont_touch of WX3053: signal is true;
	signal WX3054: std_logic; attribute dont_touch of WX3054: signal is true;
	signal WX3055: std_logic; attribute dont_touch of WX3055: signal is true;
	signal WX3056: std_logic; attribute dont_touch of WX3056: signal is true;
	signal WX3057: std_logic; attribute dont_touch of WX3057: signal is true;
	signal WX3058: std_logic; attribute dont_touch of WX3058: signal is true;
	signal WX3059: std_logic; attribute dont_touch of WX3059: signal is true;
	signal WX3060: std_logic; attribute dont_touch of WX3060: signal is true;
	signal WX3061: std_logic; attribute dont_touch of WX3061: signal is true;
	signal WX3062: std_logic; attribute dont_touch of WX3062: signal is true;
	signal WX3063: std_logic; attribute dont_touch of WX3063: signal is true;
	signal WX3064: std_logic; attribute dont_touch of WX3064: signal is true;
	signal WX3065: std_logic; attribute dont_touch of WX3065: signal is true;
	signal WX3066: std_logic; attribute dont_touch of WX3066: signal is true;
	signal WX3067: std_logic; attribute dont_touch of WX3067: signal is true;
	signal WX3068: std_logic; attribute dont_touch of WX3068: signal is true;
	signal WX3069: std_logic; attribute dont_touch of WX3069: signal is true;
	signal WX3070: std_logic; attribute dont_touch of WX3070: signal is true;
	signal WX3071: std_logic; attribute dont_touch of WX3071: signal is true;
	signal WX3072: std_logic; attribute dont_touch of WX3072: signal is true;
	signal WX3073: std_logic; attribute dont_touch of WX3073: signal is true;
	signal WX3074: std_logic; attribute dont_touch of WX3074: signal is true;
	signal WX3075: std_logic; attribute dont_touch of WX3075: signal is true;
	signal WX3076: std_logic; attribute dont_touch of WX3076: signal is true;
	signal WX3077: std_logic; attribute dont_touch of WX3077: signal is true;
	signal WX3078: std_logic; attribute dont_touch of WX3078: signal is true;
	signal WX3079: std_logic; attribute dont_touch of WX3079: signal is true;
	signal WX3080: std_logic; attribute dont_touch of WX3080: signal is true;
	signal WX3081: std_logic; attribute dont_touch of WX3081: signal is true;
	signal WX3082: std_logic; attribute dont_touch of WX3082: signal is true;
	signal WX3083: std_logic; attribute dont_touch of WX3083: signal is true;
	signal WX3084: std_logic; attribute dont_touch of WX3084: signal is true;
	signal WX3085: std_logic; attribute dont_touch of WX3085: signal is true;
	signal WX3086: std_logic; attribute dont_touch of WX3086: signal is true;
	signal WX3087: std_logic; attribute dont_touch of WX3087: signal is true;
	signal WX3088: std_logic; attribute dont_touch of WX3088: signal is true;
	signal WX3089: std_logic; attribute dont_touch of WX3089: signal is true;
	signal WX3090: std_logic; attribute dont_touch of WX3090: signal is true;
	signal WX3091: std_logic; attribute dont_touch of WX3091: signal is true;
	signal WX3092: std_logic; attribute dont_touch of WX3092: signal is true;
	signal WX3093: std_logic; attribute dont_touch of WX3093: signal is true;
	signal WX3094: std_logic; attribute dont_touch of WX3094: signal is true;
	signal WX3095: std_logic; attribute dont_touch of WX3095: signal is true;
	signal WX3096: std_logic; attribute dont_touch of WX3096: signal is true;
	signal WX3097: std_logic; attribute dont_touch of WX3097: signal is true;
	signal WX3098: std_logic; attribute dont_touch of WX3098: signal is true;
	signal WX3099: std_logic; attribute dont_touch of WX3099: signal is true;
	signal WX3100: std_logic; attribute dont_touch of WX3100: signal is true;
	signal WX3101: std_logic; attribute dont_touch of WX3101: signal is true;
	signal WX3102: std_logic; attribute dont_touch of WX3102: signal is true;
	signal WX3103: std_logic; attribute dont_touch of WX3103: signal is true;
	signal WX3104: std_logic; attribute dont_touch of WX3104: signal is true;
	signal WX3105: std_logic; attribute dont_touch of WX3105: signal is true;
	signal WX3106: std_logic; attribute dont_touch of WX3106: signal is true;
	signal WX3107: std_logic; attribute dont_touch of WX3107: signal is true;
	signal WX3108: std_logic; attribute dont_touch of WX3108: signal is true;
	signal WX3109: std_logic; attribute dont_touch of WX3109: signal is true;
	signal WX3110: std_logic; attribute dont_touch of WX3110: signal is true;
	signal WX3111: std_logic; attribute dont_touch of WX3111: signal is true;
	signal WX3112: std_logic; attribute dont_touch of WX3112: signal is true;
	signal WX3113: std_logic; attribute dont_touch of WX3113: signal is true;
	signal WX3114: std_logic; attribute dont_touch of WX3114: signal is true;
	signal WX3115: std_logic; attribute dont_touch of WX3115: signal is true;
	signal WX3116: std_logic; attribute dont_touch of WX3116: signal is true;
	signal WX3117: std_logic; attribute dont_touch of WX3117: signal is true;
	signal WX3118: std_logic; attribute dont_touch of WX3118: signal is true;
	signal WX3119: std_logic; attribute dont_touch of WX3119: signal is true;
	signal WX3120: std_logic; attribute dont_touch of WX3120: signal is true;
	signal WX3121: std_logic; attribute dont_touch of WX3121: signal is true;
	signal WX3122: std_logic; attribute dont_touch of WX3122: signal is true;
	signal WX3123: std_logic; attribute dont_touch of WX3123: signal is true;
	signal WX3124: std_logic; attribute dont_touch of WX3124: signal is true;
	signal WX3125: std_logic; attribute dont_touch of WX3125: signal is true;
	signal WX3126: std_logic; attribute dont_touch of WX3126: signal is true;
	signal WX3127: std_logic; attribute dont_touch of WX3127: signal is true;
	signal WX3128: std_logic; attribute dont_touch of WX3128: signal is true;
	signal WX3129: std_logic; attribute dont_touch of WX3129: signal is true;
	signal WX3130: std_logic; attribute dont_touch of WX3130: signal is true;
	signal WX3131: std_logic; attribute dont_touch of WX3131: signal is true;
	signal WX3132: std_logic; attribute dont_touch of WX3132: signal is true;
	signal WX3133: std_logic; attribute dont_touch of WX3133: signal is true;
	signal WX3134: std_logic; attribute dont_touch of WX3134: signal is true;
	signal WX3135: std_logic; attribute dont_touch of WX3135: signal is true;
	signal WX3136: std_logic; attribute dont_touch of WX3136: signal is true;
	signal WX3137: std_logic; attribute dont_touch of WX3137: signal is true;
	signal WX3138: std_logic; attribute dont_touch of WX3138: signal is true;
	signal WX3139: std_logic; attribute dont_touch of WX3139: signal is true;
	signal WX3140: std_logic; attribute dont_touch of WX3140: signal is true;
	signal WX3141: std_logic; attribute dont_touch of WX3141: signal is true;
	signal WX3142: std_logic; attribute dont_touch of WX3142: signal is true;
	signal WX3143: std_logic; attribute dont_touch of WX3143: signal is true;
	signal WX3144: std_logic; attribute dont_touch of WX3144: signal is true;
	signal WX3145: std_logic; attribute dont_touch of WX3145: signal is true;
	signal WX3146: std_logic; attribute dont_touch of WX3146: signal is true;
	signal WX3147: std_logic; attribute dont_touch of WX3147: signal is true;
	signal WX3148: std_logic; attribute dont_touch of WX3148: signal is true;
	signal WX3149: std_logic; attribute dont_touch of WX3149: signal is true;
	signal WX3150: std_logic; attribute dont_touch of WX3150: signal is true;
	signal WX3151: std_logic; attribute dont_touch of WX3151: signal is true;
	signal WX3152: std_logic; attribute dont_touch of WX3152: signal is true;
	signal WX3153: std_logic; attribute dont_touch of WX3153: signal is true;
	signal WX3154: std_logic; attribute dont_touch of WX3154: signal is true;
	signal WX3155: std_logic; attribute dont_touch of WX3155: signal is true;
	signal WX3156: std_logic; attribute dont_touch of WX3156: signal is true;
	signal WX3157: std_logic; attribute dont_touch of WX3157: signal is true;
	signal WX3158: std_logic; attribute dont_touch of WX3158: signal is true;
	signal WX3159: std_logic; attribute dont_touch of WX3159: signal is true;
	signal WX3160: std_logic; attribute dont_touch of WX3160: signal is true;
	signal WX3161: std_logic; attribute dont_touch of WX3161: signal is true;
	signal WX3162: std_logic; attribute dont_touch of WX3162: signal is true;
	signal WX3163: std_logic; attribute dont_touch of WX3163: signal is true;
	signal WX3164: std_logic; attribute dont_touch of WX3164: signal is true;
	signal WX3165: std_logic; attribute dont_touch of WX3165: signal is true;
	signal WX3166: std_logic; attribute dont_touch of WX3166: signal is true;
	signal WX3167: std_logic; attribute dont_touch of WX3167: signal is true;
	signal WX3168: std_logic; attribute dont_touch of WX3168: signal is true;
	signal WX3169: std_logic; attribute dont_touch of WX3169: signal is true;
	signal WX3170: std_logic; attribute dont_touch of WX3170: signal is true;
	signal WX3171: std_logic; attribute dont_touch of WX3171: signal is true;
	signal WX3172: std_logic; attribute dont_touch of WX3172: signal is true;
	signal WX3173: std_logic; attribute dont_touch of WX3173: signal is true;
	signal WX3174: std_logic; attribute dont_touch of WX3174: signal is true;
	signal WX3175: std_logic; attribute dont_touch of WX3175: signal is true;
	signal WX3176: std_logic; attribute dont_touch of WX3176: signal is true;
	signal WX3177: std_logic; attribute dont_touch of WX3177: signal is true;
	signal WX3178: std_logic; attribute dont_touch of WX3178: signal is true;
	signal WX3179: std_logic; attribute dont_touch of WX3179: signal is true;
	signal WX3180: std_logic; attribute dont_touch of WX3180: signal is true;
	signal WX3181: std_logic; attribute dont_touch of WX3181: signal is true;
	signal WX3182: std_logic; attribute dont_touch of WX3182: signal is true;
	signal WX3183: std_logic; attribute dont_touch of WX3183: signal is true;
	signal WX3184: std_logic; attribute dont_touch of WX3184: signal is true;
	signal WX3185: std_logic; attribute dont_touch of WX3185: signal is true;
	signal WX3186: std_logic; attribute dont_touch of WX3186: signal is true;
	signal WX3187: std_logic; attribute dont_touch of WX3187: signal is true;
	signal WX3188: std_logic; attribute dont_touch of WX3188: signal is true;
	signal WX3189: std_logic; attribute dont_touch of WX3189: signal is true;
	signal WX3190: std_logic; attribute dont_touch of WX3190: signal is true;
	signal WX3191: std_logic; attribute dont_touch of WX3191: signal is true;
	signal WX3192: std_logic; attribute dont_touch of WX3192: signal is true;
	signal WX3193: std_logic; attribute dont_touch of WX3193: signal is true;
	signal WX3194: std_logic; attribute dont_touch of WX3194: signal is true;
	signal WX3195: std_logic; attribute dont_touch of WX3195: signal is true;
	signal WX3196: std_logic; attribute dont_touch of WX3196: signal is true;
	signal WX3197: std_logic; attribute dont_touch of WX3197: signal is true;
	signal WX3198: std_logic; attribute dont_touch of WX3198: signal is true;
	signal WX3199: std_logic; attribute dont_touch of WX3199: signal is true;
	signal WX3200: std_logic; attribute dont_touch of WX3200: signal is true;
	signal WX3201: std_logic; attribute dont_touch of WX3201: signal is true;
	signal WX3202: std_logic; attribute dont_touch of WX3202: signal is true;
	signal WX3203: std_logic; attribute dont_touch of WX3203: signal is true;
	signal WX3204: std_logic; attribute dont_touch of WX3204: signal is true;
	signal WX3205: std_logic; attribute dont_touch of WX3205: signal is true;
	signal WX3206: std_logic; attribute dont_touch of WX3206: signal is true;
	signal WX3207: std_logic; attribute dont_touch of WX3207: signal is true;
	signal WX3208: std_logic; attribute dont_touch of WX3208: signal is true;
	signal WX3209: std_logic; attribute dont_touch of WX3209: signal is true;
	signal WX3210: std_logic; attribute dont_touch of WX3210: signal is true;
	signal WX3211: std_logic; attribute dont_touch of WX3211: signal is true;
	signal WX3212: std_logic; attribute dont_touch of WX3212: signal is true;
	signal WX3213: std_logic; attribute dont_touch of WX3213: signal is true;
	signal WX3214: std_logic; attribute dont_touch of WX3214: signal is true;
	signal WX3215: std_logic; attribute dont_touch of WX3215: signal is true;
	signal WX3216: std_logic; attribute dont_touch of WX3216: signal is true;
	signal WX3217: std_logic; attribute dont_touch of WX3217: signal is true;
	signal WX3218: std_logic; attribute dont_touch of WX3218: signal is true;
	signal WX3219: std_logic; attribute dont_touch of WX3219: signal is true;
	signal WX3220: std_logic; attribute dont_touch of WX3220: signal is true;
	signal WX3221: std_logic; attribute dont_touch of WX3221: signal is true;
	signal WX3222: std_logic; attribute dont_touch of WX3222: signal is true;
	signal WX3223: std_logic; attribute dont_touch of WX3223: signal is true;
	signal WX3224: std_logic; attribute dont_touch of WX3224: signal is true;
	signal WX3225: std_logic; attribute dont_touch of WX3225: signal is true;
	signal WX3226: std_logic; attribute dont_touch of WX3226: signal is true;
	signal WX3227: std_logic; attribute dont_touch of WX3227: signal is true;
	signal WX3228: std_logic; attribute dont_touch of WX3228: signal is true;
	signal WX3229: std_logic; attribute dont_touch of WX3229: signal is true;
	signal WX3230: std_logic; attribute dont_touch of WX3230: signal is true;
	signal WX3231: std_logic; attribute dont_touch of WX3231: signal is true;
	signal WX3232: std_logic; attribute dont_touch of WX3232: signal is true;
	signal WX3233: std_logic; attribute dont_touch of WX3233: signal is true;
	signal WX3234: std_logic; attribute dont_touch of WX3234: signal is true;
	signal WX3235: std_logic; attribute dont_touch of WX3235: signal is true;
	signal WX3236: std_logic; attribute dont_touch of WX3236: signal is true;
	signal WX3237: std_logic; attribute dont_touch of WX3237: signal is true;
	signal WX3238: std_logic; attribute dont_touch of WX3238: signal is true;
	signal WX3239: std_logic; attribute dont_touch of WX3239: signal is true;
	signal WX3240: std_logic; attribute dont_touch of WX3240: signal is true;
	signal WX3241: std_logic; attribute dont_touch of WX3241: signal is true;
	signal WX3242: std_logic; attribute dont_touch of WX3242: signal is true;
	signal WX3243: std_logic; attribute dont_touch of WX3243: signal is true;
	signal WX3244: std_logic; attribute dont_touch of WX3244: signal is true;
	signal WX3245: std_logic; attribute dont_touch of WX3245: signal is true;
	signal WX3246: std_logic; attribute dont_touch of WX3246: signal is true;
	signal WX3247: std_logic; attribute dont_touch of WX3247: signal is true;
	signal WX3248: std_logic; attribute dont_touch of WX3248: signal is true;
	signal WX3249: std_logic; attribute dont_touch of WX3249: signal is true;
	signal WX3250: std_logic; attribute dont_touch of WX3250: signal is true;
	signal WX3251: std_logic; attribute dont_touch of WX3251: signal is true;
	signal WX3252: std_logic; attribute dont_touch of WX3252: signal is true;
	signal WX3253: std_logic; attribute dont_touch of WX3253: signal is true;
	signal WX3254: std_logic; attribute dont_touch of WX3254: signal is true;
	signal WX3255: std_logic; attribute dont_touch of WX3255: signal is true;
	signal WX3256: std_logic; attribute dont_touch of WX3256: signal is true;
	signal WX3257: std_logic; attribute dont_touch of WX3257: signal is true;
	signal WX3258: std_logic; attribute dont_touch of WX3258: signal is true;
	signal WX3259: std_logic; attribute dont_touch of WX3259: signal is true;
	signal WX3260: std_logic; attribute dont_touch of WX3260: signal is true;
	signal WX3261: std_logic; attribute dont_touch of WX3261: signal is true;
	signal WX3262: std_logic; attribute dont_touch of WX3262: signal is true;
	signal WX3263: std_logic; attribute dont_touch of WX3263: signal is true;
	signal WX3264: std_logic; attribute dont_touch of WX3264: signal is true;
	signal WX3265: std_logic; attribute dont_touch of WX3265: signal is true;
	signal WX3266: std_logic; attribute dont_touch of WX3266: signal is true;
	signal WX3267: std_logic; attribute dont_touch of WX3267: signal is true;
	signal WX3268: std_logic; attribute dont_touch of WX3268: signal is true;
	signal WX3269: std_logic; attribute dont_touch of WX3269: signal is true;
	signal WX3270: std_logic; attribute dont_touch of WX3270: signal is true;
	signal WX3271: std_logic; attribute dont_touch of WX3271: signal is true;
	signal WX3272: std_logic; attribute dont_touch of WX3272: signal is true;
	signal WX3273: std_logic; attribute dont_touch of WX3273: signal is true;
	signal WX3274: std_logic; attribute dont_touch of WX3274: signal is true;
	signal WX3275: std_logic; attribute dont_touch of WX3275: signal is true;
	signal WX3276: std_logic; attribute dont_touch of WX3276: signal is true;
	signal WX3277: std_logic; attribute dont_touch of WX3277: signal is true;
	signal WX3278: std_logic; attribute dont_touch of WX3278: signal is true;
	signal WX3279: std_logic; attribute dont_touch of WX3279: signal is true;
	signal WX3280: std_logic; attribute dont_touch of WX3280: signal is true;
	signal WX3281: std_logic; attribute dont_touch of WX3281: signal is true;
	signal WX3282: std_logic; attribute dont_touch of WX3282: signal is true;
	signal WX3283: std_logic; attribute dont_touch of WX3283: signal is true;
	signal WX3284: std_logic; attribute dont_touch of WX3284: signal is true;
	signal WX3285: std_logic; attribute dont_touch of WX3285: signal is true;
	signal WX3286: std_logic; attribute dont_touch of WX3286: signal is true;
	signal WX3287: std_logic; attribute dont_touch of WX3287: signal is true;
	signal WX3288: std_logic; attribute dont_touch of WX3288: signal is true;
	signal WX3289: std_logic; attribute dont_touch of WX3289: signal is true;
	signal WX3290: std_logic; attribute dont_touch of WX3290: signal is true;
	signal WX3291: std_logic; attribute dont_touch of WX3291: signal is true;
	signal WX3292: std_logic; attribute dont_touch of WX3292: signal is true;
	signal WX3293: std_logic; attribute dont_touch of WX3293: signal is true;
	signal WX3294: std_logic; attribute dont_touch of WX3294: signal is true;
	signal WX3295: std_logic; attribute dont_touch of WX3295: signal is true;
	signal WX3296: std_logic; attribute dont_touch of WX3296: signal is true;
	signal WX3297: std_logic; attribute dont_touch of WX3297: signal is true;
	signal WX3298: std_logic; attribute dont_touch of WX3298: signal is true;
	signal WX3299: std_logic; attribute dont_touch of WX3299: signal is true;
	signal WX3300: std_logic; attribute dont_touch of WX3300: signal is true;
	signal WX3301: std_logic; attribute dont_touch of WX3301: signal is true;
	signal WX3302: std_logic; attribute dont_touch of WX3302: signal is true;
	signal WX3303: std_logic; attribute dont_touch of WX3303: signal is true;
	signal WX3304: std_logic; attribute dont_touch of WX3304: signal is true;
	signal WX3305: std_logic; attribute dont_touch of WX3305: signal is true;
	signal WX3306: std_logic; attribute dont_touch of WX3306: signal is true;
	signal WX3307: std_logic; attribute dont_touch of WX3307: signal is true;
	signal WX3308: std_logic; attribute dont_touch of WX3308: signal is true;
	signal WX3309: std_logic; attribute dont_touch of WX3309: signal is true;
	signal WX3310: std_logic; attribute dont_touch of WX3310: signal is true;
	signal WX3311: std_logic; attribute dont_touch of WX3311: signal is true;
	signal WX3312: std_logic; attribute dont_touch of WX3312: signal is true;
	signal WX3313: std_logic; attribute dont_touch of WX3313: signal is true;
	signal WX3314: std_logic; attribute dont_touch of WX3314: signal is true;
	signal WX3315: std_logic; attribute dont_touch of WX3315: signal is true;
	signal WX3316: std_logic; attribute dont_touch of WX3316: signal is true;
	signal WX3317: std_logic; attribute dont_touch of WX3317: signal is true;
	signal WX3318: std_logic; attribute dont_touch of WX3318: signal is true;
	signal WX3319: std_logic; attribute dont_touch of WX3319: signal is true;
	signal WX3320: std_logic; attribute dont_touch of WX3320: signal is true;
	signal WX3321: std_logic; attribute dont_touch of WX3321: signal is true;
	signal WX3322: std_logic; attribute dont_touch of WX3322: signal is true;
	signal WX3323: std_logic; attribute dont_touch of WX3323: signal is true;
	signal WX3324: std_logic; attribute dont_touch of WX3324: signal is true;
	signal WX3325: std_logic; attribute dont_touch of WX3325: signal is true;
	signal WX3326: std_logic; attribute dont_touch of WX3326: signal is true;
	signal WX3327: std_logic; attribute dont_touch of WX3327: signal is true;
	signal WX3328: std_logic; attribute dont_touch of WX3328: signal is true;
	signal WX3329: std_logic; attribute dont_touch of WX3329: signal is true;
	signal WX3330: std_logic; attribute dont_touch of WX3330: signal is true;
	signal WX3331: std_logic; attribute dont_touch of WX3331: signal is true;
	signal WX3332: std_logic; attribute dont_touch of WX3332: signal is true;
	signal WX3333: std_logic; attribute dont_touch of WX3333: signal is true;
	signal WX3334: std_logic; attribute dont_touch of WX3334: signal is true;
	signal WX3335: std_logic; attribute dont_touch of WX3335: signal is true;
	signal WX3336: std_logic; attribute dont_touch of WX3336: signal is true;
	signal WX3337: std_logic; attribute dont_touch of WX3337: signal is true;
	signal WX3338: std_logic; attribute dont_touch of WX3338: signal is true;
	signal WX3339: std_logic; attribute dont_touch of WX3339: signal is true;
	signal WX3340: std_logic; attribute dont_touch of WX3340: signal is true;
	signal WX3341: std_logic; attribute dont_touch of WX3341: signal is true;
	signal WX3342: std_logic; attribute dont_touch of WX3342: signal is true;
	signal WX3343: std_logic; attribute dont_touch of WX3343: signal is true;
	signal WX3344: std_logic; attribute dont_touch of WX3344: signal is true;
	signal WX3345: std_logic; attribute dont_touch of WX3345: signal is true;
	signal WX3346: std_logic; attribute dont_touch of WX3346: signal is true;
	signal WX3347: std_logic; attribute dont_touch of WX3347: signal is true;
	signal WX3348: std_logic; attribute dont_touch of WX3348: signal is true;
	signal WX3349: std_logic; attribute dont_touch of WX3349: signal is true;
	signal WX3350: std_logic; attribute dont_touch of WX3350: signal is true;
	signal WX3351: std_logic; attribute dont_touch of WX3351: signal is true;
	signal WX3352: std_logic; attribute dont_touch of WX3352: signal is true;
	signal WX3353: std_logic; attribute dont_touch of WX3353: signal is true;
	signal WX3354: std_logic; attribute dont_touch of WX3354: signal is true;
	signal WX3355: std_logic; attribute dont_touch of WX3355: signal is true;
	signal WX3356: std_logic; attribute dont_touch of WX3356: signal is true;
	signal WX3357: std_logic; attribute dont_touch of WX3357: signal is true;
	signal WX3358: std_logic; attribute dont_touch of WX3358: signal is true;
	signal WX3359: std_logic; attribute dont_touch of WX3359: signal is true;
	signal WX3360: std_logic; attribute dont_touch of WX3360: signal is true;
	signal WX3361: std_logic; attribute dont_touch of WX3361: signal is true;
	signal WX3362: std_logic; attribute dont_touch of WX3362: signal is true;
	signal WX3363: std_logic; attribute dont_touch of WX3363: signal is true;
	signal WX3364: std_logic; attribute dont_touch of WX3364: signal is true;
	signal WX3365: std_logic; attribute dont_touch of WX3365: signal is true;
	signal WX3366: std_logic; attribute dont_touch of WX3366: signal is true;
	signal WX3367: std_logic; attribute dont_touch of WX3367: signal is true;
	signal WX3368: std_logic; attribute dont_touch of WX3368: signal is true;
	signal WX3369: std_logic; attribute dont_touch of WX3369: signal is true;
	signal WX3370: std_logic; attribute dont_touch of WX3370: signal is true;
	signal WX3371: std_logic; attribute dont_touch of WX3371: signal is true;
	signal WX3372: std_logic; attribute dont_touch of WX3372: signal is true;
	signal WX3373: std_logic; attribute dont_touch of WX3373: signal is true;
	signal WX3374: std_logic; attribute dont_touch of WX3374: signal is true;
	signal WX3375: std_logic; attribute dont_touch of WX3375: signal is true;
	signal WX3376: std_logic; attribute dont_touch of WX3376: signal is true;
	signal WX3377: std_logic; attribute dont_touch of WX3377: signal is true;
	signal WX3378: std_logic; attribute dont_touch of WX3378: signal is true;
	signal WX3379: std_logic; attribute dont_touch of WX3379: signal is true;
	signal WX3380: std_logic; attribute dont_touch of WX3380: signal is true;
	signal WX3381: std_logic; attribute dont_touch of WX3381: signal is true;
	signal WX3382: std_logic; attribute dont_touch of WX3382: signal is true;
	signal WX3383: std_logic; attribute dont_touch of WX3383: signal is true;
	signal WX3384: std_logic; attribute dont_touch of WX3384: signal is true;
	signal WX3385: std_logic; attribute dont_touch of WX3385: signal is true;
	signal WX3386: std_logic; attribute dont_touch of WX3386: signal is true;
	signal WX3387: std_logic; attribute dont_touch of WX3387: signal is true;
	signal WX3388: std_logic; attribute dont_touch of WX3388: signal is true;
	signal WX3389: std_logic; attribute dont_touch of WX3389: signal is true;
	signal WX3390: std_logic; attribute dont_touch of WX3390: signal is true;
	signal WX3391: std_logic; attribute dont_touch of WX3391: signal is true;
	signal WX3392: std_logic; attribute dont_touch of WX3392: signal is true;
	signal WX3393: std_logic; attribute dont_touch of WX3393: signal is true;
	signal WX3394: std_logic; attribute dont_touch of WX3394: signal is true;
	signal WX3395: std_logic; attribute dont_touch of WX3395: signal is true;
	signal WX3396: std_logic; attribute dont_touch of WX3396: signal is true;
	signal WX3397: std_logic; attribute dont_touch of WX3397: signal is true;
	signal WX3398: std_logic; attribute dont_touch of WX3398: signal is true;
	signal WX3399: std_logic; attribute dont_touch of WX3399: signal is true;
	signal WX3400: std_logic; attribute dont_touch of WX3400: signal is true;
	signal WX3401: std_logic; attribute dont_touch of WX3401: signal is true;
	signal WX3402: std_logic; attribute dont_touch of WX3402: signal is true;
	signal WX3403: std_logic; attribute dont_touch of WX3403: signal is true;
	signal WX3404: std_logic; attribute dont_touch of WX3404: signal is true;
	signal WX3405: std_logic; attribute dont_touch of WX3405: signal is true;
	signal WX3406: std_logic; attribute dont_touch of WX3406: signal is true;
	signal WX3407: std_logic; attribute dont_touch of WX3407: signal is true;
	signal WX3408: std_logic; attribute dont_touch of WX3408: signal is true;
	signal WX3409: std_logic; attribute dont_touch of WX3409: signal is true;
	signal WX3410: std_logic; attribute dont_touch of WX3410: signal is true;
	signal WX3411: std_logic; attribute dont_touch of WX3411: signal is true;
	signal WX3412: std_logic; attribute dont_touch of WX3412: signal is true;
	signal WX3413: std_logic; attribute dont_touch of WX3413: signal is true;
	signal WX3414: std_logic; attribute dont_touch of WX3414: signal is true;
	signal WX3415: std_logic; attribute dont_touch of WX3415: signal is true;
	signal WX3416: std_logic; attribute dont_touch of WX3416: signal is true;
	signal WX3417: std_logic; attribute dont_touch of WX3417: signal is true;
	signal WX3418: std_logic; attribute dont_touch of WX3418: signal is true;
	signal WX3419: std_logic; attribute dont_touch of WX3419: signal is true;
	signal WX3420: std_logic; attribute dont_touch of WX3420: signal is true;
	signal WX3421: std_logic; attribute dont_touch of WX3421: signal is true;
	signal WX3422: std_logic; attribute dont_touch of WX3422: signal is true;
	signal WX3423: std_logic; attribute dont_touch of WX3423: signal is true;
	signal WX3424: std_logic; attribute dont_touch of WX3424: signal is true;
	signal WX3425: std_logic; attribute dont_touch of WX3425: signal is true;
	signal WX3426: std_logic; attribute dont_touch of WX3426: signal is true;
	signal WX3427: std_logic; attribute dont_touch of WX3427: signal is true;
	signal WX3428: std_logic; attribute dont_touch of WX3428: signal is true;
	signal WX3429: std_logic; attribute dont_touch of WX3429: signal is true;
	signal WX3430: std_logic; attribute dont_touch of WX3430: signal is true;
	signal WX3431: std_logic; attribute dont_touch of WX3431: signal is true;
	signal WX3432: std_logic; attribute dont_touch of WX3432: signal is true;
	signal WX3433: std_logic; attribute dont_touch of WX3433: signal is true;
	signal WX3434: std_logic; attribute dont_touch of WX3434: signal is true;
	signal WX3435: std_logic; attribute dont_touch of WX3435: signal is true;
	signal WX3436: std_logic; attribute dont_touch of WX3436: signal is true;
	signal WX3437: std_logic; attribute dont_touch of WX3437: signal is true;
	signal WX3438: std_logic; attribute dont_touch of WX3438: signal is true;
	signal WX3439: std_logic; attribute dont_touch of WX3439: signal is true;
	signal WX3440: std_logic; attribute dont_touch of WX3440: signal is true;
	signal WX3441: std_logic; attribute dont_touch of WX3441: signal is true;
	signal WX3442: std_logic; attribute dont_touch of WX3442: signal is true;
	signal WX3443: std_logic; attribute dont_touch of WX3443: signal is true;
	signal WX3444: std_logic; attribute dont_touch of WX3444: signal is true;
	signal WX3445: std_logic; attribute dont_touch of WX3445: signal is true;
	signal WX3446: std_logic; attribute dont_touch of WX3446: signal is true;
	signal WX3447: std_logic; attribute dont_touch of WX3447: signal is true;
	signal WX3448: std_logic; attribute dont_touch of WX3448: signal is true;
	signal WX3449: std_logic; attribute dont_touch of WX3449: signal is true;
	signal WX3450: std_logic; attribute dont_touch of WX3450: signal is true;
	signal WX3451: std_logic; attribute dont_touch of WX3451: signal is true;
	signal WX3452: std_logic; attribute dont_touch of WX3452: signal is true;
	signal WX3453: std_logic; attribute dont_touch of WX3453: signal is true;
	signal WX3454: std_logic; attribute dont_touch of WX3454: signal is true;
	signal WX3455: std_logic; attribute dont_touch of WX3455: signal is true;
	signal WX3456: std_logic; attribute dont_touch of WX3456: signal is true;
	signal WX3457: std_logic; attribute dont_touch of WX3457: signal is true;
	signal WX3458: std_logic; attribute dont_touch of WX3458: signal is true;
	signal WX3459: std_logic; attribute dont_touch of WX3459: signal is true;
	signal WX3460: std_logic; attribute dont_touch of WX3460: signal is true;
	signal WX3461: std_logic; attribute dont_touch of WX3461: signal is true;
	signal WX3462: std_logic; attribute dont_touch of WX3462: signal is true;
	signal WX3463: std_logic; attribute dont_touch of WX3463: signal is true;
	signal WX3464: std_logic; attribute dont_touch of WX3464: signal is true;
	signal WX3465: std_logic; attribute dont_touch of WX3465: signal is true;
	signal WX3466: std_logic; attribute dont_touch of WX3466: signal is true;
	signal WX3467: std_logic; attribute dont_touch of WX3467: signal is true;
	signal WX3468: std_logic; attribute dont_touch of WX3468: signal is true;
	signal WX3469: std_logic; attribute dont_touch of WX3469: signal is true;
	signal WX3470: std_logic; attribute dont_touch of WX3470: signal is true;
	signal WX3471: std_logic; attribute dont_touch of WX3471: signal is true;
	signal WX3472: std_logic; attribute dont_touch of WX3472: signal is true;
	signal WX3473: std_logic; attribute dont_touch of WX3473: signal is true;
	signal WX3474: std_logic; attribute dont_touch of WX3474: signal is true;
	signal WX3475: std_logic; attribute dont_touch of WX3475: signal is true;
	signal WX3476: std_logic; attribute dont_touch of WX3476: signal is true;
	signal WX3477: std_logic; attribute dont_touch of WX3477: signal is true;
	signal WX3478: std_logic; attribute dont_touch of WX3478: signal is true;
	signal WX3479: std_logic; attribute dont_touch of WX3479: signal is true;
	signal WX3480: std_logic; attribute dont_touch of WX3480: signal is true;
	signal WX3481: std_logic; attribute dont_touch of WX3481: signal is true;
	signal WX3482: std_logic; attribute dont_touch of WX3482: signal is true;
	signal WX3483: std_logic; attribute dont_touch of WX3483: signal is true;
	signal WX3484: std_logic; attribute dont_touch of WX3484: signal is true;
	signal WX3485: std_logic; attribute dont_touch of WX3485: signal is true;
	signal WX3486: std_logic; attribute dont_touch of WX3486: signal is true;
	signal WX3487: std_logic; attribute dont_touch of WX3487: signal is true;
	signal WX3488: std_logic; attribute dont_touch of WX3488: signal is true;
	signal WX3489: std_logic; attribute dont_touch of WX3489: signal is true;
	signal WX3490: std_logic; attribute dont_touch of WX3490: signal is true;
	signal WX3491: std_logic; attribute dont_touch of WX3491: signal is true;
	signal WX3492: std_logic; attribute dont_touch of WX3492: signal is true;
	signal WX3493: std_logic; attribute dont_touch of WX3493: signal is true;
	signal WX3494: std_logic; attribute dont_touch of WX3494: signal is true;
	signal WX3495: std_logic; attribute dont_touch of WX3495: signal is true;
	signal WX3496: std_logic; attribute dont_touch of WX3496: signal is true;
	signal WX3497: std_logic; attribute dont_touch of WX3497: signal is true;
	signal WX3498: std_logic; attribute dont_touch of WX3498: signal is true;
	signal WX3499: std_logic; attribute dont_touch of WX3499: signal is true;
	signal WX3500: std_logic; attribute dont_touch of WX3500: signal is true;
	signal WX3501: std_logic; attribute dont_touch of WX3501: signal is true;
	signal WX3502: std_logic; attribute dont_touch of WX3502: signal is true;
	signal WX3503: std_logic; attribute dont_touch of WX3503: signal is true;
	signal WX3504: std_logic; attribute dont_touch of WX3504: signal is true;
	signal WX3505: std_logic; attribute dont_touch of WX3505: signal is true;
	signal WX3506: std_logic; attribute dont_touch of WX3506: signal is true;
	signal WX3507: std_logic; attribute dont_touch of WX3507: signal is true;
	signal WX3508: std_logic; attribute dont_touch of WX3508: signal is true;
	signal WX3509: std_logic; attribute dont_touch of WX3509: signal is true;
	signal WX3510: std_logic; attribute dont_touch of WX3510: signal is true;
	signal WX3511: std_logic; attribute dont_touch of WX3511: signal is true;
	signal WX3512: std_logic; attribute dont_touch of WX3512: signal is true;
	signal WX3513: std_logic; attribute dont_touch of WX3513: signal is true;
	signal WX3514: std_logic; attribute dont_touch of WX3514: signal is true;
	signal WX3515: std_logic; attribute dont_touch of WX3515: signal is true;
	signal WX3516: std_logic; attribute dont_touch of WX3516: signal is true;
	signal WX3517: std_logic; attribute dont_touch of WX3517: signal is true;
	signal WX3518: std_logic; attribute dont_touch of WX3518: signal is true;
	signal WX3519: std_logic; attribute dont_touch of WX3519: signal is true;
	signal WX3520: std_logic; attribute dont_touch of WX3520: signal is true;
	signal WX3521: std_logic; attribute dont_touch of WX3521: signal is true;
	signal WX3522: std_logic; attribute dont_touch of WX3522: signal is true;
	signal WX3523: std_logic; attribute dont_touch of WX3523: signal is true;
	signal WX3524: std_logic; attribute dont_touch of WX3524: signal is true;
	signal WX3525: std_logic; attribute dont_touch of WX3525: signal is true;
	signal WX3526: std_logic; attribute dont_touch of WX3526: signal is true;
	signal WX3527: std_logic; attribute dont_touch of WX3527: signal is true;
	signal WX3528: std_logic; attribute dont_touch of WX3528: signal is true;
	signal WX3529: std_logic; attribute dont_touch of WX3529: signal is true;
	signal WX3530: std_logic; attribute dont_touch of WX3530: signal is true;
	signal WX3531: std_logic; attribute dont_touch of WX3531: signal is true;
	signal WX3532: std_logic; attribute dont_touch of WX3532: signal is true;
	signal WX3533: std_logic; attribute dont_touch of WX3533: signal is true;
	signal WX3534: std_logic; attribute dont_touch of WX3534: signal is true;
	signal WX3535: std_logic; attribute dont_touch of WX3535: signal is true;
	signal WX3536: std_logic; attribute dont_touch of WX3536: signal is true;
	signal WX3537: std_logic; attribute dont_touch of WX3537: signal is true;
	signal WX3538: std_logic; attribute dont_touch of WX3538: signal is true;
	signal WX3539: std_logic; attribute dont_touch of WX3539: signal is true;
	signal WX3540: std_logic; attribute dont_touch of WX3540: signal is true;
	signal WX3541: std_logic; attribute dont_touch of WX3541: signal is true;
	signal WX3542: std_logic; attribute dont_touch of WX3542: signal is true;
	signal WX3543: std_logic; attribute dont_touch of WX3543: signal is true;
	signal WX3544: std_logic; attribute dont_touch of WX3544: signal is true;
	signal WX3545: std_logic; attribute dont_touch of WX3545: signal is true;
	signal WX3546: std_logic; attribute dont_touch of WX3546: signal is true;
	signal WX3547: std_logic; attribute dont_touch of WX3547: signal is true;
	signal WX3548: std_logic; attribute dont_touch of WX3548: signal is true;
	signal WX3549: std_logic; attribute dont_touch of WX3549: signal is true;
	signal WX3550: std_logic; attribute dont_touch of WX3550: signal is true;
	signal WX3551: std_logic; attribute dont_touch of WX3551: signal is true;
	signal WX3552: std_logic; attribute dont_touch of WX3552: signal is true;
	signal WX3553: std_logic; attribute dont_touch of WX3553: signal is true;
	signal WX3554: std_logic; attribute dont_touch of WX3554: signal is true;
	signal WX3555: std_logic; attribute dont_touch of WX3555: signal is true;
	signal WX3556: std_logic; attribute dont_touch of WX3556: signal is true;
	signal WX3557: std_logic; attribute dont_touch of WX3557: signal is true;
	signal WX3558: std_logic; attribute dont_touch of WX3558: signal is true;
	signal WX3559: std_logic; attribute dont_touch of WX3559: signal is true;
	signal WX3560: std_logic; attribute dont_touch of WX3560: signal is true;
	signal WX3561: std_logic; attribute dont_touch of WX3561: signal is true;
	signal WX3562: std_logic; attribute dont_touch of WX3562: signal is true;
	signal WX3563: std_logic; attribute dont_touch of WX3563: signal is true;
	signal WX3564: std_logic; attribute dont_touch of WX3564: signal is true;
	signal WX3565: std_logic; attribute dont_touch of WX3565: signal is true;
	signal WX3566: std_logic; attribute dont_touch of WX3566: signal is true;
	signal WX3567: std_logic; attribute dont_touch of WX3567: signal is true;
	signal WX3568: std_logic; attribute dont_touch of WX3568: signal is true;
	signal WX3569: std_logic; attribute dont_touch of WX3569: signal is true;
	signal WX3570: std_logic; attribute dont_touch of WX3570: signal is true;
	signal WX3571: std_logic; attribute dont_touch of WX3571: signal is true;
	signal WX3572: std_logic; attribute dont_touch of WX3572: signal is true;
	signal WX3573: std_logic; attribute dont_touch of WX3573: signal is true;
	signal WX3574: std_logic; attribute dont_touch of WX3574: signal is true;
	signal WX3575: std_logic; attribute dont_touch of WX3575: signal is true;
	signal WX3576: std_logic; attribute dont_touch of WX3576: signal is true;
	signal WX3577: std_logic; attribute dont_touch of WX3577: signal is true;
	signal WX3578: std_logic; attribute dont_touch of WX3578: signal is true;
	signal WX3579: std_logic; attribute dont_touch of WX3579: signal is true;
	signal WX3580: std_logic; attribute dont_touch of WX3580: signal is true;
	signal WX3581: std_logic; attribute dont_touch of WX3581: signal is true;
	signal WX3582: std_logic; attribute dont_touch of WX3582: signal is true;
	signal WX3583: std_logic; attribute dont_touch of WX3583: signal is true;
	signal WX3584: std_logic; attribute dont_touch of WX3584: signal is true;
	signal WX3585: std_logic; attribute dont_touch of WX3585: signal is true;
	signal WX3586: std_logic; attribute dont_touch of WX3586: signal is true;
	signal WX3587: std_logic; attribute dont_touch of WX3587: signal is true;
	signal WX3588: std_logic; attribute dont_touch of WX3588: signal is true;
	signal WX3589: std_logic; attribute dont_touch of WX3589: signal is true;
	signal WX3590: std_logic; attribute dont_touch of WX3590: signal is true;
	signal WX3591: std_logic; attribute dont_touch of WX3591: signal is true;
	signal WX3592: std_logic; attribute dont_touch of WX3592: signal is true;
	signal WX3593: std_logic; attribute dont_touch of WX3593: signal is true;
	signal WX3594: std_logic; attribute dont_touch of WX3594: signal is true;
	signal WX3595: std_logic; attribute dont_touch of WX3595: signal is true;
	signal WX3596: std_logic; attribute dont_touch of WX3596: signal is true;
	signal WX3597: std_logic; attribute dont_touch of WX3597: signal is true;
	signal WX3598: std_logic; attribute dont_touch of WX3598: signal is true;
	signal WX3599: std_logic; attribute dont_touch of WX3599: signal is true;
	signal WX3600: std_logic; attribute dont_touch of WX3600: signal is true;
	signal WX3601: std_logic; attribute dont_touch of WX3601: signal is true;
	signal WX3602: std_logic; attribute dont_touch of WX3602: signal is true;
	signal WX3603: std_logic; attribute dont_touch of WX3603: signal is true;
	signal WX3604: std_logic; attribute dont_touch of WX3604: signal is true;
	signal WX3605: std_logic; attribute dont_touch of WX3605: signal is true;
	signal WX3606: std_logic; attribute dont_touch of WX3606: signal is true;
	signal WX3607: std_logic; attribute dont_touch of WX3607: signal is true;
	signal WX3608: std_logic; attribute dont_touch of WX3608: signal is true;
	signal WX3609: std_logic; attribute dont_touch of WX3609: signal is true;
	signal WX3610: std_logic; attribute dont_touch of WX3610: signal is true;
	signal WX3611: std_logic; attribute dont_touch of WX3611: signal is true;
	signal WX3612: std_logic; attribute dont_touch of WX3612: signal is true;
	signal WX3613: std_logic; attribute dont_touch of WX3613: signal is true;
	signal WX3614: std_logic; attribute dont_touch of WX3614: signal is true;
	signal WX3615: std_logic; attribute dont_touch of WX3615: signal is true;
	signal WX3616: std_logic; attribute dont_touch of WX3616: signal is true;
	signal WX3617: std_logic; attribute dont_touch of WX3617: signal is true;
	signal WX3618: std_logic; attribute dont_touch of WX3618: signal is true;
	signal WX3619: std_logic; attribute dont_touch of WX3619: signal is true;
	signal WX3620: std_logic; attribute dont_touch of WX3620: signal is true;
	signal WX3621: std_logic; attribute dont_touch of WX3621: signal is true;
	signal WX3622: std_logic; attribute dont_touch of WX3622: signal is true;
	signal WX3623: std_logic; attribute dont_touch of WX3623: signal is true;
	signal WX3624: std_logic; attribute dont_touch of WX3624: signal is true;
	signal WX3625: std_logic; attribute dont_touch of WX3625: signal is true;
	signal WX3626: std_logic; attribute dont_touch of WX3626: signal is true;
	signal WX3627: std_logic; attribute dont_touch of WX3627: signal is true;
	signal WX3628: std_logic; attribute dont_touch of WX3628: signal is true;
	signal WX3629: std_logic; attribute dont_touch of WX3629: signal is true;
	signal WX3630: std_logic; attribute dont_touch of WX3630: signal is true;
	signal WX3631: std_logic; attribute dont_touch of WX3631: signal is true;
	signal WX3632: std_logic; attribute dont_touch of WX3632: signal is true;
	signal WX3633: std_logic; attribute dont_touch of WX3633: signal is true;
	signal WX3634: std_logic; attribute dont_touch of WX3634: signal is true;
	signal WX3635: std_logic; attribute dont_touch of WX3635: signal is true;
	signal WX3636: std_logic; attribute dont_touch of WX3636: signal is true;
	signal WX3637: std_logic; attribute dont_touch of WX3637: signal is true;
	signal WX3638: std_logic; attribute dont_touch of WX3638: signal is true;
	signal WX3639: std_logic; attribute dont_touch of WX3639: signal is true;
	signal WX3640: std_logic; attribute dont_touch of WX3640: signal is true;
	signal WX3641: std_logic; attribute dont_touch of WX3641: signal is true;
	signal WX3642: std_logic; attribute dont_touch of WX3642: signal is true;
	signal WX3643: std_logic; attribute dont_touch of WX3643: signal is true;
	signal WX3644: std_logic; attribute dont_touch of WX3644: signal is true;
	signal WX3645: std_logic; attribute dont_touch of WX3645: signal is true;
	signal WX3646: std_logic; attribute dont_touch of WX3646: signal is true;
	signal WX3647: std_logic; attribute dont_touch of WX3647: signal is true;
	signal WX3648: std_logic; attribute dont_touch of WX3648: signal is true;
	signal WX3649: std_logic; attribute dont_touch of WX3649: signal is true;
	signal WX3650: std_logic; attribute dont_touch of WX3650: signal is true;
	signal WX3651: std_logic; attribute dont_touch of WX3651: signal is true;
	signal WX3652: std_logic; attribute dont_touch of WX3652: signal is true;
	signal WX3653: std_logic; attribute dont_touch of WX3653: signal is true;
	signal WX3654: std_logic; attribute dont_touch of WX3654: signal is true;
	signal WX3655: std_logic; attribute dont_touch of WX3655: signal is true;
	signal WX3656: std_logic; attribute dont_touch of WX3656: signal is true;
	signal WX3657: std_logic; attribute dont_touch of WX3657: signal is true;
	signal WX3658: std_logic; attribute dont_touch of WX3658: signal is true;
	signal WX3659: std_logic; attribute dont_touch of WX3659: signal is true;
	signal WX3660: std_logic; attribute dont_touch of WX3660: signal is true;
	signal WX3661: std_logic; attribute dont_touch of WX3661: signal is true;
	signal WX3662: std_logic; attribute dont_touch of WX3662: signal is true;
	signal WX3663: std_logic; attribute dont_touch of WX3663: signal is true;
	signal WX3664: std_logic; attribute dont_touch of WX3664: signal is true;
	signal WX3665: std_logic; attribute dont_touch of WX3665: signal is true;
	signal WX3666: std_logic; attribute dont_touch of WX3666: signal is true;
	signal WX3667: std_logic; attribute dont_touch of WX3667: signal is true;
	signal WX3668: std_logic; attribute dont_touch of WX3668: signal is true;
	signal WX3669: std_logic; attribute dont_touch of WX3669: signal is true;
	signal WX3670: std_logic; attribute dont_touch of WX3670: signal is true;
	signal WX3671: std_logic; attribute dont_touch of WX3671: signal is true;
	signal WX3672: std_logic; attribute dont_touch of WX3672: signal is true;
	signal WX3673: std_logic; attribute dont_touch of WX3673: signal is true;
	signal WX3674: std_logic; attribute dont_touch of WX3674: signal is true;
	signal WX3675: std_logic; attribute dont_touch of WX3675: signal is true;
	signal WX3676: std_logic; attribute dont_touch of WX3676: signal is true;
	signal WX3677: std_logic; attribute dont_touch of WX3677: signal is true;
	signal WX3678: std_logic; attribute dont_touch of WX3678: signal is true;
	signal WX3679: std_logic; attribute dont_touch of WX3679: signal is true;
	signal WX3680: std_logic; attribute dont_touch of WX3680: signal is true;
	signal WX3681: std_logic; attribute dont_touch of WX3681: signal is true;
	signal WX3682: std_logic; attribute dont_touch of WX3682: signal is true;
	signal WX3683: std_logic; attribute dont_touch of WX3683: signal is true;
	signal WX3684: std_logic; attribute dont_touch of WX3684: signal is true;
	signal WX3685: std_logic; attribute dont_touch of WX3685: signal is true;
	signal WX3686: std_logic; attribute dont_touch of WX3686: signal is true;
	signal WX3687: std_logic; attribute dont_touch of WX3687: signal is true;
	signal WX3688: std_logic; attribute dont_touch of WX3688: signal is true;
	signal WX3689: std_logic; attribute dont_touch of WX3689: signal is true;
	signal WX3690: std_logic; attribute dont_touch of WX3690: signal is true;
	signal WX3691: std_logic; attribute dont_touch of WX3691: signal is true;
	signal WX3692: std_logic; attribute dont_touch of WX3692: signal is true;
	signal WX3693: std_logic; attribute dont_touch of WX3693: signal is true;
	signal WX3694: std_logic; attribute dont_touch of WX3694: signal is true;
	signal WX3695: std_logic; attribute dont_touch of WX3695: signal is true;
	signal WX3696: std_logic; attribute dont_touch of WX3696: signal is true;
	signal WX3697: std_logic; attribute dont_touch of WX3697: signal is true;
	signal WX3698: std_logic; attribute dont_touch of WX3698: signal is true;
	signal WX3699: std_logic; attribute dont_touch of WX3699: signal is true;
	signal WX3700: std_logic; attribute dont_touch of WX3700: signal is true;
	signal WX3701: std_logic; attribute dont_touch of WX3701: signal is true;
	signal WX3702: std_logic; attribute dont_touch of WX3702: signal is true;
	signal WX3703: std_logic; attribute dont_touch of WX3703: signal is true;
	signal WX3704: std_logic; attribute dont_touch of WX3704: signal is true;
	signal WX3705: std_logic; attribute dont_touch of WX3705: signal is true;
	signal WX3706: std_logic; attribute dont_touch of WX3706: signal is true;
	signal WX3707: std_logic; attribute dont_touch of WX3707: signal is true;
	signal WX3708: std_logic; attribute dont_touch of WX3708: signal is true;
	signal WX3709: std_logic; attribute dont_touch of WX3709: signal is true;
	signal WX3710: std_logic; attribute dont_touch of WX3710: signal is true;
	signal WX3711: std_logic; attribute dont_touch of WX3711: signal is true;
	signal WX3712: std_logic; attribute dont_touch of WX3712: signal is true;
	signal WX3713: std_logic; attribute dont_touch of WX3713: signal is true;
	signal WX3714: std_logic; attribute dont_touch of WX3714: signal is true;
	signal WX3715: std_logic; attribute dont_touch of WX3715: signal is true;
	signal WX3716: std_logic; attribute dont_touch of WX3716: signal is true;
	signal WX3717: std_logic; attribute dont_touch of WX3717: signal is true;
	signal WX3718: std_logic; attribute dont_touch of WX3718: signal is true;
	signal WX3719: std_logic; attribute dont_touch of WX3719: signal is true;
	signal WX3720: std_logic; attribute dont_touch of WX3720: signal is true;
	signal WX3721: std_logic; attribute dont_touch of WX3721: signal is true;
	signal WX3722: std_logic; attribute dont_touch of WX3722: signal is true;
	signal WX3723: std_logic; attribute dont_touch of WX3723: signal is true;
	signal WX3724: std_logic; attribute dont_touch of WX3724: signal is true;
	signal WX3725: std_logic; attribute dont_touch of WX3725: signal is true;
	signal WX3726: std_logic; attribute dont_touch of WX3726: signal is true;
	signal WX3727: std_logic; attribute dont_touch of WX3727: signal is true;
	signal WX3728: std_logic; attribute dont_touch of WX3728: signal is true;
	signal WX3729: std_logic; attribute dont_touch of WX3729: signal is true;
	signal WX3730: std_logic; attribute dont_touch of WX3730: signal is true;
	signal WX3731: std_logic; attribute dont_touch of WX3731: signal is true;
	signal WX3732: std_logic; attribute dont_touch of WX3732: signal is true;
	signal WX3733: std_logic; attribute dont_touch of WX3733: signal is true;
	signal WX3734: std_logic; attribute dont_touch of WX3734: signal is true;
	signal WX3735: std_logic; attribute dont_touch of WX3735: signal is true;
	signal WX3736: std_logic; attribute dont_touch of WX3736: signal is true;
	signal WX3737: std_logic; attribute dont_touch of WX3737: signal is true;
	signal WX3738: std_logic; attribute dont_touch of WX3738: signal is true;
	signal WX3739: std_logic; attribute dont_touch of WX3739: signal is true;
	signal WX3740: std_logic; attribute dont_touch of WX3740: signal is true;
	signal WX3741: std_logic; attribute dont_touch of WX3741: signal is true;
	signal WX3742: std_logic; attribute dont_touch of WX3742: signal is true;
	signal WX3743: std_logic; attribute dont_touch of WX3743: signal is true;
	signal WX3744: std_logic; attribute dont_touch of WX3744: signal is true;
	signal WX3745: std_logic; attribute dont_touch of WX3745: signal is true;
	signal WX3746: std_logic; attribute dont_touch of WX3746: signal is true;
	signal WX3747: std_logic; attribute dont_touch of WX3747: signal is true;
	signal WX3748: std_logic; attribute dont_touch of WX3748: signal is true;
	signal WX3749: std_logic; attribute dont_touch of WX3749: signal is true;
	signal WX3750: std_logic; attribute dont_touch of WX3750: signal is true;
	signal WX3751: std_logic; attribute dont_touch of WX3751: signal is true;
	signal WX3752: std_logic; attribute dont_touch of WX3752: signal is true;
	signal WX3753: std_logic; attribute dont_touch of WX3753: signal is true;
	signal WX3754: std_logic; attribute dont_touch of WX3754: signal is true;
	signal WX3755: std_logic; attribute dont_touch of WX3755: signal is true;
	signal WX3756: std_logic; attribute dont_touch of WX3756: signal is true;
	signal WX3757: std_logic; attribute dont_touch of WX3757: signal is true;
	signal WX3758: std_logic; attribute dont_touch of WX3758: signal is true;
	signal WX3759: std_logic; attribute dont_touch of WX3759: signal is true;
	signal WX3760: std_logic; attribute dont_touch of WX3760: signal is true;
	signal WX3761: std_logic; attribute dont_touch of WX3761: signal is true;
	signal WX3762: std_logic; attribute dont_touch of WX3762: signal is true;
	signal WX3763: std_logic; attribute dont_touch of WX3763: signal is true;
	signal WX3764: std_logic; attribute dont_touch of WX3764: signal is true;
	signal WX3765: std_logic; attribute dont_touch of WX3765: signal is true;
	signal WX3766: std_logic; attribute dont_touch of WX3766: signal is true;
	signal WX3767: std_logic; attribute dont_touch of WX3767: signal is true;
	signal WX3768: std_logic; attribute dont_touch of WX3768: signal is true;
	signal WX3769: std_logic; attribute dont_touch of WX3769: signal is true;
	signal WX3770: std_logic; attribute dont_touch of WX3770: signal is true;
	signal WX3771: std_logic; attribute dont_touch of WX3771: signal is true;
	signal WX3772: std_logic; attribute dont_touch of WX3772: signal is true;
	signal WX3773: std_logic; attribute dont_touch of WX3773: signal is true;
	signal WX3774: std_logic; attribute dont_touch of WX3774: signal is true;
	signal WX3775: std_logic; attribute dont_touch of WX3775: signal is true;
	signal WX3776: std_logic; attribute dont_touch of WX3776: signal is true;
	signal WX3777: std_logic; attribute dont_touch of WX3777: signal is true;
	signal WX3778: std_logic; attribute dont_touch of WX3778: signal is true;
	signal WX3779: std_logic; attribute dont_touch of WX3779: signal is true;
	signal WX3780: std_logic; attribute dont_touch of WX3780: signal is true;
	signal WX3781: std_logic; attribute dont_touch of WX3781: signal is true;
	signal WX3782: std_logic; attribute dont_touch of WX3782: signal is true;
	signal WX3783: std_logic; attribute dont_touch of WX3783: signal is true;
	signal WX3784: std_logic; attribute dont_touch of WX3784: signal is true;
	signal WX3785: std_logic; attribute dont_touch of WX3785: signal is true;
	signal WX3786: std_logic; attribute dont_touch of WX3786: signal is true;
	signal WX3787: std_logic; attribute dont_touch of WX3787: signal is true;
	signal WX3788: std_logic; attribute dont_touch of WX3788: signal is true;
	signal WX3789: std_logic; attribute dont_touch of WX3789: signal is true;
	signal WX3790: std_logic; attribute dont_touch of WX3790: signal is true;
	signal WX3791: std_logic; attribute dont_touch of WX3791: signal is true;
	signal WX3792: std_logic; attribute dont_touch of WX3792: signal is true;
	signal WX3793: std_logic; attribute dont_touch of WX3793: signal is true;
	signal WX3794: std_logic; attribute dont_touch of WX3794: signal is true;
	signal WX3795: std_logic; attribute dont_touch of WX3795: signal is true;
	signal WX3796: std_logic; attribute dont_touch of WX3796: signal is true;
	signal WX3797: std_logic; attribute dont_touch of WX3797: signal is true;
	signal WX3798: std_logic; attribute dont_touch of WX3798: signal is true;
	signal WX3799: std_logic; attribute dont_touch of WX3799: signal is true;
	signal WX3800: std_logic; attribute dont_touch of WX3800: signal is true;
	signal WX3801: std_logic; attribute dont_touch of WX3801: signal is true;
	signal WX3802: std_logic; attribute dont_touch of WX3802: signal is true;
	signal WX3803: std_logic; attribute dont_touch of WX3803: signal is true;
	signal WX3804: std_logic; attribute dont_touch of WX3804: signal is true;
	signal WX3805: std_logic; attribute dont_touch of WX3805: signal is true;
	signal WX3806: std_logic; attribute dont_touch of WX3806: signal is true;
	signal WX3807: std_logic; attribute dont_touch of WX3807: signal is true;
	signal WX3808: std_logic; attribute dont_touch of WX3808: signal is true;
	signal WX3809: std_logic; attribute dont_touch of WX3809: signal is true;
	signal WX3810: std_logic; attribute dont_touch of WX3810: signal is true;
	signal WX3811: std_logic; attribute dont_touch of WX3811: signal is true;
	signal WX3812: std_logic; attribute dont_touch of WX3812: signal is true;
	signal WX3813: std_logic; attribute dont_touch of WX3813: signal is true;
	signal WX3814: std_logic; attribute dont_touch of WX3814: signal is true;
	signal WX3815: std_logic; attribute dont_touch of WX3815: signal is true;
	signal WX3816: std_logic; attribute dont_touch of WX3816: signal is true;
	signal WX3817: std_logic; attribute dont_touch of WX3817: signal is true;
	signal WX3818: std_logic; attribute dont_touch of WX3818: signal is true;
	signal WX3819: std_logic; attribute dont_touch of WX3819: signal is true;
	signal WX3820: std_logic; attribute dont_touch of WX3820: signal is true;
	signal WX3821: std_logic; attribute dont_touch of WX3821: signal is true;
	signal WX3822: std_logic; attribute dont_touch of WX3822: signal is true;
	signal WX3823: std_logic; attribute dont_touch of WX3823: signal is true;
	signal WX3824: std_logic; attribute dont_touch of WX3824: signal is true;
	signal WX3825: std_logic; attribute dont_touch of WX3825: signal is true;
	signal WX3826: std_logic; attribute dont_touch of WX3826: signal is true;
	signal WX3827: std_logic; attribute dont_touch of WX3827: signal is true;
	signal WX3828: std_logic; attribute dont_touch of WX3828: signal is true;
	signal WX3829: std_logic; attribute dont_touch of WX3829: signal is true;
	signal WX3830: std_logic; attribute dont_touch of WX3830: signal is true;
	signal WX3831: std_logic; attribute dont_touch of WX3831: signal is true;
	signal WX3832: std_logic; attribute dont_touch of WX3832: signal is true;
	signal WX3833: std_logic; attribute dont_touch of WX3833: signal is true;
	signal WX3834: std_logic; attribute dont_touch of WX3834: signal is true;
	signal WX3835: std_logic; attribute dont_touch of WX3835: signal is true;
	signal WX3836: std_logic; attribute dont_touch of WX3836: signal is true;
	signal WX3837: std_logic; attribute dont_touch of WX3837: signal is true;
	signal WX3838: std_logic; attribute dont_touch of WX3838: signal is true;
	signal WX3839: std_logic; attribute dont_touch of WX3839: signal is true;
	signal WX3840: std_logic; attribute dont_touch of WX3840: signal is true;
	signal WX3841: std_logic; attribute dont_touch of WX3841: signal is true;
	signal WX3842: std_logic; attribute dont_touch of WX3842: signal is true;
	signal WX3843: std_logic; attribute dont_touch of WX3843: signal is true;
	signal WX3844: std_logic; attribute dont_touch of WX3844: signal is true;
	signal WX3845: std_logic; attribute dont_touch of WX3845: signal is true;
	signal WX3846: std_logic; attribute dont_touch of WX3846: signal is true;
	signal WX3847: std_logic; attribute dont_touch of WX3847: signal is true;
	signal WX3848: std_logic; attribute dont_touch of WX3848: signal is true;
	signal WX3849: std_logic; attribute dont_touch of WX3849: signal is true;
	signal WX3850: std_logic; attribute dont_touch of WX3850: signal is true;
	signal WX3852: std_logic; attribute dont_touch of WX3852: signal is true;
	signal WX3854: std_logic; attribute dont_touch of WX3854: signal is true;
	signal WX3856: std_logic; attribute dont_touch of WX3856: signal is true;
	signal WX3858: std_logic; attribute dont_touch of WX3858: signal is true;
	signal WX3860: std_logic; attribute dont_touch of WX3860: signal is true;
	signal WX3862: std_logic; attribute dont_touch of WX3862: signal is true;
	signal WX3864: std_logic; attribute dont_touch of WX3864: signal is true;
	signal WX3866: std_logic; attribute dont_touch of WX3866: signal is true;
	signal WX3868: std_logic; attribute dont_touch of WX3868: signal is true;
	signal WX3870: std_logic; attribute dont_touch of WX3870: signal is true;
	signal WX3872: std_logic; attribute dont_touch of WX3872: signal is true;
	signal WX3874: std_logic; attribute dont_touch of WX3874: signal is true;
	signal WX3876: std_logic; attribute dont_touch of WX3876: signal is true;
	signal WX3878: std_logic; attribute dont_touch of WX3878: signal is true;
	signal WX3880: std_logic; attribute dont_touch of WX3880: signal is true;
	signal WX3882: std_logic; attribute dont_touch of WX3882: signal is true;
	signal WX3884: std_logic; attribute dont_touch of WX3884: signal is true;
	signal WX3886: std_logic; attribute dont_touch of WX3886: signal is true;
	signal WX3888: std_logic; attribute dont_touch of WX3888: signal is true;
	signal WX3890: std_logic; attribute dont_touch of WX3890: signal is true;
	signal WX3892: std_logic; attribute dont_touch of WX3892: signal is true;
	signal WX3894: std_logic; attribute dont_touch of WX3894: signal is true;
	signal WX3896: std_logic; attribute dont_touch of WX3896: signal is true;
	signal WX3898: std_logic; attribute dont_touch of WX3898: signal is true;
	signal WX3900: std_logic; attribute dont_touch of WX3900: signal is true;
	signal WX3902: std_logic; attribute dont_touch of WX3902: signal is true;
	signal WX3904: std_logic; attribute dont_touch of WX3904: signal is true;
	signal WX3906: std_logic; attribute dont_touch of WX3906: signal is true;
	signal WX3908: std_logic; attribute dont_touch of WX3908: signal is true;
	signal WX3910: std_logic; attribute dont_touch of WX3910: signal is true;
	signal WX3912: std_logic; attribute dont_touch of WX3912: signal is true;
	signal WX3914: std_logic; attribute dont_touch of WX3914: signal is true;
	signal WX3915: std_logic; attribute dont_touch of WX3915: signal is true;
	signal WX3916: std_logic; attribute dont_touch of WX3916: signal is true;
	signal WX3917: std_logic; attribute dont_touch of WX3917: signal is true;
	signal WX3918: std_logic; attribute dont_touch of WX3918: signal is true;
	signal WX3919: std_logic; attribute dont_touch of WX3919: signal is true;
	signal WX3920: std_logic; attribute dont_touch of WX3920: signal is true;
	signal WX3921: std_logic; attribute dont_touch of WX3921: signal is true;
	signal WX3922: std_logic; attribute dont_touch of WX3922: signal is true;
	signal WX3923: std_logic; attribute dont_touch of WX3923: signal is true;
	signal WX3924: std_logic; attribute dont_touch of WX3924: signal is true;
	signal WX3925: std_logic; attribute dont_touch of WX3925: signal is true;
	signal WX3926: std_logic; attribute dont_touch of WX3926: signal is true;
	signal WX3927: std_logic; attribute dont_touch of WX3927: signal is true;
	signal WX3928: std_logic; attribute dont_touch of WX3928: signal is true;
	signal WX3929: std_logic; attribute dont_touch of WX3929: signal is true;
	signal WX3930: std_logic; attribute dont_touch of WX3930: signal is true;
	signal WX3931: std_logic; attribute dont_touch of WX3931: signal is true;
	signal WX3932: std_logic; attribute dont_touch of WX3932: signal is true;
	signal WX3933: std_logic; attribute dont_touch of WX3933: signal is true;
	signal WX3934: std_logic; attribute dont_touch of WX3934: signal is true;
	signal WX3935: std_logic; attribute dont_touch of WX3935: signal is true;
	signal WX3936: std_logic; attribute dont_touch of WX3936: signal is true;
	signal WX3937: std_logic; attribute dont_touch of WX3937: signal is true;
	signal WX3938: std_logic; attribute dont_touch of WX3938: signal is true;
	signal WX3939: std_logic; attribute dont_touch of WX3939: signal is true;
	signal WX3940: std_logic; attribute dont_touch of WX3940: signal is true;
	signal WX3941: std_logic; attribute dont_touch of WX3941: signal is true;
	signal WX3942: std_logic; attribute dont_touch of WX3942: signal is true;
	signal WX3943: std_logic; attribute dont_touch of WX3943: signal is true;
	signal WX3944: std_logic; attribute dont_touch of WX3944: signal is true;
	signal WX3945: std_logic; attribute dont_touch of WX3945: signal is true;
	signal WX3946: std_logic; attribute dont_touch of WX3946: signal is true;
	signal WX3947: std_logic; attribute dont_touch of WX3947: signal is true;
	signal WX3948: std_logic; attribute dont_touch of WX3948: signal is true;
	signal WX3949: std_logic; attribute dont_touch of WX3949: signal is true;
	signal WX3950: std_logic; attribute dont_touch of WX3950: signal is true;
	signal WX3951: std_logic; attribute dont_touch of WX3951: signal is true;
	signal WX3952: std_logic; attribute dont_touch of WX3952: signal is true;
	signal WX3953: std_logic; attribute dont_touch of WX3953: signal is true;
	signal WX3954: std_logic; attribute dont_touch of WX3954: signal is true;
	signal WX3955: std_logic; attribute dont_touch of WX3955: signal is true;
	signal WX3956: std_logic; attribute dont_touch of WX3956: signal is true;
	signal WX3957: std_logic; attribute dont_touch of WX3957: signal is true;
	signal WX3958: std_logic; attribute dont_touch of WX3958: signal is true;
	signal WX3959: std_logic; attribute dont_touch of WX3959: signal is true;
	signal WX3960: std_logic; attribute dont_touch of WX3960: signal is true;
	signal WX3961: std_logic; attribute dont_touch of WX3961: signal is true;
	signal WX3962: std_logic; attribute dont_touch of WX3962: signal is true;
	signal WX3963: std_logic; attribute dont_touch of WX3963: signal is true;
	signal WX3964: std_logic; attribute dont_touch of WX3964: signal is true;
	signal WX3965: std_logic; attribute dont_touch of WX3965: signal is true;
	signal WX3966: std_logic; attribute dont_touch of WX3966: signal is true;
	signal WX3967: std_logic; attribute dont_touch of WX3967: signal is true;
	signal WX3968: std_logic; attribute dont_touch of WX3968: signal is true;
	signal WX3969: std_logic; attribute dont_touch of WX3969: signal is true;
	signal WX3970: std_logic; attribute dont_touch of WX3970: signal is true;
	signal WX3971: std_logic; attribute dont_touch of WX3971: signal is true;
	signal WX3972: std_logic; attribute dont_touch of WX3972: signal is true;
	signal WX3973: std_logic; attribute dont_touch of WX3973: signal is true;
	signal WX3974: std_logic; attribute dont_touch of WX3974: signal is true;
	signal WX3975: std_logic; attribute dont_touch of WX3975: signal is true;
	signal WX3976: std_logic; attribute dont_touch of WX3976: signal is true;
	signal WX3977: std_logic; attribute dont_touch of WX3977: signal is true;
	signal WX3978: std_logic; attribute dont_touch of WX3978: signal is true;
	signal WX3979: std_logic; attribute dont_touch of WX3979: signal is true;
	signal WX3980: std_logic; attribute dont_touch of WX3980: signal is true;
	signal WX3981: std_logic; attribute dont_touch of WX3981: signal is true;
	signal WX3982: std_logic; attribute dont_touch of WX3982: signal is true;
	signal WX3983: std_logic; attribute dont_touch of WX3983: signal is true;
	signal WX3984: std_logic; attribute dont_touch of WX3984: signal is true;
	signal WX3985: std_logic; attribute dont_touch of WX3985: signal is true;
	signal WX3986: std_logic; attribute dont_touch of WX3986: signal is true;
	signal WX3987: std_logic; attribute dont_touch of WX3987: signal is true;
	signal WX3988: std_logic; attribute dont_touch of WX3988: signal is true;
	signal WX3989: std_logic; attribute dont_touch of WX3989: signal is true;
	signal WX3990: std_logic; attribute dont_touch of WX3990: signal is true;
	signal WX3991: std_logic; attribute dont_touch of WX3991: signal is true;
	signal WX3992: std_logic; attribute dont_touch of WX3992: signal is true;
	signal WX3993: std_logic; attribute dont_touch of WX3993: signal is true;
	signal WX3994: std_logic; attribute dont_touch of WX3994: signal is true;
	signal WX3995: std_logic; attribute dont_touch of WX3995: signal is true;
	signal WX3996: std_logic; attribute dont_touch of WX3996: signal is true;
	signal WX3997: std_logic; attribute dont_touch of WX3997: signal is true;
	signal WX3998: std_logic; attribute dont_touch of WX3998: signal is true;
	signal WX3999: std_logic; attribute dont_touch of WX3999: signal is true;
	signal WX4000: std_logic; attribute dont_touch of WX4000: signal is true;
	signal WX4001: std_logic; attribute dont_touch of WX4001: signal is true;
	signal WX4002: std_logic; attribute dont_touch of WX4002: signal is true;
	signal WX4003: std_logic; attribute dont_touch of WX4003: signal is true;
	signal WX4004: std_logic; attribute dont_touch of WX4004: signal is true;
	signal WX4005: std_logic; attribute dont_touch of WX4005: signal is true;
	signal WX4006: std_logic; attribute dont_touch of WX4006: signal is true;
	signal WX4007: std_logic; attribute dont_touch of WX4007: signal is true;
	signal WX4008: std_logic; attribute dont_touch of WX4008: signal is true;
	signal WX4009: std_logic; attribute dont_touch of WX4009: signal is true;
	signal WX4010: std_logic; attribute dont_touch of WX4010: signal is true;
	signal WX4011: std_logic; attribute dont_touch of WX4011: signal is true;
	signal WX4012: std_logic; attribute dont_touch of WX4012: signal is true;
	signal WX4013: std_logic; attribute dont_touch of WX4013: signal is true;
	signal WX4014: std_logic; attribute dont_touch of WX4014: signal is true;
	signal WX4015: std_logic; attribute dont_touch of WX4015: signal is true;
	signal WX4016: std_logic; attribute dont_touch of WX4016: signal is true;
	signal WX4017: std_logic; attribute dont_touch of WX4017: signal is true;
	signal WX4018: std_logic; attribute dont_touch of WX4018: signal is true;
	signal WX4019: std_logic; attribute dont_touch of WX4019: signal is true;
	signal WX4020: std_logic; attribute dont_touch of WX4020: signal is true;
	signal WX4021: std_logic; attribute dont_touch of WX4021: signal is true;
	signal WX4022: std_logic; attribute dont_touch of WX4022: signal is true;
	signal WX4023: std_logic; attribute dont_touch of WX4023: signal is true;
	signal WX4024: std_logic; attribute dont_touch of WX4024: signal is true;
	signal WX4025: std_logic; attribute dont_touch of WX4025: signal is true;
	signal WX4026: std_logic; attribute dont_touch of WX4026: signal is true;
	signal WX4027: std_logic; attribute dont_touch of WX4027: signal is true;
	signal WX4028: std_logic; attribute dont_touch of WX4028: signal is true;
	signal WX4029: std_logic; attribute dont_touch of WX4029: signal is true;
	signal WX4030: std_logic; attribute dont_touch of WX4030: signal is true;
	signal WX4031: std_logic; attribute dont_touch of WX4031: signal is true;
	signal WX4032: std_logic; attribute dont_touch of WX4032: signal is true;
	signal WX4033: std_logic; attribute dont_touch of WX4033: signal is true;
	signal WX4034: std_logic; attribute dont_touch of WX4034: signal is true;
	signal WX4035: std_logic; attribute dont_touch of WX4035: signal is true;
	signal WX4036: std_logic; attribute dont_touch of WX4036: signal is true;
	signal WX4037: std_logic; attribute dont_touch of WX4037: signal is true;
	signal WX4038: std_logic; attribute dont_touch of WX4038: signal is true;
	signal WX4039: std_logic; attribute dont_touch of WX4039: signal is true;
	signal WX4040: std_logic; attribute dont_touch of WX4040: signal is true;
	signal WX4041: std_logic; attribute dont_touch of WX4041: signal is true;
	signal WX4042: std_logic; attribute dont_touch of WX4042: signal is true;
	signal WX4043: std_logic; attribute dont_touch of WX4043: signal is true;
	signal WX4044: std_logic; attribute dont_touch of WX4044: signal is true;
	signal WX4045: std_logic; attribute dont_touch of WX4045: signal is true;
	signal WX4046: std_logic; attribute dont_touch of WX4046: signal is true;
	signal WX4047: std_logic; attribute dont_touch of WX4047: signal is true;
	signal WX4048: std_logic; attribute dont_touch of WX4048: signal is true;
	signal WX4049: std_logic; attribute dont_touch of WX4049: signal is true;
	signal WX4050: std_logic; attribute dont_touch of WX4050: signal is true;
	signal WX4051: std_logic; attribute dont_touch of WX4051: signal is true;
	signal WX4052: std_logic; attribute dont_touch of WX4052: signal is true;
	signal WX4053: std_logic; attribute dont_touch of WX4053: signal is true;
	signal WX4054: std_logic; attribute dont_touch of WX4054: signal is true;
	signal WX4055: std_logic; attribute dont_touch of WX4055: signal is true;
	signal WX4056: std_logic; attribute dont_touch of WX4056: signal is true;
	signal WX4057: std_logic; attribute dont_touch of WX4057: signal is true;
	signal WX4058: std_logic; attribute dont_touch of WX4058: signal is true;
	signal WX4059: std_logic; attribute dont_touch of WX4059: signal is true;
	signal WX4060: std_logic; attribute dont_touch of WX4060: signal is true;
	signal WX4061: std_logic; attribute dont_touch of WX4061: signal is true;
	signal WX4062: std_logic; attribute dont_touch of WX4062: signal is true;
	signal WX4063: std_logic; attribute dont_touch of WX4063: signal is true;
	signal WX4064: std_logic; attribute dont_touch of WX4064: signal is true;
	signal WX4065: std_logic; attribute dont_touch of WX4065: signal is true;
	signal WX4066: std_logic; attribute dont_touch of WX4066: signal is true;
	signal WX4067: std_logic; attribute dont_touch of WX4067: signal is true;
	signal WX4068: std_logic; attribute dont_touch of WX4068: signal is true;
	signal WX4069: std_logic; attribute dont_touch of WX4069: signal is true;
	signal WX4070: std_logic; attribute dont_touch of WX4070: signal is true;
	signal WX4071: std_logic; attribute dont_touch of WX4071: signal is true;
	signal WX4072: std_logic; attribute dont_touch of WX4072: signal is true;
	signal WX4073: std_logic; attribute dont_touch of WX4073: signal is true;
	signal WX4074: std_logic; attribute dont_touch of WX4074: signal is true;
	signal WX4075: std_logic; attribute dont_touch of WX4075: signal is true;
	signal WX4076: std_logic; attribute dont_touch of WX4076: signal is true;
	signal WX4077: std_logic; attribute dont_touch of WX4077: signal is true;
	signal WX4078: std_logic; attribute dont_touch of WX4078: signal is true;
	signal WX4079: std_logic; attribute dont_touch of WX4079: signal is true;
	signal WX4080: std_logic; attribute dont_touch of WX4080: signal is true;
	signal WX4081: std_logic; attribute dont_touch of WX4081: signal is true;
	signal WX4082: std_logic; attribute dont_touch of WX4082: signal is true;
	signal WX4083: std_logic; attribute dont_touch of WX4083: signal is true;
	signal WX4084: std_logic; attribute dont_touch of WX4084: signal is true;
	signal WX4085: std_logic; attribute dont_touch of WX4085: signal is true;
	signal WX4086: std_logic; attribute dont_touch of WX4086: signal is true;
	signal WX4087: std_logic; attribute dont_touch of WX4087: signal is true;
	signal WX4088: std_logic; attribute dont_touch of WX4088: signal is true;
	signal WX4089: std_logic; attribute dont_touch of WX4089: signal is true;
	signal WX4090: std_logic; attribute dont_touch of WX4090: signal is true;
	signal WX4091: std_logic; attribute dont_touch of WX4091: signal is true;
	signal WX4092: std_logic; attribute dont_touch of WX4092: signal is true;
	signal WX4093: std_logic; attribute dont_touch of WX4093: signal is true;
	signal WX4094: std_logic; attribute dont_touch of WX4094: signal is true;
	signal WX4095: std_logic; attribute dont_touch of WX4095: signal is true;
	signal WX4096: std_logic; attribute dont_touch of WX4096: signal is true;
	signal WX4097: std_logic; attribute dont_touch of WX4097: signal is true;
	signal WX4098: std_logic; attribute dont_touch of WX4098: signal is true;
	signal WX4099: std_logic; attribute dont_touch of WX4099: signal is true;
	signal WX4100: std_logic; attribute dont_touch of WX4100: signal is true;
	signal WX4101: std_logic; attribute dont_touch of WX4101: signal is true;
	signal WX4102: std_logic; attribute dont_touch of WX4102: signal is true;
	signal WX4103: std_logic; attribute dont_touch of WX4103: signal is true;
	signal WX4104: std_logic; attribute dont_touch of WX4104: signal is true;
	signal WX4105: std_logic; attribute dont_touch of WX4105: signal is true;
	signal WX4106: std_logic; attribute dont_touch of WX4106: signal is true;
	signal WX4107: std_logic; attribute dont_touch of WX4107: signal is true;
	signal WX4108: std_logic; attribute dont_touch of WX4108: signal is true;
	signal WX4109: std_logic; attribute dont_touch of WX4109: signal is true;
	signal WX4110: std_logic; attribute dont_touch of WX4110: signal is true;
	signal WX4111: std_logic; attribute dont_touch of WX4111: signal is true;
	signal WX4112: std_logic; attribute dont_touch of WX4112: signal is true;
	signal WX4113: std_logic; attribute dont_touch of WX4113: signal is true;
	signal WX4114: std_logic; attribute dont_touch of WX4114: signal is true;
	signal WX4115: std_logic; attribute dont_touch of WX4115: signal is true;
	signal WX4116: std_logic; attribute dont_touch of WX4116: signal is true;
	signal WX4117: std_logic; attribute dont_touch of WX4117: signal is true;
	signal WX4118: std_logic; attribute dont_touch of WX4118: signal is true;
	signal WX4119: std_logic; attribute dont_touch of WX4119: signal is true;
	signal WX4120: std_logic; attribute dont_touch of WX4120: signal is true;
	signal WX4121: std_logic; attribute dont_touch of WX4121: signal is true;
	signal WX4122: std_logic; attribute dont_touch of WX4122: signal is true;
	signal WX4123: std_logic; attribute dont_touch of WX4123: signal is true;
	signal WX4124: std_logic; attribute dont_touch of WX4124: signal is true;
	signal WX4125: std_logic; attribute dont_touch of WX4125: signal is true;
	signal WX4126: std_logic; attribute dont_touch of WX4126: signal is true;
	signal WX4127: std_logic; attribute dont_touch of WX4127: signal is true;
	signal WX4128: std_logic; attribute dont_touch of WX4128: signal is true;
	signal WX4129: std_logic; attribute dont_touch of WX4129: signal is true;
	signal WX4130: std_logic; attribute dont_touch of WX4130: signal is true;
	signal WX4131: std_logic; attribute dont_touch of WX4131: signal is true;
	signal WX4132: std_logic; attribute dont_touch of WX4132: signal is true;
	signal WX4133: std_logic; attribute dont_touch of WX4133: signal is true;
	signal WX4134: std_logic; attribute dont_touch of WX4134: signal is true;
	signal WX4135: std_logic; attribute dont_touch of WX4135: signal is true;
	signal WX4136: std_logic; attribute dont_touch of WX4136: signal is true;
	signal WX4137: std_logic; attribute dont_touch of WX4137: signal is true;
	signal WX4138: std_logic; attribute dont_touch of WX4138: signal is true;
	signal WX4139: std_logic; attribute dont_touch of WX4139: signal is true;
	signal WX4140: std_logic; attribute dont_touch of WX4140: signal is true;
	signal WX4141: std_logic; attribute dont_touch of WX4141: signal is true;
	signal WX4142: std_logic; attribute dont_touch of WX4142: signal is true;
	signal WX4143: std_logic; attribute dont_touch of WX4143: signal is true;
	signal WX4144: std_logic; attribute dont_touch of WX4144: signal is true;
	signal WX4145: std_logic; attribute dont_touch of WX4145: signal is true;
	signal WX4146: std_logic; attribute dont_touch of WX4146: signal is true;
	signal WX4147: std_logic; attribute dont_touch of WX4147: signal is true;
	signal WX4148: std_logic; attribute dont_touch of WX4148: signal is true;
	signal WX4149: std_logic; attribute dont_touch of WX4149: signal is true;
	signal WX4150: std_logic; attribute dont_touch of WX4150: signal is true;
	signal WX4151: std_logic; attribute dont_touch of WX4151: signal is true;
	signal WX4152: std_logic; attribute dont_touch of WX4152: signal is true;
	signal WX4153: std_logic; attribute dont_touch of WX4153: signal is true;
	signal WX4154: std_logic; attribute dont_touch of WX4154: signal is true;
	signal WX4155: std_logic; attribute dont_touch of WX4155: signal is true;
	signal WX4156: std_logic; attribute dont_touch of WX4156: signal is true;
	signal WX4157: std_logic; attribute dont_touch of WX4157: signal is true;
	signal WX4158: std_logic; attribute dont_touch of WX4158: signal is true;
	signal WX4159: std_logic; attribute dont_touch of WX4159: signal is true;
	signal WX4160: std_logic; attribute dont_touch of WX4160: signal is true;
	signal WX4161: std_logic; attribute dont_touch of WX4161: signal is true;
	signal WX4162: std_logic; attribute dont_touch of WX4162: signal is true;
	signal WX4163: std_logic; attribute dont_touch of WX4163: signal is true;
	signal WX4164: std_logic; attribute dont_touch of WX4164: signal is true;
	signal WX4165: std_logic; attribute dont_touch of WX4165: signal is true;
	signal WX4166: std_logic; attribute dont_touch of WX4166: signal is true;
	signal WX4167: std_logic; attribute dont_touch of WX4167: signal is true;
	signal WX4168: std_logic; attribute dont_touch of WX4168: signal is true;
	signal WX4169: std_logic; attribute dont_touch of WX4169: signal is true;
	signal WX4170: std_logic; attribute dont_touch of WX4170: signal is true;
	signal WX4171: std_logic; attribute dont_touch of WX4171: signal is true;
	signal WX4172: std_logic; attribute dont_touch of WX4172: signal is true;
	signal WX4173: std_logic; attribute dont_touch of WX4173: signal is true;
	signal WX4174: std_logic; attribute dont_touch of WX4174: signal is true;
	signal WX4175: std_logic; attribute dont_touch of WX4175: signal is true;
	signal WX4176: std_logic; attribute dont_touch of WX4176: signal is true;
	signal WX4177: std_logic; attribute dont_touch of WX4177: signal is true;
	signal WX4178: std_logic; attribute dont_touch of WX4178: signal is true;
	signal WX4179: std_logic; attribute dont_touch of WX4179: signal is true;
	signal WX4180: std_logic; attribute dont_touch of WX4180: signal is true;
	signal WX4181: std_logic; attribute dont_touch of WX4181: signal is true;
	signal WX4182: std_logic; attribute dont_touch of WX4182: signal is true;
	signal WX4183: std_logic; attribute dont_touch of WX4183: signal is true;
	signal WX4184: std_logic; attribute dont_touch of WX4184: signal is true;
	signal WX4185: std_logic; attribute dont_touch of WX4185: signal is true;
	signal WX4186: std_logic; attribute dont_touch of WX4186: signal is true;
	signal WX4187: std_logic; attribute dont_touch of WX4187: signal is true;
	signal WX4188: std_logic; attribute dont_touch of WX4188: signal is true;
	signal WX4189: std_logic; attribute dont_touch of WX4189: signal is true;
	signal WX4190: std_logic; attribute dont_touch of WX4190: signal is true;
	signal WX4191: std_logic; attribute dont_touch of WX4191: signal is true;
	signal WX4192: std_logic; attribute dont_touch of WX4192: signal is true;
	signal WX4193: std_logic; attribute dont_touch of WX4193: signal is true;
	signal WX4194: std_logic; attribute dont_touch of WX4194: signal is true;
	signal WX4195: std_logic; attribute dont_touch of WX4195: signal is true;
	signal WX4196: std_logic; attribute dont_touch of WX4196: signal is true;
	signal WX4197: std_logic; attribute dont_touch of WX4197: signal is true;
	signal WX4198: std_logic; attribute dont_touch of WX4198: signal is true;
	signal WX4199: std_logic; attribute dont_touch of WX4199: signal is true;
	signal WX4200: std_logic; attribute dont_touch of WX4200: signal is true;
	signal WX4201: std_logic; attribute dont_touch of WX4201: signal is true;
	signal WX4202: std_logic; attribute dont_touch of WX4202: signal is true;
	signal WX4203: std_logic; attribute dont_touch of WX4203: signal is true;
	signal WX4204: std_logic; attribute dont_touch of WX4204: signal is true;
	signal WX4205: std_logic; attribute dont_touch of WX4205: signal is true;
	signal WX4206: std_logic; attribute dont_touch of WX4206: signal is true;
	signal WX4207: std_logic; attribute dont_touch of WX4207: signal is true;
	signal WX4208: std_logic; attribute dont_touch of WX4208: signal is true;
	signal WX4209: std_logic; attribute dont_touch of WX4209: signal is true;
	signal WX4210: std_logic; attribute dont_touch of WX4210: signal is true;
	signal WX4211: std_logic; attribute dont_touch of WX4211: signal is true;
	signal WX4212: std_logic; attribute dont_touch of WX4212: signal is true;
	signal WX4213: std_logic; attribute dont_touch of WX4213: signal is true;
	signal WX4214: std_logic; attribute dont_touch of WX4214: signal is true;
	signal WX4215: std_logic; attribute dont_touch of WX4215: signal is true;
	signal WX4216: std_logic; attribute dont_touch of WX4216: signal is true;
	signal WX4217: std_logic; attribute dont_touch of WX4217: signal is true;
	signal WX4218: std_logic; attribute dont_touch of WX4218: signal is true;
	signal WX4219: std_logic; attribute dont_touch of WX4219: signal is true;
	signal WX4220: std_logic; attribute dont_touch of WX4220: signal is true;
	signal WX4221: std_logic; attribute dont_touch of WX4221: signal is true;
	signal WX4222: std_logic; attribute dont_touch of WX4222: signal is true;
	signal WX4223: std_logic; attribute dont_touch of WX4223: signal is true;
	signal WX4224: std_logic; attribute dont_touch of WX4224: signal is true;
	signal WX4225: std_logic; attribute dont_touch of WX4225: signal is true;
	signal WX4226: std_logic; attribute dont_touch of WX4226: signal is true;
	signal WX4227: std_logic; attribute dont_touch of WX4227: signal is true;
	signal WX4228: std_logic; attribute dont_touch of WX4228: signal is true;
	signal WX4229: std_logic; attribute dont_touch of WX4229: signal is true;
	signal WX4230: std_logic; attribute dont_touch of WX4230: signal is true;
	signal WX4231: std_logic; attribute dont_touch of WX4231: signal is true;
	signal WX4232: std_logic; attribute dont_touch of WX4232: signal is true;
	signal WX4233: std_logic; attribute dont_touch of WX4233: signal is true;
	signal WX4234: std_logic; attribute dont_touch of WX4234: signal is true;
	signal WX4235: std_logic; attribute dont_touch of WX4235: signal is true;
	signal WX4236: std_logic; attribute dont_touch of WX4236: signal is true;
	signal WX4237: std_logic; attribute dont_touch of WX4237: signal is true;
	signal WX4238: std_logic; attribute dont_touch of WX4238: signal is true;
	signal WX4239: std_logic; attribute dont_touch of WX4239: signal is true;
	signal WX4240: std_logic; attribute dont_touch of WX4240: signal is true;
	signal WX4241: std_logic; attribute dont_touch of WX4241: signal is true;
	signal WX4242: std_logic; attribute dont_touch of WX4242: signal is true;
	signal WX4243: std_logic; attribute dont_touch of WX4243: signal is true;
	signal WX4244: std_logic; attribute dont_touch of WX4244: signal is true;
	signal WX4245: std_logic; attribute dont_touch of WX4245: signal is true;
	signal WX4246: std_logic; attribute dont_touch of WX4246: signal is true;
	signal WX4247: std_logic; attribute dont_touch of WX4247: signal is true;
	signal WX4248: std_logic; attribute dont_touch of WX4248: signal is true;
	signal WX4249: std_logic; attribute dont_touch of WX4249: signal is true;
	signal WX4250: std_logic; attribute dont_touch of WX4250: signal is true;
	signal WX4251: std_logic; attribute dont_touch of WX4251: signal is true;
	signal WX4252: std_logic; attribute dont_touch of WX4252: signal is true;
	signal WX4253: std_logic; attribute dont_touch of WX4253: signal is true;
	signal WX4254: std_logic; attribute dont_touch of WX4254: signal is true;
	signal WX4255: std_logic; attribute dont_touch of WX4255: signal is true;
	signal WX4256: std_logic; attribute dont_touch of WX4256: signal is true;
	signal WX4257: std_logic; attribute dont_touch of WX4257: signal is true;
	signal WX4258: std_logic; attribute dont_touch of WX4258: signal is true;
	signal WX4259: std_logic; attribute dont_touch of WX4259: signal is true;
	signal WX4260: std_logic; attribute dont_touch of WX4260: signal is true;
	signal WX4261: std_logic; attribute dont_touch of WX4261: signal is true;
	signal WX4262: std_logic; attribute dont_touch of WX4262: signal is true;
	signal WX4263: std_logic; attribute dont_touch of WX4263: signal is true;
	signal WX4264: std_logic; attribute dont_touch of WX4264: signal is true;
	signal WX4265: std_logic; attribute dont_touch of WX4265: signal is true;
	signal WX4266: std_logic; attribute dont_touch of WX4266: signal is true;
	signal WX4267: std_logic; attribute dont_touch of WX4267: signal is true;
	signal WX4268: std_logic; attribute dont_touch of WX4268: signal is true;
	signal WX4269: std_logic; attribute dont_touch of WX4269: signal is true;
	signal WX4270: std_logic; attribute dont_touch of WX4270: signal is true;
	signal WX4271: std_logic; attribute dont_touch of WX4271: signal is true;
	signal WX4272: std_logic; attribute dont_touch of WX4272: signal is true;
	signal WX4273: std_logic; attribute dont_touch of WX4273: signal is true;
	signal WX4274: std_logic; attribute dont_touch of WX4274: signal is true;
	signal WX4275: std_logic; attribute dont_touch of WX4275: signal is true;
	signal WX4276: std_logic; attribute dont_touch of WX4276: signal is true;
	signal WX4277: std_logic; attribute dont_touch of WX4277: signal is true;
	signal WX4278: std_logic; attribute dont_touch of WX4278: signal is true;
	signal WX4279: std_logic; attribute dont_touch of WX4279: signal is true;
	signal WX4280: std_logic; attribute dont_touch of WX4280: signal is true;
	signal WX4281: std_logic; attribute dont_touch of WX4281: signal is true;
	signal WX4282: std_logic; attribute dont_touch of WX4282: signal is true;
	signal WX4283: std_logic; attribute dont_touch of WX4283: signal is true;
	signal WX4284: std_logic; attribute dont_touch of WX4284: signal is true;
	signal WX4285: std_logic; attribute dont_touch of WX4285: signal is true;
	signal WX4286: std_logic; attribute dont_touch of WX4286: signal is true;
	signal WX4287: std_logic; attribute dont_touch of WX4287: signal is true;
	signal WX4288: std_logic; attribute dont_touch of WX4288: signal is true;
	signal WX4289: std_logic; attribute dont_touch of WX4289: signal is true;
	signal WX4290: std_logic; attribute dont_touch of WX4290: signal is true;
	signal WX4291: std_logic; attribute dont_touch of WX4291: signal is true;
	signal WX4292: std_logic; attribute dont_touch of WX4292: signal is true;
	signal WX4293: std_logic; attribute dont_touch of WX4293: signal is true;
	signal WX4294: std_logic; attribute dont_touch of WX4294: signal is true;
	signal WX4295: std_logic; attribute dont_touch of WX4295: signal is true;
	signal WX4296: std_logic; attribute dont_touch of WX4296: signal is true;
	signal WX4297: std_logic; attribute dont_touch of WX4297: signal is true;
	signal WX4298: std_logic; attribute dont_touch of WX4298: signal is true;
	signal WX4299: std_logic; attribute dont_touch of WX4299: signal is true;
	signal WX4300: std_logic; attribute dont_touch of WX4300: signal is true;
	signal WX4301: std_logic; attribute dont_touch of WX4301: signal is true;
	signal WX4302: std_logic; attribute dont_touch of WX4302: signal is true;
	signal WX4303: std_logic; attribute dont_touch of WX4303: signal is true;
	signal WX4304: std_logic; attribute dont_touch of WX4304: signal is true;
	signal WX4305: std_logic; attribute dont_touch of WX4305: signal is true;
	signal WX4306: std_logic; attribute dont_touch of WX4306: signal is true;
	signal WX4307: std_logic; attribute dont_touch of WX4307: signal is true;
	signal WX4308: std_logic; attribute dont_touch of WX4308: signal is true;
	signal WX4309: std_logic; attribute dont_touch of WX4309: signal is true;
	signal WX4310: std_logic; attribute dont_touch of WX4310: signal is true;
	signal WX4311: std_logic; attribute dont_touch of WX4311: signal is true;
	signal WX4312: std_logic; attribute dont_touch of WX4312: signal is true;
	signal WX4313: std_logic; attribute dont_touch of WX4313: signal is true;
	signal WX4314: std_logic; attribute dont_touch of WX4314: signal is true;
	signal WX4315: std_logic; attribute dont_touch of WX4315: signal is true;
	signal WX4316: std_logic; attribute dont_touch of WX4316: signal is true;
	signal WX4317: std_logic; attribute dont_touch of WX4317: signal is true;
	signal WX4318: std_logic; attribute dont_touch of WX4318: signal is true;
	signal WX4319: std_logic; attribute dont_touch of WX4319: signal is true;
	signal WX4320: std_logic; attribute dont_touch of WX4320: signal is true;
	signal WX4321: std_logic; attribute dont_touch of WX4321: signal is true;
	signal WX4322: std_logic; attribute dont_touch of WX4322: signal is true;
	signal WX4323: std_logic; attribute dont_touch of WX4323: signal is true;
	signal WX4324: std_logic; attribute dont_touch of WX4324: signal is true;
	signal WX4325: std_logic; attribute dont_touch of WX4325: signal is true;
	signal WX4326: std_logic; attribute dont_touch of WX4326: signal is true;
	signal WX4327: std_logic; attribute dont_touch of WX4327: signal is true;
	signal WX4328: std_logic; attribute dont_touch of WX4328: signal is true;
	signal WX4329: std_logic; attribute dont_touch of WX4329: signal is true;
	signal WX4330: std_logic; attribute dont_touch of WX4330: signal is true;
	signal WX4331: std_logic; attribute dont_touch of WX4331: signal is true;
	signal WX4332: std_logic; attribute dont_touch of WX4332: signal is true;
	signal WX4333: std_logic; attribute dont_touch of WX4333: signal is true;
	signal WX4334: std_logic; attribute dont_touch of WX4334: signal is true;
	signal WX4335: std_logic; attribute dont_touch of WX4335: signal is true;
	signal WX4336: std_logic; attribute dont_touch of WX4336: signal is true;
	signal WX4337: std_logic; attribute dont_touch of WX4337: signal is true;
	signal WX4338: std_logic; attribute dont_touch of WX4338: signal is true;
	signal WX4339: std_logic; attribute dont_touch of WX4339: signal is true;
	signal WX4340: std_logic; attribute dont_touch of WX4340: signal is true;
	signal WX4341: std_logic; attribute dont_touch of WX4341: signal is true;
	signal WX4342: std_logic; attribute dont_touch of WX4342: signal is true;
	signal WX4343: std_logic; attribute dont_touch of WX4343: signal is true;
	signal WX4344: std_logic; attribute dont_touch of WX4344: signal is true;
	signal WX4345: std_logic; attribute dont_touch of WX4345: signal is true;
	signal WX4346: std_logic; attribute dont_touch of WX4346: signal is true;
	signal WX4347: std_logic; attribute dont_touch of WX4347: signal is true;
	signal WX4348: std_logic; attribute dont_touch of WX4348: signal is true;
	signal WX4349: std_logic; attribute dont_touch of WX4349: signal is true;
	signal WX4350: std_logic; attribute dont_touch of WX4350: signal is true;
	signal WX4351: std_logic; attribute dont_touch of WX4351: signal is true;
	signal WX4352: std_logic; attribute dont_touch of WX4352: signal is true;
	signal WX4353: std_logic; attribute dont_touch of WX4353: signal is true;
	signal WX4354: std_logic; attribute dont_touch of WX4354: signal is true;
	signal WX4355: std_logic; attribute dont_touch of WX4355: signal is true;
	signal WX4356: std_logic; attribute dont_touch of WX4356: signal is true;
	signal WX4357: std_logic; attribute dont_touch of WX4357: signal is true;
	signal WX4358: std_logic; attribute dont_touch of WX4358: signal is true;
	signal WX4359: std_logic; attribute dont_touch of WX4359: signal is true;
	signal WX4360: std_logic; attribute dont_touch of WX4360: signal is true;
	signal WX4361: std_logic; attribute dont_touch of WX4361: signal is true;
	signal WX4362: std_logic; attribute dont_touch of WX4362: signal is true;
	signal WX4363: std_logic; attribute dont_touch of WX4363: signal is true;
	signal WX4364: std_logic; attribute dont_touch of WX4364: signal is true;
	signal WX4365: std_logic; attribute dont_touch of WX4365: signal is true;
	signal WX4366: std_logic; attribute dont_touch of WX4366: signal is true;
	signal WX4367: std_logic; attribute dont_touch of WX4367: signal is true;
	signal WX4368: std_logic; attribute dont_touch of WX4368: signal is true;
	signal WX4369: std_logic; attribute dont_touch of WX4369: signal is true;
	signal WX4370: std_logic; attribute dont_touch of WX4370: signal is true;
	signal WX4371: std_logic; attribute dont_touch of WX4371: signal is true;
	signal WX4372: std_logic; attribute dont_touch of WX4372: signal is true;
	signal WX4373: std_logic; attribute dont_touch of WX4373: signal is true;
	signal WX4374: std_logic; attribute dont_touch of WX4374: signal is true;
	signal WX4375: std_logic; attribute dont_touch of WX4375: signal is true;
	signal WX4376: std_logic; attribute dont_touch of WX4376: signal is true;
	signal WX4377: std_logic; attribute dont_touch of WX4377: signal is true;
	signal WX4378: std_logic; attribute dont_touch of WX4378: signal is true;
	signal WX4379: std_logic; attribute dont_touch of WX4379: signal is true;
	signal WX4380: std_logic; attribute dont_touch of WX4380: signal is true;
	signal WX4381: std_logic; attribute dont_touch of WX4381: signal is true;
	signal WX4382: std_logic; attribute dont_touch of WX4382: signal is true;
	signal WX4383: std_logic; attribute dont_touch of WX4383: signal is true;
	signal WX4384: std_logic; attribute dont_touch of WX4384: signal is true;
	signal WX4385: std_logic; attribute dont_touch of WX4385: signal is true;
	signal WX4386: std_logic; attribute dont_touch of WX4386: signal is true;
	signal WX4387: std_logic; attribute dont_touch of WX4387: signal is true;
	signal WX4388: std_logic; attribute dont_touch of WX4388: signal is true;
	signal WX4389: std_logic; attribute dont_touch of WX4389: signal is true;
	signal WX4390: std_logic; attribute dont_touch of WX4390: signal is true;
	signal WX4391: std_logic; attribute dont_touch of WX4391: signal is true;
	signal WX4392: std_logic; attribute dont_touch of WX4392: signal is true;
	signal WX4393: std_logic; attribute dont_touch of WX4393: signal is true;
	signal WX4394: std_logic; attribute dont_touch of WX4394: signal is true;
	signal WX4395: std_logic; attribute dont_touch of WX4395: signal is true;
	signal WX4396: std_logic; attribute dont_touch of WX4396: signal is true;
	signal WX4397: std_logic; attribute dont_touch of WX4397: signal is true;
	signal WX4398: std_logic; attribute dont_touch of WX4398: signal is true;
	signal WX4399: std_logic; attribute dont_touch of WX4399: signal is true;
	signal WX4400: std_logic; attribute dont_touch of WX4400: signal is true;
	signal WX4401: std_logic; attribute dont_touch of WX4401: signal is true;
	signal WX4402: std_logic; attribute dont_touch of WX4402: signal is true;
	signal WX4403: std_logic; attribute dont_touch of WX4403: signal is true;
	signal WX4404: std_logic; attribute dont_touch of WX4404: signal is true;
	signal WX4405: std_logic; attribute dont_touch of WX4405: signal is true;
	signal WX4406: std_logic; attribute dont_touch of WX4406: signal is true;
	signal WX4407: std_logic; attribute dont_touch of WX4407: signal is true;
	signal WX4408: std_logic; attribute dont_touch of WX4408: signal is true;
	signal WX4409: std_logic; attribute dont_touch of WX4409: signal is true;
	signal WX4410: std_logic; attribute dont_touch of WX4410: signal is true;
	signal WX4411: std_logic; attribute dont_touch of WX4411: signal is true;
	signal WX4412: std_logic; attribute dont_touch of WX4412: signal is true;
	signal WX4413: std_logic; attribute dont_touch of WX4413: signal is true;
	signal WX4414: std_logic; attribute dont_touch of WX4414: signal is true;
	signal WX4415: std_logic; attribute dont_touch of WX4415: signal is true;
	signal WX4416: std_logic; attribute dont_touch of WX4416: signal is true;
	signal WX4417: std_logic; attribute dont_touch of WX4417: signal is true;
	signal WX4418: std_logic; attribute dont_touch of WX4418: signal is true;
	signal WX4419: std_logic; attribute dont_touch of WX4419: signal is true;
	signal WX4420: std_logic; attribute dont_touch of WX4420: signal is true;
	signal WX4421: std_logic; attribute dont_touch of WX4421: signal is true;
	signal WX4422: std_logic; attribute dont_touch of WX4422: signal is true;
	signal WX4423: std_logic; attribute dont_touch of WX4423: signal is true;
	signal WX4424: std_logic; attribute dont_touch of WX4424: signal is true;
	signal WX4425: std_logic; attribute dont_touch of WX4425: signal is true;
	signal WX4426: std_logic; attribute dont_touch of WX4426: signal is true;
	signal WX4427: std_logic; attribute dont_touch of WX4427: signal is true;
	signal WX4428: std_logic; attribute dont_touch of WX4428: signal is true;
	signal WX4429: std_logic; attribute dont_touch of WX4429: signal is true;
	signal WX4430: std_logic; attribute dont_touch of WX4430: signal is true;
	signal WX4431: std_logic; attribute dont_touch of WX4431: signal is true;
	signal WX4432: std_logic; attribute dont_touch of WX4432: signal is true;
	signal WX4433: std_logic; attribute dont_touch of WX4433: signal is true;
	signal WX4434: std_logic; attribute dont_touch of WX4434: signal is true;
	signal WX4435: std_logic; attribute dont_touch of WX4435: signal is true;
	signal WX4436: std_logic; attribute dont_touch of WX4436: signal is true;
	signal WX4437: std_logic; attribute dont_touch of WX4437: signal is true;
	signal WX4438: std_logic; attribute dont_touch of WX4438: signal is true;
	signal WX4439: std_logic; attribute dont_touch of WX4439: signal is true;
	signal WX4440: std_logic; attribute dont_touch of WX4440: signal is true;
	signal WX4441: std_logic; attribute dont_touch of WX4441: signal is true;
	signal WX4442: std_logic; attribute dont_touch of WX4442: signal is true;
	signal WX4443: std_logic; attribute dont_touch of WX4443: signal is true;
	signal WX4444: std_logic; attribute dont_touch of WX4444: signal is true;
	signal WX4445: std_logic; attribute dont_touch of WX4445: signal is true;
	signal WX4446: std_logic; attribute dont_touch of WX4446: signal is true;
	signal WX4447: std_logic; attribute dont_touch of WX4447: signal is true;
	signal WX4448: std_logic; attribute dont_touch of WX4448: signal is true;
	signal WX4449: std_logic; attribute dont_touch of WX4449: signal is true;
	signal WX4450: std_logic; attribute dont_touch of WX4450: signal is true;
	signal WX4451: std_logic; attribute dont_touch of WX4451: signal is true;
	signal WX4452: std_logic; attribute dont_touch of WX4452: signal is true;
	signal WX4453: std_logic; attribute dont_touch of WX4453: signal is true;
	signal WX4454: std_logic; attribute dont_touch of WX4454: signal is true;
	signal WX4455: std_logic; attribute dont_touch of WX4455: signal is true;
	signal WX4456: std_logic; attribute dont_touch of WX4456: signal is true;
	signal WX4457: std_logic; attribute dont_touch of WX4457: signal is true;
	signal WX4458: std_logic; attribute dont_touch of WX4458: signal is true;
	signal WX4459: std_logic; attribute dont_touch of WX4459: signal is true;
	signal WX4460: std_logic; attribute dont_touch of WX4460: signal is true;
	signal WX4461: std_logic; attribute dont_touch of WX4461: signal is true;
	signal WX4462: std_logic; attribute dont_touch of WX4462: signal is true;
	signal WX4463: std_logic; attribute dont_touch of WX4463: signal is true;
	signal WX4464: std_logic; attribute dont_touch of WX4464: signal is true;
	signal WX4465: std_logic; attribute dont_touch of WX4465: signal is true;
	signal WX4466: std_logic; attribute dont_touch of WX4466: signal is true;
	signal WX4467: std_logic; attribute dont_touch of WX4467: signal is true;
	signal WX4468: std_logic; attribute dont_touch of WX4468: signal is true;
	signal WX4469: std_logic; attribute dont_touch of WX4469: signal is true;
	signal WX4470: std_logic; attribute dont_touch of WX4470: signal is true;
	signal WX4471: std_logic; attribute dont_touch of WX4471: signal is true;
	signal WX4472: std_logic; attribute dont_touch of WX4472: signal is true;
	signal WX4473: std_logic; attribute dont_touch of WX4473: signal is true;
	signal WX4474: std_logic; attribute dont_touch of WX4474: signal is true;
	signal WX4475: std_logic; attribute dont_touch of WX4475: signal is true;
	signal WX4476: std_logic; attribute dont_touch of WX4476: signal is true;
	signal WX4477: std_logic; attribute dont_touch of WX4477: signal is true;
	signal WX4478: std_logic; attribute dont_touch of WX4478: signal is true;
	signal WX4479: std_logic; attribute dont_touch of WX4479: signal is true;
	signal WX4480: std_logic; attribute dont_touch of WX4480: signal is true;
	signal WX4481: std_logic; attribute dont_touch of WX4481: signal is true;
	signal WX4482: std_logic; attribute dont_touch of WX4482: signal is true;
	signal WX4483: std_logic; attribute dont_touch of WX4483: signal is true;
	signal WX4484: std_logic; attribute dont_touch of WX4484: signal is true;
	signal WX4485: std_logic; attribute dont_touch of WX4485: signal is true;
	signal WX4486: std_logic; attribute dont_touch of WX4486: signal is true;
	signal WX4487: std_logic; attribute dont_touch of WX4487: signal is true;
	signal WX4488: std_logic; attribute dont_touch of WX4488: signal is true;
	signal WX4489: std_logic; attribute dont_touch of WX4489: signal is true;
	signal WX4490: std_logic; attribute dont_touch of WX4490: signal is true;
	signal WX4491: std_logic; attribute dont_touch of WX4491: signal is true;
	signal WX4492: std_logic; attribute dont_touch of WX4492: signal is true;
	signal WX4493: std_logic; attribute dont_touch of WX4493: signal is true;
	signal WX4494: std_logic; attribute dont_touch of WX4494: signal is true;
	signal WX4495: std_logic; attribute dont_touch of WX4495: signal is true;
	signal WX4496: std_logic; attribute dont_touch of WX4496: signal is true;
	signal WX4497: std_logic; attribute dont_touch of WX4497: signal is true;
	signal WX4498: std_logic; attribute dont_touch of WX4498: signal is true;
	signal WX4499: std_logic; attribute dont_touch of WX4499: signal is true;
	signal WX4500: std_logic; attribute dont_touch of WX4500: signal is true;
	signal WX4501: std_logic; attribute dont_touch of WX4501: signal is true;
	signal WX4502: std_logic; attribute dont_touch of WX4502: signal is true;
	signal WX4503: std_logic; attribute dont_touch of WX4503: signal is true;
	signal WX4504: std_logic; attribute dont_touch of WX4504: signal is true;
	signal WX4505: std_logic; attribute dont_touch of WX4505: signal is true;
	signal WX4506: std_logic; attribute dont_touch of WX4506: signal is true;
	signal WX4507: std_logic; attribute dont_touch of WX4507: signal is true;
	signal WX4508: std_logic; attribute dont_touch of WX4508: signal is true;
	signal WX4509: std_logic; attribute dont_touch of WX4509: signal is true;
	signal WX4510: std_logic; attribute dont_touch of WX4510: signal is true;
	signal WX4511: std_logic; attribute dont_touch of WX4511: signal is true;
	signal WX4512: std_logic; attribute dont_touch of WX4512: signal is true;
	signal WX4513: std_logic; attribute dont_touch of WX4513: signal is true;
	signal WX4514: std_logic; attribute dont_touch of WX4514: signal is true;
	signal WX4515: std_logic; attribute dont_touch of WX4515: signal is true;
	signal WX4516: std_logic; attribute dont_touch of WX4516: signal is true;
	signal WX4517: std_logic; attribute dont_touch of WX4517: signal is true;
	signal WX4518: std_logic; attribute dont_touch of WX4518: signal is true;
	signal WX4519: std_logic; attribute dont_touch of WX4519: signal is true;
	signal WX4520: std_logic; attribute dont_touch of WX4520: signal is true;
	signal WX4521: std_logic; attribute dont_touch of WX4521: signal is true;
	signal WX4522: std_logic; attribute dont_touch of WX4522: signal is true;
	signal WX4523: std_logic; attribute dont_touch of WX4523: signal is true;
	signal WX4524: std_logic; attribute dont_touch of WX4524: signal is true;
	signal WX4525: std_logic; attribute dont_touch of WX4525: signal is true;
	signal WX4526: std_logic; attribute dont_touch of WX4526: signal is true;
	signal WX4527: std_logic; attribute dont_touch of WX4527: signal is true;
	signal WX4528: std_logic; attribute dont_touch of WX4528: signal is true;
	signal WX4529: std_logic; attribute dont_touch of WX4529: signal is true;
	signal WX4530: std_logic; attribute dont_touch of WX4530: signal is true;
	signal WX4531: std_logic; attribute dont_touch of WX4531: signal is true;
	signal WX4532: std_logic; attribute dont_touch of WX4532: signal is true;
	signal WX4533: std_logic; attribute dont_touch of WX4533: signal is true;
	signal WX4534: std_logic; attribute dont_touch of WX4534: signal is true;
	signal WX4535: std_logic; attribute dont_touch of WX4535: signal is true;
	signal WX4536: std_logic; attribute dont_touch of WX4536: signal is true;
	signal WX4537: std_logic; attribute dont_touch of WX4537: signal is true;
	signal WX4538: std_logic; attribute dont_touch of WX4538: signal is true;
	signal WX4539: std_logic; attribute dont_touch of WX4539: signal is true;
	signal WX4540: std_logic; attribute dont_touch of WX4540: signal is true;
	signal WX4541: std_logic; attribute dont_touch of WX4541: signal is true;
	signal WX4542: std_logic; attribute dont_touch of WX4542: signal is true;
	signal WX4543: std_logic; attribute dont_touch of WX4543: signal is true;
	signal WX4544: std_logic; attribute dont_touch of WX4544: signal is true;
	signal WX4545: std_logic; attribute dont_touch of WX4545: signal is true;
	signal WX4546: std_logic; attribute dont_touch of WX4546: signal is true;
	signal WX4547: std_logic; attribute dont_touch of WX4547: signal is true;
	signal WX4548: std_logic; attribute dont_touch of WX4548: signal is true;
	signal WX4549: std_logic; attribute dont_touch of WX4549: signal is true;
	signal WX4550: std_logic; attribute dont_touch of WX4550: signal is true;
	signal WX4551: std_logic; attribute dont_touch of WX4551: signal is true;
	signal WX4552: std_logic; attribute dont_touch of WX4552: signal is true;
	signal WX4553: std_logic; attribute dont_touch of WX4553: signal is true;
	signal WX4554: std_logic; attribute dont_touch of WX4554: signal is true;
	signal WX4555: std_logic; attribute dont_touch of WX4555: signal is true;
	signal WX4556: std_logic; attribute dont_touch of WX4556: signal is true;
	signal WX4557: std_logic; attribute dont_touch of WX4557: signal is true;
	signal WX4558: std_logic; attribute dont_touch of WX4558: signal is true;
	signal WX4559: std_logic; attribute dont_touch of WX4559: signal is true;
	signal WX4560: std_logic; attribute dont_touch of WX4560: signal is true;
	signal WX4561: std_logic; attribute dont_touch of WX4561: signal is true;
	signal WX4562: std_logic; attribute dont_touch of WX4562: signal is true;
	signal WX4563: std_logic; attribute dont_touch of WX4563: signal is true;
	signal WX4564: std_logic; attribute dont_touch of WX4564: signal is true;
	signal WX4565: std_logic; attribute dont_touch of WX4565: signal is true;
	signal WX4566: std_logic; attribute dont_touch of WX4566: signal is true;
	signal WX4567: std_logic; attribute dont_touch of WX4567: signal is true;
	signal WX4568: std_logic; attribute dont_touch of WX4568: signal is true;
	signal WX4569: std_logic; attribute dont_touch of WX4569: signal is true;
	signal WX4570: std_logic; attribute dont_touch of WX4570: signal is true;
	signal WX4571: std_logic; attribute dont_touch of WX4571: signal is true;
	signal WX4572: std_logic; attribute dont_touch of WX4572: signal is true;
	signal WX4573: std_logic; attribute dont_touch of WX4573: signal is true;
	signal WX4574: std_logic; attribute dont_touch of WX4574: signal is true;
	signal WX4575: std_logic; attribute dont_touch of WX4575: signal is true;
	signal WX4576: std_logic; attribute dont_touch of WX4576: signal is true;
	signal WX4577: std_logic; attribute dont_touch of WX4577: signal is true;
	signal WX4578: std_logic; attribute dont_touch of WX4578: signal is true;
	signal WX4579: std_logic; attribute dont_touch of WX4579: signal is true;
	signal WX4580: std_logic; attribute dont_touch of WX4580: signal is true;
	signal WX4581: std_logic; attribute dont_touch of WX4581: signal is true;
	signal WX4582: std_logic; attribute dont_touch of WX4582: signal is true;
	signal WX4583: std_logic; attribute dont_touch of WX4583: signal is true;
	signal WX4584: std_logic; attribute dont_touch of WX4584: signal is true;
	signal WX4585: std_logic; attribute dont_touch of WX4585: signal is true;
	signal WX4586: std_logic; attribute dont_touch of WX4586: signal is true;
	signal WX4587: std_logic; attribute dont_touch of WX4587: signal is true;
	signal WX4588: std_logic; attribute dont_touch of WX4588: signal is true;
	signal WX4589: std_logic; attribute dont_touch of WX4589: signal is true;
	signal WX4590: std_logic; attribute dont_touch of WX4590: signal is true;
	signal WX4591: std_logic; attribute dont_touch of WX4591: signal is true;
	signal WX4592: std_logic; attribute dont_touch of WX4592: signal is true;
	signal WX4593: std_logic; attribute dont_touch of WX4593: signal is true;
	signal WX4594: std_logic; attribute dont_touch of WX4594: signal is true;
	signal WX4595: std_logic; attribute dont_touch of WX4595: signal is true;
	signal WX4596: std_logic; attribute dont_touch of WX4596: signal is true;
	signal WX4597: std_logic; attribute dont_touch of WX4597: signal is true;
	signal WX4598: std_logic; attribute dont_touch of WX4598: signal is true;
	signal WX4599: std_logic; attribute dont_touch of WX4599: signal is true;
	signal WX4600: std_logic; attribute dont_touch of WX4600: signal is true;
	signal WX4601: std_logic; attribute dont_touch of WX4601: signal is true;
	signal WX4602: std_logic; attribute dont_touch of WX4602: signal is true;
	signal WX4603: std_logic; attribute dont_touch of WX4603: signal is true;
	signal WX4604: std_logic; attribute dont_touch of WX4604: signal is true;
	signal WX4605: std_logic; attribute dont_touch of WX4605: signal is true;
	signal WX4606: std_logic; attribute dont_touch of WX4606: signal is true;
	signal WX4607: std_logic; attribute dont_touch of WX4607: signal is true;
	signal WX4608: std_logic; attribute dont_touch of WX4608: signal is true;
	signal WX4609: std_logic; attribute dont_touch of WX4609: signal is true;
	signal WX4610: std_logic; attribute dont_touch of WX4610: signal is true;
	signal WX4611: std_logic; attribute dont_touch of WX4611: signal is true;
	signal WX4612: std_logic; attribute dont_touch of WX4612: signal is true;
	signal WX4613: std_logic; attribute dont_touch of WX4613: signal is true;
	signal WX4614: std_logic; attribute dont_touch of WX4614: signal is true;
	signal WX4615: std_logic; attribute dont_touch of WX4615: signal is true;
	signal WX4616: std_logic; attribute dont_touch of WX4616: signal is true;
	signal WX4617: std_logic; attribute dont_touch of WX4617: signal is true;
	signal WX4618: std_logic; attribute dont_touch of WX4618: signal is true;
	signal WX4619: std_logic; attribute dont_touch of WX4619: signal is true;
	signal WX4620: std_logic; attribute dont_touch of WX4620: signal is true;
	signal WX4621: std_logic; attribute dont_touch of WX4621: signal is true;
	signal WX4622: std_logic; attribute dont_touch of WX4622: signal is true;
	signal WX4623: std_logic; attribute dont_touch of WX4623: signal is true;
	signal WX4624: std_logic; attribute dont_touch of WX4624: signal is true;
	signal WX4625: std_logic; attribute dont_touch of WX4625: signal is true;
	signal WX4626: std_logic; attribute dont_touch of WX4626: signal is true;
	signal WX4627: std_logic; attribute dont_touch of WX4627: signal is true;
	signal WX4628: std_logic; attribute dont_touch of WX4628: signal is true;
	signal WX4629: std_logic; attribute dont_touch of WX4629: signal is true;
	signal WX4630: std_logic; attribute dont_touch of WX4630: signal is true;
	signal WX4631: std_logic; attribute dont_touch of WX4631: signal is true;
	signal WX4632: std_logic; attribute dont_touch of WX4632: signal is true;
	signal WX4633: std_logic; attribute dont_touch of WX4633: signal is true;
	signal WX4634: std_logic; attribute dont_touch of WX4634: signal is true;
	signal WX4635: std_logic; attribute dont_touch of WX4635: signal is true;
	signal WX4636: std_logic; attribute dont_touch of WX4636: signal is true;
	signal WX4637: std_logic; attribute dont_touch of WX4637: signal is true;
	signal WX4638: std_logic; attribute dont_touch of WX4638: signal is true;
	signal WX4639: std_logic; attribute dont_touch of WX4639: signal is true;
	signal WX4640: std_logic; attribute dont_touch of WX4640: signal is true;
	signal WX4641: std_logic; attribute dont_touch of WX4641: signal is true;
	signal WX4642: std_logic; attribute dont_touch of WX4642: signal is true;
	signal WX4643: std_logic; attribute dont_touch of WX4643: signal is true;
	signal WX4644: std_logic; attribute dont_touch of WX4644: signal is true;
	signal WX4645: std_logic; attribute dont_touch of WX4645: signal is true;
	signal WX4646: std_logic; attribute dont_touch of WX4646: signal is true;
	signal WX4647: std_logic; attribute dont_touch of WX4647: signal is true;
	signal WX4648: std_logic; attribute dont_touch of WX4648: signal is true;
	signal WX4649: std_logic; attribute dont_touch of WX4649: signal is true;
	signal WX4650: std_logic; attribute dont_touch of WX4650: signal is true;
	signal WX4651: std_logic; attribute dont_touch of WX4651: signal is true;
	signal WX4652: std_logic; attribute dont_touch of WX4652: signal is true;
	signal WX4653: std_logic; attribute dont_touch of WX4653: signal is true;
	signal WX4654: std_logic; attribute dont_touch of WX4654: signal is true;
	signal WX4655: std_logic; attribute dont_touch of WX4655: signal is true;
	signal WX4656: std_logic; attribute dont_touch of WX4656: signal is true;
	signal WX4657: std_logic; attribute dont_touch of WX4657: signal is true;
	signal WX4658: std_logic; attribute dont_touch of WX4658: signal is true;
	signal WX4659: std_logic; attribute dont_touch of WX4659: signal is true;
	signal WX4660: std_logic; attribute dont_touch of WX4660: signal is true;
	signal WX4661: std_logic; attribute dont_touch of WX4661: signal is true;
	signal WX4662: std_logic; attribute dont_touch of WX4662: signal is true;
	signal WX4663: std_logic; attribute dont_touch of WX4663: signal is true;
	signal WX4664: std_logic; attribute dont_touch of WX4664: signal is true;
	signal WX4665: std_logic; attribute dont_touch of WX4665: signal is true;
	signal WX4666: std_logic; attribute dont_touch of WX4666: signal is true;
	signal WX4667: std_logic; attribute dont_touch of WX4667: signal is true;
	signal WX4668: std_logic; attribute dont_touch of WX4668: signal is true;
	signal WX4669: std_logic; attribute dont_touch of WX4669: signal is true;
	signal WX4670: std_logic; attribute dont_touch of WX4670: signal is true;
	signal WX4671: std_logic; attribute dont_touch of WX4671: signal is true;
	signal WX4672: std_logic; attribute dont_touch of WX4672: signal is true;
	signal WX4673: std_logic; attribute dont_touch of WX4673: signal is true;
	signal WX4674: std_logic; attribute dont_touch of WX4674: signal is true;
	signal WX4675: std_logic; attribute dont_touch of WX4675: signal is true;
	signal WX4676: std_logic; attribute dont_touch of WX4676: signal is true;
	signal WX4677: std_logic; attribute dont_touch of WX4677: signal is true;
	signal WX4678: std_logic; attribute dont_touch of WX4678: signal is true;
	signal WX4679: std_logic; attribute dont_touch of WX4679: signal is true;
	signal WX4680: std_logic; attribute dont_touch of WX4680: signal is true;
	signal WX4681: std_logic; attribute dont_touch of WX4681: signal is true;
	signal WX4682: std_logic; attribute dont_touch of WX4682: signal is true;
	signal WX4683: std_logic; attribute dont_touch of WX4683: signal is true;
	signal WX4684: std_logic; attribute dont_touch of WX4684: signal is true;
	signal WX4685: std_logic; attribute dont_touch of WX4685: signal is true;
	signal WX4686: std_logic; attribute dont_touch of WX4686: signal is true;
	signal WX4687: std_logic; attribute dont_touch of WX4687: signal is true;
	signal WX4688: std_logic; attribute dont_touch of WX4688: signal is true;
	signal WX4689: std_logic; attribute dont_touch of WX4689: signal is true;
	signal WX4690: std_logic; attribute dont_touch of WX4690: signal is true;
	signal WX4691: std_logic; attribute dont_touch of WX4691: signal is true;
	signal WX4692: std_logic; attribute dont_touch of WX4692: signal is true;
	signal WX4693: std_logic; attribute dont_touch of WX4693: signal is true;
	signal WX4694: std_logic; attribute dont_touch of WX4694: signal is true;
	signal WX4695: std_logic; attribute dont_touch of WX4695: signal is true;
	signal WX4696: std_logic; attribute dont_touch of WX4696: signal is true;
	signal WX4697: std_logic; attribute dont_touch of WX4697: signal is true;
	signal WX4698: std_logic; attribute dont_touch of WX4698: signal is true;
	signal WX4699: std_logic; attribute dont_touch of WX4699: signal is true;
	signal WX4700: std_logic; attribute dont_touch of WX4700: signal is true;
	signal WX4701: std_logic; attribute dont_touch of WX4701: signal is true;
	signal WX4702: std_logic; attribute dont_touch of WX4702: signal is true;
	signal WX4703: std_logic; attribute dont_touch of WX4703: signal is true;
	signal WX4704: std_logic; attribute dont_touch of WX4704: signal is true;
	signal WX4705: std_logic; attribute dont_touch of WX4705: signal is true;
	signal WX4706: std_logic; attribute dont_touch of WX4706: signal is true;
	signal WX4707: std_logic; attribute dont_touch of WX4707: signal is true;
	signal WX4708: std_logic; attribute dont_touch of WX4708: signal is true;
	signal WX4709: std_logic; attribute dont_touch of WX4709: signal is true;
	signal WX4710: std_logic; attribute dont_touch of WX4710: signal is true;
	signal WX4711: std_logic; attribute dont_touch of WX4711: signal is true;
	signal WX4712: std_logic; attribute dont_touch of WX4712: signal is true;
	signal WX4713: std_logic; attribute dont_touch of WX4713: signal is true;
	signal WX4714: std_logic; attribute dont_touch of WX4714: signal is true;
	signal WX4715: std_logic; attribute dont_touch of WX4715: signal is true;
	signal WX4716: std_logic; attribute dont_touch of WX4716: signal is true;
	signal WX4717: std_logic; attribute dont_touch of WX4717: signal is true;
	signal WX4718: std_logic; attribute dont_touch of WX4718: signal is true;
	signal WX4719: std_logic; attribute dont_touch of WX4719: signal is true;
	signal WX4720: std_logic; attribute dont_touch of WX4720: signal is true;
	signal WX4721: std_logic; attribute dont_touch of WX4721: signal is true;
	signal WX4722: std_logic; attribute dont_touch of WX4722: signal is true;
	signal WX4723: std_logic; attribute dont_touch of WX4723: signal is true;
	signal WX4724: std_logic; attribute dont_touch of WX4724: signal is true;
	signal WX4725: std_logic; attribute dont_touch of WX4725: signal is true;
	signal WX4726: std_logic; attribute dont_touch of WX4726: signal is true;
	signal WX4727: std_logic; attribute dont_touch of WX4727: signal is true;
	signal WX4728: std_logic; attribute dont_touch of WX4728: signal is true;
	signal WX4729: std_logic; attribute dont_touch of WX4729: signal is true;
	signal WX4730: std_logic; attribute dont_touch of WX4730: signal is true;
	signal WX4731: std_logic; attribute dont_touch of WX4731: signal is true;
	signal WX4732: std_logic; attribute dont_touch of WX4732: signal is true;
	signal WX4733: std_logic; attribute dont_touch of WX4733: signal is true;
	signal WX4734: std_logic; attribute dont_touch of WX4734: signal is true;
	signal WX4735: std_logic; attribute dont_touch of WX4735: signal is true;
	signal WX4736: std_logic; attribute dont_touch of WX4736: signal is true;
	signal WX4737: std_logic; attribute dont_touch of WX4737: signal is true;
	signal WX4738: std_logic; attribute dont_touch of WX4738: signal is true;
	signal WX4739: std_logic; attribute dont_touch of WX4739: signal is true;
	signal WX4740: std_logic; attribute dont_touch of WX4740: signal is true;
	signal WX4741: std_logic; attribute dont_touch of WX4741: signal is true;
	signal WX4742: std_logic; attribute dont_touch of WX4742: signal is true;
	signal WX4743: std_logic; attribute dont_touch of WX4743: signal is true;
	signal WX4744: std_logic; attribute dont_touch of WX4744: signal is true;
	signal WX4745: std_logic; attribute dont_touch of WX4745: signal is true;
	signal WX4746: std_logic; attribute dont_touch of WX4746: signal is true;
	signal WX4747: std_logic; attribute dont_touch of WX4747: signal is true;
	signal WX4748: std_logic; attribute dont_touch of WX4748: signal is true;
	signal WX4749: std_logic; attribute dont_touch of WX4749: signal is true;
	signal WX4750: std_logic; attribute dont_touch of WX4750: signal is true;
	signal WX4751: std_logic; attribute dont_touch of WX4751: signal is true;
	signal WX4752: std_logic; attribute dont_touch of WX4752: signal is true;
	signal WX4753: std_logic; attribute dont_touch of WX4753: signal is true;
	signal WX4754: std_logic; attribute dont_touch of WX4754: signal is true;
	signal WX4755: std_logic; attribute dont_touch of WX4755: signal is true;
	signal WX4756: std_logic; attribute dont_touch of WX4756: signal is true;
	signal WX4757: std_logic; attribute dont_touch of WX4757: signal is true;
	signal WX4758: std_logic; attribute dont_touch of WX4758: signal is true;
	signal WX4759: std_logic; attribute dont_touch of WX4759: signal is true;
	signal WX4760: std_logic; attribute dont_touch of WX4760: signal is true;
	signal WX4761: std_logic; attribute dont_touch of WX4761: signal is true;
	signal WX4762: std_logic; attribute dont_touch of WX4762: signal is true;
	signal WX4763: std_logic; attribute dont_touch of WX4763: signal is true;
	signal WX4764: std_logic; attribute dont_touch of WX4764: signal is true;
	signal WX4765: std_logic; attribute dont_touch of WX4765: signal is true;
	signal WX4766: std_logic; attribute dont_touch of WX4766: signal is true;
	signal WX4767: std_logic; attribute dont_touch of WX4767: signal is true;
	signal WX4768: std_logic; attribute dont_touch of WX4768: signal is true;
	signal WX4769: std_logic; attribute dont_touch of WX4769: signal is true;
	signal WX4770: std_logic; attribute dont_touch of WX4770: signal is true;
	signal WX4771: std_logic; attribute dont_touch of WX4771: signal is true;
	signal WX4772: std_logic; attribute dont_touch of WX4772: signal is true;
	signal WX4773: std_logic; attribute dont_touch of WX4773: signal is true;
	signal WX4774: std_logic; attribute dont_touch of WX4774: signal is true;
	signal WX4775: std_logic; attribute dont_touch of WX4775: signal is true;
	signal WX4776: std_logic; attribute dont_touch of WX4776: signal is true;
	signal WX4777: std_logic; attribute dont_touch of WX4777: signal is true;
	signal WX4778: std_logic; attribute dont_touch of WX4778: signal is true;
	signal WX4779: std_logic; attribute dont_touch of WX4779: signal is true;
	signal WX4780: std_logic; attribute dont_touch of WX4780: signal is true;
	signal WX4781: std_logic; attribute dont_touch of WX4781: signal is true;
	signal WX4782: std_logic; attribute dont_touch of WX4782: signal is true;
	signal WX4783: std_logic; attribute dont_touch of WX4783: signal is true;
	signal WX4784: std_logic; attribute dont_touch of WX4784: signal is true;
	signal WX4785: std_logic; attribute dont_touch of WX4785: signal is true;
	signal WX4786: std_logic; attribute dont_touch of WX4786: signal is true;
	signal WX4787: std_logic; attribute dont_touch of WX4787: signal is true;
	signal WX4788: std_logic; attribute dont_touch of WX4788: signal is true;
	signal WX4789: std_logic; attribute dont_touch of WX4789: signal is true;
	signal WX4790: std_logic; attribute dont_touch of WX4790: signal is true;
	signal WX4791: std_logic; attribute dont_touch of WX4791: signal is true;
	signal WX4792: std_logic; attribute dont_touch of WX4792: signal is true;
	signal WX4793: std_logic; attribute dont_touch of WX4793: signal is true;
	signal WX4794: std_logic; attribute dont_touch of WX4794: signal is true;
	signal WX4795: std_logic; attribute dont_touch of WX4795: signal is true;
	signal WX4796: std_logic; attribute dont_touch of WX4796: signal is true;
	signal WX4797: std_logic; attribute dont_touch of WX4797: signal is true;
	signal WX4798: std_logic; attribute dont_touch of WX4798: signal is true;
	signal WX4799: std_logic; attribute dont_touch of WX4799: signal is true;
	signal WX4800: std_logic; attribute dont_touch of WX4800: signal is true;
	signal WX4801: std_logic; attribute dont_touch of WX4801: signal is true;
	signal WX4802: std_logic; attribute dont_touch of WX4802: signal is true;
	signal WX4803: std_logic; attribute dont_touch of WX4803: signal is true;
	signal WX4804: std_logic; attribute dont_touch of WX4804: signal is true;
	signal WX4805: std_logic; attribute dont_touch of WX4805: signal is true;
	signal WX4806: std_logic; attribute dont_touch of WX4806: signal is true;
	signal WX4807: std_logic; attribute dont_touch of WX4807: signal is true;
	signal WX4808: std_logic; attribute dont_touch of WX4808: signal is true;
	signal WX4809: std_logic; attribute dont_touch of WX4809: signal is true;
	signal WX4810: std_logic; attribute dont_touch of WX4810: signal is true;
	signal WX4811: std_logic; attribute dont_touch of WX4811: signal is true;
	signal WX4812: std_logic; attribute dont_touch of WX4812: signal is true;
	signal WX4813: std_logic; attribute dont_touch of WX4813: signal is true;
	signal WX4814: std_logic; attribute dont_touch of WX4814: signal is true;
	signal WX4815: std_logic; attribute dont_touch of WX4815: signal is true;
	signal WX4816: std_logic; attribute dont_touch of WX4816: signal is true;
	signal WX4817: std_logic; attribute dont_touch of WX4817: signal is true;
	signal WX4818: std_logic; attribute dont_touch of WX4818: signal is true;
	signal WX4819: std_logic; attribute dont_touch of WX4819: signal is true;
	signal WX4820: std_logic; attribute dont_touch of WX4820: signal is true;
	signal WX4821: std_logic; attribute dont_touch of WX4821: signal is true;
	signal WX4822: std_logic; attribute dont_touch of WX4822: signal is true;
	signal WX4823: std_logic; attribute dont_touch of WX4823: signal is true;
	signal WX4824: std_logic; attribute dont_touch of WX4824: signal is true;
	signal WX4825: std_logic; attribute dont_touch of WX4825: signal is true;
	signal WX4826: std_logic; attribute dont_touch of WX4826: signal is true;
	signal WX4827: std_logic; attribute dont_touch of WX4827: signal is true;
	signal WX4828: std_logic; attribute dont_touch of WX4828: signal is true;
	signal WX4829: std_logic; attribute dont_touch of WX4829: signal is true;
	signal WX4830: std_logic; attribute dont_touch of WX4830: signal is true;
	signal WX4831: std_logic; attribute dont_touch of WX4831: signal is true;
	signal WX4832: std_logic; attribute dont_touch of WX4832: signal is true;
	signal WX4833: std_logic; attribute dont_touch of WX4833: signal is true;
	signal WX4834: std_logic; attribute dont_touch of WX4834: signal is true;
	signal WX4835: std_logic; attribute dont_touch of WX4835: signal is true;
	signal WX4836: std_logic; attribute dont_touch of WX4836: signal is true;
	signal WX4837: std_logic; attribute dont_touch of WX4837: signal is true;
	signal WX4838: std_logic; attribute dont_touch of WX4838: signal is true;
	signal WX4839: std_logic; attribute dont_touch of WX4839: signal is true;
	signal WX4840: std_logic; attribute dont_touch of WX4840: signal is true;
	signal WX4841: std_logic; attribute dont_touch of WX4841: signal is true;
	signal WX4842: std_logic; attribute dont_touch of WX4842: signal is true;
	signal WX4843: std_logic; attribute dont_touch of WX4843: signal is true;
	signal WX4844: std_logic; attribute dont_touch of WX4844: signal is true;
	signal WX4845: std_logic; attribute dont_touch of WX4845: signal is true;
	signal WX4846: std_logic; attribute dont_touch of WX4846: signal is true;
	signal WX4847: std_logic; attribute dont_touch of WX4847: signal is true;
	signal WX4848: std_logic; attribute dont_touch of WX4848: signal is true;
	signal WX4849: std_logic; attribute dont_touch of WX4849: signal is true;
	signal WX4850: std_logic; attribute dont_touch of WX4850: signal is true;
	signal WX4851: std_logic; attribute dont_touch of WX4851: signal is true;
	signal WX4852: std_logic; attribute dont_touch of WX4852: signal is true;
	signal WX4853: std_logic; attribute dont_touch of WX4853: signal is true;
	signal WX4854: std_logic; attribute dont_touch of WX4854: signal is true;
	signal WX4855: std_logic; attribute dont_touch of WX4855: signal is true;
	signal WX4856: std_logic; attribute dont_touch of WX4856: signal is true;
	signal WX4857: std_logic; attribute dont_touch of WX4857: signal is true;
	signal WX4858: std_logic; attribute dont_touch of WX4858: signal is true;
	signal WX4859: std_logic; attribute dont_touch of WX4859: signal is true;
	signal WX4860: std_logic; attribute dont_touch of WX4860: signal is true;
	signal WX4861: std_logic; attribute dont_touch of WX4861: signal is true;
	signal WX4862: std_logic; attribute dont_touch of WX4862: signal is true;
	signal WX4863: std_logic; attribute dont_touch of WX4863: signal is true;
	signal WX4864: std_logic; attribute dont_touch of WX4864: signal is true;
	signal WX4865: std_logic; attribute dont_touch of WX4865: signal is true;
	signal WX4866: std_logic; attribute dont_touch of WX4866: signal is true;
	signal WX4867: std_logic; attribute dont_touch of WX4867: signal is true;
	signal WX4868: std_logic; attribute dont_touch of WX4868: signal is true;
	signal WX4869: std_logic; attribute dont_touch of WX4869: signal is true;
	signal WX4870: std_logic; attribute dont_touch of WX4870: signal is true;
	signal WX4871: std_logic; attribute dont_touch of WX4871: signal is true;
	signal WX4872: std_logic; attribute dont_touch of WX4872: signal is true;
	signal WX4873: std_logic; attribute dont_touch of WX4873: signal is true;
	signal WX4874: std_logic; attribute dont_touch of WX4874: signal is true;
	signal WX4875: std_logic; attribute dont_touch of WX4875: signal is true;
	signal WX4876: std_logic; attribute dont_touch of WX4876: signal is true;
	signal WX4877: std_logic; attribute dont_touch of WX4877: signal is true;
	signal WX4878: std_logic; attribute dont_touch of WX4878: signal is true;
	signal WX4879: std_logic; attribute dont_touch of WX4879: signal is true;
	signal WX4880: std_logic; attribute dont_touch of WX4880: signal is true;
	signal WX4881: std_logic; attribute dont_touch of WX4881: signal is true;
	signal WX4882: std_logic; attribute dont_touch of WX4882: signal is true;
	signal WX4883: std_logic; attribute dont_touch of WX4883: signal is true;
	signal WX4884: std_logic; attribute dont_touch of WX4884: signal is true;
	signal WX4885: std_logic; attribute dont_touch of WX4885: signal is true;
	signal WX4886: std_logic; attribute dont_touch of WX4886: signal is true;
	signal WX4887: std_logic; attribute dont_touch of WX4887: signal is true;
	signal WX4888: std_logic; attribute dont_touch of WX4888: signal is true;
	signal WX4889: std_logic; attribute dont_touch of WX4889: signal is true;
	signal WX4890: std_logic; attribute dont_touch of WX4890: signal is true;
	signal WX4891: std_logic; attribute dont_touch of WX4891: signal is true;
	signal WX4892: std_logic; attribute dont_touch of WX4892: signal is true;
	signal WX4893: std_logic; attribute dont_touch of WX4893: signal is true;
	signal WX4894: std_logic; attribute dont_touch of WX4894: signal is true;
	signal WX4895: std_logic; attribute dont_touch of WX4895: signal is true;
	signal WX4896: std_logic; attribute dont_touch of WX4896: signal is true;
	signal WX4897: std_logic; attribute dont_touch of WX4897: signal is true;
	signal WX4898: std_logic; attribute dont_touch of WX4898: signal is true;
	signal WX4899: std_logic; attribute dont_touch of WX4899: signal is true;
	signal WX4900: std_logic; attribute dont_touch of WX4900: signal is true;
	signal WX4901: std_logic; attribute dont_touch of WX4901: signal is true;
	signal WX4902: std_logic; attribute dont_touch of WX4902: signal is true;
	signal WX4903: std_logic; attribute dont_touch of WX4903: signal is true;
	signal WX4904: std_logic; attribute dont_touch of WX4904: signal is true;
	signal WX4905: std_logic; attribute dont_touch of WX4905: signal is true;
	signal WX4906: std_logic; attribute dont_touch of WX4906: signal is true;
	signal WX4907: std_logic; attribute dont_touch of WX4907: signal is true;
	signal WX4908: std_logic; attribute dont_touch of WX4908: signal is true;
	signal WX4909: std_logic; attribute dont_touch of WX4909: signal is true;
	signal WX4910: std_logic; attribute dont_touch of WX4910: signal is true;
	signal WX4911: std_logic; attribute dont_touch of WX4911: signal is true;
	signal WX4912: std_logic; attribute dont_touch of WX4912: signal is true;
	signal WX4913: std_logic; attribute dont_touch of WX4913: signal is true;
	signal WX4914: std_logic; attribute dont_touch of WX4914: signal is true;
	signal WX4915: std_logic; attribute dont_touch of WX4915: signal is true;
	signal WX4916: std_logic; attribute dont_touch of WX4916: signal is true;
	signal WX4917: std_logic; attribute dont_touch of WX4917: signal is true;
	signal WX4918: std_logic; attribute dont_touch of WX4918: signal is true;
	signal WX4919: std_logic; attribute dont_touch of WX4919: signal is true;
	signal WX4920: std_logic; attribute dont_touch of WX4920: signal is true;
	signal WX4921: std_logic; attribute dont_touch of WX4921: signal is true;
	signal WX4922: std_logic; attribute dont_touch of WX4922: signal is true;
	signal WX4923: std_logic; attribute dont_touch of WX4923: signal is true;
	signal WX4924: std_logic; attribute dont_touch of WX4924: signal is true;
	signal WX4925: std_logic; attribute dont_touch of WX4925: signal is true;
	signal WX4926: std_logic; attribute dont_touch of WX4926: signal is true;
	signal WX4927: std_logic; attribute dont_touch of WX4927: signal is true;
	signal WX4928: std_logic; attribute dont_touch of WX4928: signal is true;
	signal WX4929: std_logic; attribute dont_touch of WX4929: signal is true;
	signal WX4930: std_logic; attribute dont_touch of WX4930: signal is true;
	signal WX4931: std_logic; attribute dont_touch of WX4931: signal is true;
	signal WX4932: std_logic; attribute dont_touch of WX4932: signal is true;
	signal WX4933: std_logic; attribute dont_touch of WX4933: signal is true;
	signal WX4934: std_logic; attribute dont_touch of WX4934: signal is true;
	signal WX4935: std_logic; attribute dont_touch of WX4935: signal is true;
	signal WX4936: std_logic; attribute dont_touch of WX4936: signal is true;
	signal WX4937: std_logic; attribute dont_touch of WX4937: signal is true;
	signal WX4938: std_logic; attribute dont_touch of WX4938: signal is true;
	signal WX4939: std_logic; attribute dont_touch of WX4939: signal is true;
	signal WX4940: std_logic; attribute dont_touch of WX4940: signal is true;
	signal WX4941: std_logic; attribute dont_touch of WX4941: signal is true;
	signal WX4942: std_logic; attribute dont_touch of WX4942: signal is true;
	signal WX4943: std_logic; attribute dont_touch of WX4943: signal is true;
	signal WX4944: std_logic; attribute dont_touch of WX4944: signal is true;
	signal WX4945: std_logic; attribute dont_touch of WX4945: signal is true;
	signal WX4946: std_logic; attribute dont_touch of WX4946: signal is true;
	signal WX4947: std_logic; attribute dont_touch of WX4947: signal is true;
	signal WX4948: std_logic; attribute dont_touch of WX4948: signal is true;
	signal WX4949: std_logic; attribute dont_touch of WX4949: signal is true;
	signal WX4950: std_logic; attribute dont_touch of WX4950: signal is true;
	signal WX4951: std_logic; attribute dont_touch of WX4951: signal is true;
	signal WX4952: std_logic; attribute dont_touch of WX4952: signal is true;
	signal WX4953: std_logic; attribute dont_touch of WX4953: signal is true;
	signal WX4954: std_logic; attribute dont_touch of WX4954: signal is true;
	signal WX4955: std_logic; attribute dont_touch of WX4955: signal is true;
	signal WX4956: std_logic; attribute dont_touch of WX4956: signal is true;
	signal WX4957: std_logic; attribute dont_touch of WX4957: signal is true;
	signal WX4958: std_logic; attribute dont_touch of WX4958: signal is true;
	signal WX4959: std_logic; attribute dont_touch of WX4959: signal is true;
	signal WX4960: std_logic; attribute dont_touch of WX4960: signal is true;
	signal WX4961: std_logic; attribute dont_touch of WX4961: signal is true;
	signal WX4962: std_logic; attribute dont_touch of WX4962: signal is true;
	signal WX4963: std_logic; attribute dont_touch of WX4963: signal is true;
	signal WX4964: std_logic; attribute dont_touch of WX4964: signal is true;
	signal WX4965: std_logic; attribute dont_touch of WX4965: signal is true;
	signal WX4966: std_logic; attribute dont_touch of WX4966: signal is true;
	signal WX4967: std_logic; attribute dont_touch of WX4967: signal is true;
	signal WX4968: std_logic; attribute dont_touch of WX4968: signal is true;
	signal WX4969: std_logic; attribute dont_touch of WX4969: signal is true;
	signal WX4970: std_logic; attribute dont_touch of WX4970: signal is true;
	signal WX4971: std_logic; attribute dont_touch of WX4971: signal is true;
	signal WX4972: std_logic; attribute dont_touch of WX4972: signal is true;
	signal WX4973: std_logic; attribute dont_touch of WX4973: signal is true;
	signal WX4974: std_logic; attribute dont_touch of WX4974: signal is true;
	signal WX4975: std_logic; attribute dont_touch of WX4975: signal is true;
	signal WX4976: std_logic; attribute dont_touch of WX4976: signal is true;
	signal WX4977: std_logic; attribute dont_touch of WX4977: signal is true;
	signal WX4978: std_logic; attribute dont_touch of WX4978: signal is true;
	signal WX4979: std_logic; attribute dont_touch of WX4979: signal is true;
	signal WX4980: std_logic; attribute dont_touch of WX4980: signal is true;
	signal WX4981: std_logic; attribute dont_touch of WX4981: signal is true;
	signal WX4982: std_logic; attribute dont_touch of WX4982: signal is true;
	signal WX4983: std_logic; attribute dont_touch of WX4983: signal is true;
	signal WX4984: std_logic; attribute dont_touch of WX4984: signal is true;
	signal WX4985: std_logic; attribute dont_touch of WX4985: signal is true;
	signal WX4986: std_logic; attribute dont_touch of WX4986: signal is true;
	signal WX4987: std_logic; attribute dont_touch of WX4987: signal is true;
	signal WX4988: std_logic; attribute dont_touch of WX4988: signal is true;
	signal WX4989: std_logic; attribute dont_touch of WX4989: signal is true;
	signal WX4990: std_logic; attribute dont_touch of WX4990: signal is true;
	signal WX4991: std_logic; attribute dont_touch of WX4991: signal is true;
	signal WX4992: std_logic; attribute dont_touch of WX4992: signal is true;
	signal WX4993: std_logic; attribute dont_touch of WX4993: signal is true;
	signal WX4994: std_logic; attribute dont_touch of WX4994: signal is true;
	signal WX4995: std_logic; attribute dont_touch of WX4995: signal is true;
	signal WX4996: std_logic; attribute dont_touch of WX4996: signal is true;
	signal WX4997: std_logic; attribute dont_touch of WX4997: signal is true;
	signal WX4998: std_logic; attribute dont_touch of WX4998: signal is true;
	signal WX4999: std_logic; attribute dont_touch of WX4999: signal is true;
	signal WX5000: std_logic; attribute dont_touch of WX5000: signal is true;
	signal WX5001: std_logic; attribute dont_touch of WX5001: signal is true;
	signal WX5002: std_logic; attribute dont_touch of WX5002: signal is true;
	signal WX5003: std_logic; attribute dont_touch of WX5003: signal is true;
	signal WX5004: std_logic; attribute dont_touch of WX5004: signal is true;
	signal WX5005: std_logic; attribute dont_touch of WX5005: signal is true;
	signal WX5006: std_logic; attribute dont_touch of WX5006: signal is true;
	signal WX5007: std_logic; attribute dont_touch of WX5007: signal is true;
	signal WX5008: std_logic; attribute dont_touch of WX5008: signal is true;
	signal WX5009: std_logic; attribute dont_touch of WX5009: signal is true;
	signal WX5010: std_logic; attribute dont_touch of WX5010: signal is true;
	signal WX5011: std_logic; attribute dont_touch of WX5011: signal is true;
	signal WX5012: std_logic; attribute dont_touch of WX5012: signal is true;
	signal WX5013: std_logic; attribute dont_touch of WX5013: signal is true;
	signal WX5014: std_logic; attribute dont_touch of WX5014: signal is true;
	signal WX5015: std_logic; attribute dont_touch of WX5015: signal is true;
	signal WX5016: std_logic; attribute dont_touch of WX5016: signal is true;
	signal WX5017: std_logic; attribute dont_touch of WX5017: signal is true;
	signal WX5018: std_logic; attribute dont_touch of WX5018: signal is true;
	signal WX5019: std_logic; attribute dont_touch of WX5019: signal is true;
	signal WX5020: std_logic; attribute dont_touch of WX5020: signal is true;
	signal WX5021: std_logic; attribute dont_touch of WX5021: signal is true;
	signal WX5022: std_logic; attribute dont_touch of WX5022: signal is true;
	signal WX5023: std_logic; attribute dont_touch of WX5023: signal is true;
	signal WX5024: std_logic; attribute dont_touch of WX5024: signal is true;
	signal WX5025: std_logic; attribute dont_touch of WX5025: signal is true;
	signal WX5026: std_logic; attribute dont_touch of WX5026: signal is true;
	signal WX5027: std_logic; attribute dont_touch of WX5027: signal is true;
	signal WX5028: std_logic; attribute dont_touch of WX5028: signal is true;
	signal WX5029: std_logic; attribute dont_touch of WX5029: signal is true;
	signal WX5030: std_logic; attribute dont_touch of WX5030: signal is true;
	signal WX5031: std_logic; attribute dont_touch of WX5031: signal is true;
	signal WX5032: std_logic; attribute dont_touch of WX5032: signal is true;
	signal WX5033: std_logic; attribute dont_touch of WX5033: signal is true;
	signal WX5034: std_logic; attribute dont_touch of WX5034: signal is true;
	signal WX5035: std_logic; attribute dont_touch of WX5035: signal is true;
	signal WX5036: std_logic; attribute dont_touch of WX5036: signal is true;
	signal WX5037: std_logic; attribute dont_touch of WX5037: signal is true;
	signal WX5038: std_logic; attribute dont_touch of WX5038: signal is true;
	signal WX5039: std_logic; attribute dont_touch of WX5039: signal is true;
	signal WX5040: std_logic; attribute dont_touch of WX5040: signal is true;
	signal WX5041: std_logic; attribute dont_touch of WX5041: signal is true;
	signal WX5042: std_logic; attribute dont_touch of WX5042: signal is true;
	signal WX5043: std_logic; attribute dont_touch of WX5043: signal is true;
	signal WX5044: std_logic; attribute dont_touch of WX5044: signal is true;
	signal WX5045: std_logic; attribute dont_touch of WX5045: signal is true;
	signal WX5046: std_logic; attribute dont_touch of WX5046: signal is true;
	signal WX5047: std_logic; attribute dont_touch of WX5047: signal is true;
	signal WX5048: std_logic; attribute dont_touch of WX5048: signal is true;
	signal WX5049: std_logic; attribute dont_touch of WX5049: signal is true;
	signal WX5050: std_logic; attribute dont_touch of WX5050: signal is true;
	signal WX5051: std_logic; attribute dont_touch of WX5051: signal is true;
	signal WX5052: std_logic; attribute dont_touch of WX5052: signal is true;
	signal WX5053: std_logic; attribute dont_touch of WX5053: signal is true;
	signal WX5054: std_logic; attribute dont_touch of WX5054: signal is true;
	signal WX5055: std_logic; attribute dont_touch of WX5055: signal is true;
	signal WX5056: std_logic; attribute dont_touch of WX5056: signal is true;
	signal WX5057: std_logic; attribute dont_touch of WX5057: signal is true;
	signal WX5058: std_logic; attribute dont_touch of WX5058: signal is true;
	signal WX5059: std_logic; attribute dont_touch of WX5059: signal is true;
	signal WX5060: std_logic; attribute dont_touch of WX5060: signal is true;
	signal WX5061: std_logic; attribute dont_touch of WX5061: signal is true;
	signal WX5062: std_logic; attribute dont_touch of WX5062: signal is true;
	signal WX5063: std_logic; attribute dont_touch of WX5063: signal is true;
	signal WX5064: std_logic; attribute dont_touch of WX5064: signal is true;
	signal WX5065: std_logic; attribute dont_touch of WX5065: signal is true;
	signal WX5066: std_logic; attribute dont_touch of WX5066: signal is true;
	signal WX5067: std_logic; attribute dont_touch of WX5067: signal is true;
	signal WX5068: std_logic; attribute dont_touch of WX5068: signal is true;
	signal WX5069: std_logic; attribute dont_touch of WX5069: signal is true;
	signal WX5070: std_logic; attribute dont_touch of WX5070: signal is true;
	signal WX5071: std_logic; attribute dont_touch of WX5071: signal is true;
	signal WX5072: std_logic; attribute dont_touch of WX5072: signal is true;
	signal WX5073: std_logic; attribute dont_touch of WX5073: signal is true;
	signal WX5074: std_logic; attribute dont_touch of WX5074: signal is true;
	signal WX5075: std_logic; attribute dont_touch of WX5075: signal is true;
	signal WX5076: std_logic; attribute dont_touch of WX5076: signal is true;
	signal WX5077: std_logic; attribute dont_touch of WX5077: signal is true;
	signal WX5078: std_logic; attribute dont_touch of WX5078: signal is true;
	signal WX5079: std_logic; attribute dont_touch of WX5079: signal is true;
	signal WX5080: std_logic; attribute dont_touch of WX5080: signal is true;
	signal WX5081: std_logic; attribute dont_touch of WX5081: signal is true;
	signal WX5082: std_logic; attribute dont_touch of WX5082: signal is true;
	signal WX5083: std_logic; attribute dont_touch of WX5083: signal is true;
	signal WX5084: std_logic; attribute dont_touch of WX5084: signal is true;
	signal WX5085: std_logic; attribute dont_touch of WX5085: signal is true;
	signal WX5086: std_logic; attribute dont_touch of WX5086: signal is true;
	signal WX5087: std_logic; attribute dont_touch of WX5087: signal is true;
	signal WX5088: std_logic; attribute dont_touch of WX5088: signal is true;
	signal WX5089: std_logic; attribute dont_touch of WX5089: signal is true;
	signal WX5090: std_logic; attribute dont_touch of WX5090: signal is true;
	signal WX5091: std_logic; attribute dont_touch of WX5091: signal is true;
	signal WX5092: std_logic; attribute dont_touch of WX5092: signal is true;
	signal WX5093: std_logic; attribute dont_touch of WX5093: signal is true;
	signal WX5094: std_logic; attribute dont_touch of WX5094: signal is true;
	signal WX5095: std_logic; attribute dont_touch of WX5095: signal is true;
	signal WX5096: std_logic; attribute dont_touch of WX5096: signal is true;
	signal WX5097: std_logic; attribute dont_touch of WX5097: signal is true;
	signal WX5098: std_logic; attribute dont_touch of WX5098: signal is true;
	signal WX5099: std_logic; attribute dont_touch of WX5099: signal is true;
	signal WX5100: std_logic; attribute dont_touch of WX5100: signal is true;
	signal WX5101: std_logic; attribute dont_touch of WX5101: signal is true;
	signal WX5102: std_logic; attribute dont_touch of WX5102: signal is true;
	signal WX5103: std_logic; attribute dont_touch of WX5103: signal is true;
	signal WX5104: std_logic; attribute dont_touch of WX5104: signal is true;
	signal WX5105: std_logic; attribute dont_touch of WX5105: signal is true;
	signal WX5106: std_logic; attribute dont_touch of WX5106: signal is true;
	signal WX5107: std_logic; attribute dont_touch of WX5107: signal is true;
	signal WX5108: std_logic; attribute dont_touch of WX5108: signal is true;
	signal WX5109: std_logic; attribute dont_touch of WX5109: signal is true;
	signal WX5110: std_logic; attribute dont_touch of WX5110: signal is true;
	signal WX5111: std_logic; attribute dont_touch of WX5111: signal is true;
	signal WX5112: std_logic; attribute dont_touch of WX5112: signal is true;
	signal WX5113: std_logic; attribute dont_touch of WX5113: signal is true;
	signal WX5114: std_logic; attribute dont_touch of WX5114: signal is true;
	signal WX5115: std_logic; attribute dont_touch of WX5115: signal is true;
	signal WX5116: std_logic; attribute dont_touch of WX5116: signal is true;
	signal WX5117: std_logic; attribute dont_touch of WX5117: signal is true;
	signal WX5118: std_logic; attribute dont_touch of WX5118: signal is true;
	signal WX5119: std_logic; attribute dont_touch of WX5119: signal is true;
	signal WX5120: std_logic; attribute dont_touch of WX5120: signal is true;
	signal WX5121: std_logic; attribute dont_touch of WX5121: signal is true;
	signal WX5122: std_logic; attribute dont_touch of WX5122: signal is true;
	signal WX5123: std_logic; attribute dont_touch of WX5123: signal is true;
	signal WX5124: std_logic; attribute dont_touch of WX5124: signal is true;
	signal WX5125: std_logic; attribute dont_touch of WX5125: signal is true;
	signal WX5126: std_logic; attribute dont_touch of WX5126: signal is true;
	signal WX5127: std_logic; attribute dont_touch of WX5127: signal is true;
	signal WX5128: std_logic; attribute dont_touch of WX5128: signal is true;
	signal WX5129: std_logic; attribute dont_touch of WX5129: signal is true;
	signal WX5130: std_logic; attribute dont_touch of WX5130: signal is true;
	signal WX5131: std_logic; attribute dont_touch of WX5131: signal is true;
	signal WX5132: std_logic; attribute dont_touch of WX5132: signal is true;
	signal WX5133: std_logic; attribute dont_touch of WX5133: signal is true;
	signal WX5134: std_logic; attribute dont_touch of WX5134: signal is true;
	signal WX5135: std_logic; attribute dont_touch of WX5135: signal is true;
	signal WX5136: std_logic; attribute dont_touch of WX5136: signal is true;
	signal WX5137: std_logic; attribute dont_touch of WX5137: signal is true;
	signal WX5138: std_logic; attribute dont_touch of WX5138: signal is true;
	signal WX5139: std_logic; attribute dont_touch of WX5139: signal is true;
	signal WX5140: std_logic; attribute dont_touch of WX5140: signal is true;
	signal WX5141: std_logic; attribute dont_touch of WX5141: signal is true;
	signal WX5142: std_logic; attribute dont_touch of WX5142: signal is true;
	signal WX5143: std_logic; attribute dont_touch of WX5143: signal is true;
	signal WX5145: std_logic; attribute dont_touch of WX5145: signal is true;
	signal WX5147: std_logic; attribute dont_touch of WX5147: signal is true;
	signal WX5149: std_logic; attribute dont_touch of WX5149: signal is true;
	signal WX5151: std_logic; attribute dont_touch of WX5151: signal is true;
	signal WX5153: std_logic; attribute dont_touch of WX5153: signal is true;
	signal WX5155: std_logic; attribute dont_touch of WX5155: signal is true;
	signal WX5157: std_logic; attribute dont_touch of WX5157: signal is true;
	signal WX5159: std_logic; attribute dont_touch of WX5159: signal is true;
	signal WX5161: std_logic; attribute dont_touch of WX5161: signal is true;
	signal WX5163: std_logic; attribute dont_touch of WX5163: signal is true;
	signal WX5165: std_logic; attribute dont_touch of WX5165: signal is true;
	signal WX5167: std_logic; attribute dont_touch of WX5167: signal is true;
	signal WX5169: std_logic; attribute dont_touch of WX5169: signal is true;
	signal WX5171: std_logic; attribute dont_touch of WX5171: signal is true;
	signal WX5173: std_logic; attribute dont_touch of WX5173: signal is true;
	signal WX5175: std_logic; attribute dont_touch of WX5175: signal is true;
	signal WX5177: std_logic; attribute dont_touch of WX5177: signal is true;
	signal WX5179: std_logic; attribute dont_touch of WX5179: signal is true;
	signal WX5181: std_logic; attribute dont_touch of WX5181: signal is true;
	signal WX5183: std_logic; attribute dont_touch of WX5183: signal is true;
	signal WX5185: std_logic; attribute dont_touch of WX5185: signal is true;
	signal WX5187: std_logic; attribute dont_touch of WX5187: signal is true;
	signal WX5189: std_logic; attribute dont_touch of WX5189: signal is true;
	signal WX5191: std_logic; attribute dont_touch of WX5191: signal is true;
	signal WX5193: std_logic; attribute dont_touch of WX5193: signal is true;
	signal WX5195: std_logic; attribute dont_touch of WX5195: signal is true;
	signal WX5197: std_logic; attribute dont_touch of WX5197: signal is true;
	signal WX5199: std_logic; attribute dont_touch of WX5199: signal is true;
	signal WX5201: std_logic; attribute dont_touch of WX5201: signal is true;
	signal WX5203: std_logic; attribute dont_touch of WX5203: signal is true;
	signal WX5205: std_logic; attribute dont_touch of WX5205: signal is true;
	signal WX5207: std_logic; attribute dont_touch of WX5207: signal is true;
	signal WX5208: std_logic; attribute dont_touch of WX5208: signal is true;
	signal WX5209: std_logic; attribute dont_touch of WX5209: signal is true;
	signal WX5210: std_logic; attribute dont_touch of WX5210: signal is true;
	signal WX5211: std_logic; attribute dont_touch of WX5211: signal is true;
	signal WX5212: std_logic; attribute dont_touch of WX5212: signal is true;
	signal WX5213: std_logic; attribute dont_touch of WX5213: signal is true;
	signal WX5214: std_logic; attribute dont_touch of WX5214: signal is true;
	signal WX5215: std_logic; attribute dont_touch of WX5215: signal is true;
	signal WX5216: std_logic; attribute dont_touch of WX5216: signal is true;
	signal WX5217: std_logic; attribute dont_touch of WX5217: signal is true;
	signal WX5218: std_logic; attribute dont_touch of WX5218: signal is true;
	signal WX5219: std_logic; attribute dont_touch of WX5219: signal is true;
	signal WX5220: std_logic; attribute dont_touch of WX5220: signal is true;
	signal WX5221: std_logic; attribute dont_touch of WX5221: signal is true;
	signal WX5222: std_logic; attribute dont_touch of WX5222: signal is true;
	signal WX5223: std_logic; attribute dont_touch of WX5223: signal is true;
	signal WX5224: std_logic; attribute dont_touch of WX5224: signal is true;
	signal WX5225: std_logic; attribute dont_touch of WX5225: signal is true;
	signal WX5226: std_logic; attribute dont_touch of WX5226: signal is true;
	signal WX5227: std_logic; attribute dont_touch of WX5227: signal is true;
	signal WX5228: std_logic; attribute dont_touch of WX5228: signal is true;
	signal WX5229: std_logic; attribute dont_touch of WX5229: signal is true;
	signal WX5230: std_logic; attribute dont_touch of WX5230: signal is true;
	signal WX5231: std_logic; attribute dont_touch of WX5231: signal is true;
	signal WX5232: std_logic; attribute dont_touch of WX5232: signal is true;
	signal WX5233: std_logic; attribute dont_touch of WX5233: signal is true;
	signal WX5234: std_logic; attribute dont_touch of WX5234: signal is true;
	signal WX5235: std_logic; attribute dont_touch of WX5235: signal is true;
	signal WX5236: std_logic; attribute dont_touch of WX5236: signal is true;
	signal WX5237: std_logic; attribute dont_touch of WX5237: signal is true;
	signal WX5238: std_logic; attribute dont_touch of WX5238: signal is true;
	signal WX5239: std_logic; attribute dont_touch of WX5239: signal is true;
	signal WX5240: std_logic; attribute dont_touch of WX5240: signal is true;
	signal WX5241: std_logic; attribute dont_touch of WX5241: signal is true;
	signal WX5242: std_logic; attribute dont_touch of WX5242: signal is true;
	signal WX5243: std_logic; attribute dont_touch of WX5243: signal is true;
	signal WX5244: std_logic; attribute dont_touch of WX5244: signal is true;
	signal WX5245: std_logic; attribute dont_touch of WX5245: signal is true;
	signal WX5246: std_logic; attribute dont_touch of WX5246: signal is true;
	signal WX5247: std_logic; attribute dont_touch of WX5247: signal is true;
	signal WX5248: std_logic; attribute dont_touch of WX5248: signal is true;
	signal WX5249: std_logic; attribute dont_touch of WX5249: signal is true;
	signal WX5250: std_logic; attribute dont_touch of WX5250: signal is true;
	signal WX5251: std_logic; attribute dont_touch of WX5251: signal is true;
	signal WX5252: std_logic; attribute dont_touch of WX5252: signal is true;
	signal WX5253: std_logic; attribute dont_touch of WX5253: signal is true;
	signal WX5254: std_logic; attribute dont_touch of WX5254: signal is true;
	signal WX5255: std_logic; attribute dont_touch of WX5255: signal is true;
	signal WX5256: std_logic; attribute dont_touch of WX5256: signal is true;
	signal WX5257: std_logic; attribute dont_touch of WX5257: signal is true;
	signal WX5258: std_logic; attribute dont_touch of WX5258: signal is true;
	signal WX5259: std_logic; attribute dont_touch of WX5259: signal is true;
	signal WX5260: std_logic; attribute dont_touch of WX5260: signal is true;
	signal WX5261: std_logic; attribute dont_touch of WX5261: signal is true;
	signal WX5262: std_logic; attribute dont_touch of WX5262: signal is true;
	signal WX5263: std_logic; attribute dont_touch of WX5263: signal is true;
	signal WX5264: std_logic; attribute dont_touch of WX5264: signal is true;
	signal WX5265: std_logic; attribute dont_touch of WX5265: signal is true;
	signal WX5266: std_logic; attribute dont_touch of WX5266: signal is true;
	signal WX5267: std_logic; attribute dont_touch of WX5267: signal is true;
	signal WX5268: std_logic; attribute dont_touch of WX5268: signal is true;
	signal WX5269: std_logic; attribute dont_touch of WX5269: signal is true;
	signal WX5270: std_logic; attribute dont_touch of WX5270: signal is true;
	signal WX5271: std_logic; attribute dont_touch of WX5271: signal is true;
	signal WX5272: std_logic; attribute dont_touch of WX5272: signal is true;
	signal WX5273: std_logic; attribute dont_touch of WX5273: signal is true;
	signal WX5274: std_logic; attribute dont_touch of WX5274: signal is true;
	signal WX5275: std_logic; attribute dont_touch of WX5275: signal is true;
	signal WX5276: std_logic; attribute dont_touch of WX5276: signal is true;
	signal WX5277: std_logic; attribute dont_touch of WX5277: signal is true;
	signal WX5278: std_logic; attribute dont_touch of WX5278: signal is true;
	signal WX5279: std_logic; attribute dont_touch of WX5279: signal is true;
	signal WX5280: std_logic; attribute dont_touch of WX5280: signal is true;
	signal WX5281: std_logic; attribute dont_touch of WX5281: signal is true;
	signal WX5282: std_logic; attribute dont_touch of WX5282: signal is true;
	signal WX5283: std_logic; attribute dont_touch of WX5283: signal is true;
	signal WX5284: std_logic; attribute dont_touch of WX5284: signal is true;
	signal WX5285: std_logic; attribute dont_touch of WX5285: signal is true;
	signal WX5286: std_logic; attribute dont_touch of WX5286: signal is true;
	signal WX5287: std_logic; attribute dont_touch of WX5287: signal is true;
	signal WX5288: std_logic; attribute dont_touch of WX5288: signal is true;
	signal WX5289: std_logic; attribute dont_touch of WX5289: signal is true;
	signal WX5290: std_logic; attribute dont_touch of WX5290: signal is true;
	signal WX5291: std_logic; attribute dont_touch of WX5291: signal is true;
	signal WX5292: std_logic; attribute dont_touch of WX5292: signal is true;
	signal WX5293: std_logic; attribute dont_touch of WX5293: signal is true;
	signal WX5294: std_logic; attribute dont_touch of WX5294: signal is true;
	signal WX5295: std_logic; attribute dont_touch of WX5295: signal is true;
	signal WX5296: std_logic; attribute dont_touch of WX5296: signal is true;
	signal WX5297: std_logic; attribute dont_touch of WX5297: signal is true;
	signal WX5298: std_logic; attribute dont_touch of WX5298: signal is true;
	signal WX5299: std_logic; attribute dont_touch of WX5299: signal is true;
	signal WX5300: std_logic; attribute dont_touch of WX5300: signal is true;
	signal WX5301: std_logic; attribute dont_touch of WX5301: signal is true;
	signal WX5302: std_logic; attribute dont_touch of WX5302: signal is true;
	signal WX5303: std_logic; attribute dont_touch of WX5303: signal is true;
	signal WX5304: std_logic; attribute dont_touch of WX5304: signal is true;
	signal WX5305: std_logic; attribute dont_touch of WX5305: signal is true;
	signal WX5306: std_logic; attribute dont_touch of WX5306: signal is true;
	signal WX5307: std_logic; attribute dont_touch of WX5307: signal is true;
	signal WX5308: std_logic; attribute dont_touch of WX5308: signal is true;
	signal WX5309: std_logic; attribute dont_touch of WX5309: signal is true;
	signal WX5310: std_logic; attribute dont_touch of WX5310: signal is true;
	signal WX5311: std_logic; attribute dont_touch of WX5311: signal is true;
	signal WX5312: std_logic; attribute dont_touch of WX5312: signal is true;
	signal WX5313: std_logic; attribute dont_touch of WX5313: signal is true;
	signal WX5314: std_logic; attribute dont_touch of WX5314: signal is true;
	signal WX5315: std_logic; attribute dont_touch of WX5315: signal is true;
	signal WX5316: std_logic; attribute dont_touch of WX5316: signal is true;
	signal WX5317: std_logic; attribute dont_touch of WX5317: signal is true;
	signal WX5318: std_logic; attribute dont_touch of WX5318: signal is true;
	signal WX5319: std_logic; attribute dont_touch of WX5319: signal is true;
	signal WX5320: std_logic; attribute dont_touch of WX5320: signal is true;
	signal WX5321: std_logic; attribute dont_touch of WX5321: signal is true;
	signal WX5322: std_logic; attribute dont_touch of WX5322: signal is true;
	signal WX5323: std_logic; attribute dont_touch of WX5323: signal is true;
	signal WX5324: std_logic; attribute dont_touch of WX5324: signal is true;
	signal WX5325: std_logic; attribute dont_touch of WX5325: signal is true;
	signal WX5326: std_logic; attribute dont_touch of WX5326: signal is true;
	signal WX5327: std_logic; attribute dont_touch of WX5327: signal is true;
	signal WX5328: std_logic; attribute dont_touch of WX5328: signal is true;
	signal WX5329: std_logic; attribute dont_touch of WX5329: signal is true;
	signal WX5330: std_logic; attribute dont_touch of WX5330: signal is true;
	signal WX5331: std_logic; attribute dont_touch of WX5331: signal is true;
	signal WX5332: std_logic; attribute dont_touch of WX5332: signal is true;
	signal WX5333: std_logic; attribute dont_touch of WX5333: signal is true;
	signal WX5334: std_logic; attribute dont_touch of WX5334: signal is true;
	signal WX5335: std_logic; attribute dont_touch of WX5335: signal is true;
	signal WX5336: std_logic; attribute dont_touch of WX5336: signal is true;
	signal WX5337: std_logic; attribute dont_touch of WX5337: signal is true;
	signal WX5338: std_logic; attribute dont_touch of WX5338: signal is true;
	signal WX5339: std_logic; attribute dont_touch of WX5339: signal is true;
	signal WX5340: std_logic; attribute dont_touch of WX5340: signal is true;
	signal WX5341: std_logic; attribute dont_touch of WX5341: signal is true;
	signal WX5342: std_logic; attribute dont_touch of WX5342: signal is true;
	signal WX5343: std_logic; attribute dont_touch of WX5343: signal is true;
	signal WX5344: std_logic; attribute dont_touch of WX5344: signal is true;
	signal WX5345: std_logic; attribute dont_touch of WX5345: signal is true;
	signal WX5346: std_logic; attribute dont_touch of WX5346: signal is true;
	signal WX5347: std_logic; attribute dont_touch of WX5347: signal is true;
	signal WX5348: std_logic; attribute dont_touch of WX5348: signal is true;
	signal WX5349: std_logic; attribute dont_touch of WX5349: signal is true;
	signal WX5350: std_logic; attribute dont_touch of WX5350: signal is true;
	signal WX5351: std_logic; attribute dont_touch of WX5351: signal is true;
	signal WX5352: std_logic; attribute dont_touch of WX5352: signal is true;
	signal WX5353: std_logic; attribute dont_touch of WX5353: signal is true;
	signal WX5354: std_logic; attribute dont_touch of WX5354: signal is true;
	signal WX5355: std_logic; attribute dont_touch of WX5355: signal is true;
	signal WX5356: std_logic; attribute dont_touch of WX5356: signal is true;
	signal WX5357: std_logic; attribute dont_touch of WX5357: signal is true;
	signal WX5358: std_logic; attribute dont_touch of WX5358: signal is true;
	signal WX5359: std_logic; attribute dont_touch of WX5359: signal is true;
	signal WX5360: std_logic; attribute dont_touch of WX5360: signal is true;
	signal WX5361: std_logic; attribute dont_touch of WX5361: signal is true;
	signal WX5362: std_logic; attribute dont_touch of WX5362: signal is true;
	signal WX5363: std_logic; attribute dont_touch of WX5363: signal is true;
	signal WX5364: std_logic; attribute dont_touch of WX5364: signal is true;
	signal WX5365: std_logic; attribute dont_touch of WX5365: signal is true;
	signal WX5366: std_logic; attribute dont_touch of WX5366: signal is true;
	signal WX5367: std_logic; attribute dont_touch of WX5367: signal is true;
	signal WX5368: std_logic; attribute dont_touch of WX5368: signal is true;
	signal WX5369: std_logic; attribute dont_touch of WX5369: signal is true;
	signal WX5370: std_logic; attribute dont_touch of WX5370: signal is true;
	signal WX5371: std_logic; attribute dont_touch of WX5371: signal is true;
	signal WX5372: std_logic; attribute dont_touch of WX5372: signal is true;
	signal WX5373: std_logic; attribute dont_touch of WX5373: signal is true;
	signal WX5374: std_logic; attribute dont_touch of WX5374: signal is true;
	signal WX5375: std_logic; attribute dont_touch of WX5375: signal is true;
	signal WX5376: std_logic; attribute dont_touch of WX5376: signal is true;
	signal WX5377: std_logic; attribute dont_touch of WX5377: signal is true;
	signal WX5378: std_logic; attribute dont_touch of WX5378: signal is true;
	signal WX5379: std_logic; attribute dont_touch of WX5379: signal is true;
	signal WX5380: std_logic; attribute dont_touch of WX5380: signal is true;
	signal WX5381: std_logic; attribute dont_touch of WX5381: signal is true;
	signal WX5382: std_logic; attribute dont_touch of WX5382: signal is true;
	signal WX5383: std_logic; attribute dont_touch of WX5383: signal is true;
	signal WX5384: std_logic; attribute dont_touch of WX5384: signal is true;
	signal WX5385: std_logic; attribute dont_touch of WX5385: signal is true;
	signal WX5386: std_logic; attribute dont_touch of WX5386: signal is true;
	signal WX5387: std_logic; attribute dont_touch of WX5387: signal is true;
	signal WX5388: std_logic; attribute dont_touch of WX5388: signal is true;
	signal WX5389: std_logic; attribute dont_touch of WX5389: signal is true;
	signal WX5390: std_logic; attribute dont_touch of WX5390: signal is true;
	signal WX5391: std_logic; attribute dont_touch of WX5391: signal is true;
	signal WX5392: std_logic; attribute dont_touch of WX5392: signal is true;
	signal WX5393: std_logic; attribute dont_touch of WX5393: signal is true;
	signal WX5394: std_logic; attribute dont_touch of WX5394: signal is true;
	signal WX5395: std_logic; attribute dont_touch of WX5395: signal is true;
	signal WX5396: std_logic; attribute dont_touch of WX5396: signal is true;
	signal WX5397: std_logic; attribute dont_touch of WX5397: signal is true;
	signal WX5398: std_logic; attribute dont_touch of WX5398: signal is true;
	signal WX5399: std_logic; attribute dont_touch of WX5399: signal is true;
	signal WX5400: std_logic; attribute dont_touch of WX5400: signal is true;
	signal WX5401: std_logic; attribute dont_touch of WX5401: signal is true;
	signal WX5402: std_logic; attribute dont_touch of WX5402: signal is true;
	signal WX5403: std_logic; attribute dont_touch of WX5403: signal is true;
	signal WX5404: std_logic; attribute dont_touch of WX5404: signal is true;
	signal WX5405: std_logic; attribute dont_touch of WX5405: signal is true;
	signal WX5406: std_logic; attribute dont_touch of WX5406: signal is true;
	signal WX5407: std_logic; attribute dont_touch of WX5407: signal is true;
	signal WX5408: std_logic; attribute dont_touch of WX5408: signal is true;
	signal WX5409: std_logic; attribute dont_touch of WX5409: signal is true;
	signal WX5410: std_logic; attribute dont_touch of WX5410: signal is true;
	signal WX5411: std_logic; attribute dont_touch of WX5411: signal is true;
	signal WX5412: std_logic; attribute dont_touch of WX5412: signal is true;
	signal WX5413: std_logic; attribute dont_touch of WX5413: signal is true;
	signal WX5414: std_logic; attribute dont_touch of WX5414: signal is true;
	signal WX5415: std_logic; attribute dont_touch of WX5415: signal is true;
	signal WX5416: std_logic; attribute dont_touch of WX5416: signal is true;
	signal WX5417: std_logic; attribute dont_touch of WX5417: signal is true;
	signal WX5418: std_logic; attribute dont_touch of WX5418: signal is true;
	signal WX5419: std_logic; attribute dont_touch of WX5419: signal is true;
	signal WX5420: std_logic; attribute dont_touch of WX5420: signal is true;
	signal WX5421: std_logic; attribute dont_touch of WX5421: signal is true;
	signal WX5422: std_logic; attribute dont_touch of WX5422: signal is true;
	signal WX5423: std_logic; attribute dont_touch of WX5423: signal is true;
	signal WX5424: std_logic; attribute dont_touch of WX5424: signal is true;
	signal WX5425: std_logic; attribute dont_touch of WX5425: signal is true;
	signal WX5426: std_logic; attribute dont_touch of WX5426: signal is true;
	signal WX5427: std_logic; attribute dont_touch of WX5427: signal is true;
	signal WX5428: std_logic; attribute dont_touch of WX5428: signal is true;
	signal WX5429: std_logic; attribute dont_touch of WX5429: signal is true;
	signal WX5430: std_logic; attribute dont_touch of WX5430: signal is true;
	signal WX5431: std_logic; attribute dont_touch of WX5431: signal is true;
	signal WX5432: std_logic; attribute dont_touch of WX5432: signal is true;
	signal WX5433: std_logic; attribute dont_touch of WX5433: signal is true;
	signal WX5434: std_logic; attribute dont_touch of WX5434: signal is true;
	signal WX5435: std_logic; attribute dont_touch of WX5435: signal is true;
	signal WX5436: std_logic; attribute dont_touch of WX5436: signal is true;
	signal WX5437: std_logic; attribute dont_touch of WX5437: signal is true;
	signal WX5438: std_logic; attribute dont_touch of WX5438: signal is true;
	signal WX5439: std_logic; attribute dont_touch of WX5439: signal is true;
	signal WX5440: std_logic; attribute dont_touch of WX5440: signal is true;
	signal WX5441: std_logic; attribute dont_touch of WX5441: signal is true;
	signal WX5442: std_logic; attribute dont_touch of WX5442: signal is true;
	signal WX5443: std_logic; attribute dont_touch of WX5443: signal is true;
	signal WX5444: std_logic; attribute dont_touch of WX5444: signal is true;
	signal WX5445: std_logic; attribute dont_touch of WX5445: signal is true;
	signal WX5446: std_logic; attribute dont_touch of WX5446: signal is true;
	signal WX5447: std_logic; attribute dont_touch of WX5447: signal is true;
	signal WX5448: std_logic; attribute dont_touch of WX5448: signal is true;
	signal WX5449: std_logic; attribute dont_touch of WX5449: signal is true;
	signal WX5450: std_logic; attribute dont_touch of WX5450: signal is true;
	signal WX5451: std_logic; attribute dont_touch of WX5451: signal is true;
	signal WX5452: std_logic; attribute dont_touch of WX5452: signal is true;
	signal WX5453: std_logic; attribute dont_touch of WX5453: signal is true;
	signal WX5454: std_logic; attribute dont_touch of WX5454: signal is true;
	signal WX5455: std_logic; attribute dont_touch of WX5455: signal is true;
	signal WX5456: std_logic; attribute dont_touch of WX5456: signal is true;
	signal WX5457: std_logic; attribute dont_touch of WX5457: signal is true;
	signal WX5458: std_logic; attribute dont_touch of WX5458: signal is true;
	signal WX5459: std_logic; attribute dont_touch of WX5459: signal is true;
	signal WX5460: std_logic; attribute dont_touch of WX5460: signal is true;
	signal WX5461: std_logic; attribute dont_touch of WX5461: signal is true;
	signal WX5462: std_logic; attribute dont_touch of WX5462: signal is true;
	signal WX5463: std_logic; attribute dont_touch of WX5463: signal is true;
	signal WX5464: std_logic; attribute dont_touch of WX5464: signal is true;
	signal WX5465: std_logic; attribute dont_touch of WX5465: signal is true;
	signal WX5466: std_logic; attribute dont_touch of WX5466: signal is true;
	signal WX5467: std_logic; attribute dont_touch of WX5467: signal is true;
	signal WX5468: std_logic; attribute dont_touch of WX5468: signal is true;
	signal WX5469: std_logic; attribute dont_touch of WX5469: signal is true;
	signal WX5470: std_logic; attribute dont_touch of WX5470: signal is true;
	signal WX5471: std_logic; attribute dont_touch of WX5471: signal is true;
	signal WX5472: std_logic; attribute dont_touch of WX5472: signal is true;
	signal WX5473: std_logic; attribute dont_touch of WX5473: signal is true;
	signal WX5474: std_logic; attribute dont_touch of WX5474: signal is true;
	signal WX5475: std_logic; attribute dont_touch of WX5475: signal is true;
	signal WX5476: std_logic; attribute dont_touch of WX5476: signal is true;
	signal WX5477: std_logic; attribute dont_touch of WX5477: signal is true;
	signal WX5478: std_logic; attribute dont_touch of WX5478: signal is true;
	signal WX5479: std_logic; attribute dont_touch of WX5479: signal is true;
	signal WX5480: std_logic; attribute dont_touch of WX5480: signal is true;
	signal WX5481: std_logic; attribute dont_touch of WX5481: signal is true;
	signal WX5482: std_logic; attribute dont_touch of WX5482: signal is true;
	signal WX5483: std_logic; attribute dont_touch of WX5483: signal is true;
	signal WX5484: std_logic; attribute dont_touch of WX5484: signal is true;
	signal WX5485: std_logic; attribute dont_touch of WX5485: signal is true;
	signal WX5486: std_logic; attribute dont_touch of WX5486: signal is true;
	signal WX5487: std_logic; attribute dont_touch of WX5487: signal is true;
	signal WX5488: std_logic; attribute dont_touch of WX5488: signal is true;
	signal WX5489: std_logic; attribute dont_touch of WX5489: signal is true;
	signal WX5490: std_logic; attribute dont_touch of WX5490: signal is true;
	signal WX5491: std_logic; attribute dont_touch of WX5491: signal is true;
	signal WX5492: std_logic; attribute dont_touch of WX5492: signal is true;
	signal WX5493: std_logic; attribute dont_touch of WX5493: signal is true;
	signal WX5494: std_logic; attribute dont_touch of WX5494: signal is true;
	signal WX5495: std_logic; attribute dont_touch of WX5495: signal is true;
	signal WX5496: std_logic; attribute dont_touch of WX5496: signal is true;
	signal WX5497: std_logic; attribute dont_touch of WX5497: signal is true;
	signal WX5498: std_logic; attribute dont_touch of WX5498: signal is true;
	signal WX5499: std_logic; attribute dont_touch of WX5499: signal is true;
	signal WX5500: std_logic; attribute dont_touch of WX5500: signal is true;
	signal WX5501: std_logic; attribute dont_touch of WX5501: signal is true;
	signal WX5502: std_logic; attribute dont_touch of WX5502: signal is true;
	signal WX5503: std_logic; attribute dont_touch of WX5503: signal is true;
	signal WX5504: std_logic; attribute dont_touch of WX5504: signal is true;
	signal WX5505: std_logic; attribute dont_touch of WX5505: signal is true;
	signal WX5506: std_logic; attribute dont_touch of WX5506: signal is true;
	signal WX5507: std_logic; attribute dont_touch of WX5507: signal is true;
	signal WX5508: std_logic; attribute dont_touch of WX5508: signal is true;
	signal WX5509: std_logic; attribute dont_touch of WX5509: signal is true;
	signal WX5510: std_logic; attribute dont_touch of WX5510: signal is true;
	signal WX5511: std_logic; attribute dont_touch of WX5511: signal is true;
	signal WX5512: std_logic; attribute dont_touch of WX5512: signal is true;
	signal WX5513: std_logic; attribute dont_touch of WX5513: signal is true;
	signal WX5514: std_logic; attribute dont_touch of WX5514: signal is true;
	signal WX5515: std_logic; attribute dont_touch of WX5515: signal is true;
	signal WX5516: std_logic; attribute dont_touch of WX5516: signal is true;
	signal WX5517: std_logic; attribute dont_touch of WX5517: signal is true;
	signal WX5518: std_logic; attribute dont_touch of WX5518: signal is true;
	signal WX5519: std_logic; attribute dont_touch of WX5519: signal is true;
	signal WX5520: std_logic; attribute dont_touch of WX5520: signal is true;
	signal WX5521: std_logic; attribute dont_touch of WX5521: signal is true;
	signal WX5522: std_logic; attribute dont_touch of WX5522: signal is true;
	signal WX5523: std_logic; attribute dont_touch of WX5523: signal is true;
	signal WX5524: std_logic; attribute dont_touch of WX5524: signal is true;
	signal WX5525: std_logic; attribute dont_touch of WX5525: signal is true;
	signal WX5526: std_logic; attribute dont_touch of WX5526: signal is true;
	signal WX5527: std_logic; attribute dont_touch of WX5527: signal is true;
	signal WX5528: std_logic; attribute dont_touch of WX5528: signal is true;
	signal WX5529: std_logic; attribute dont_touch of WX5529: signal is true;
	signal WX5530: std_logic; attribute dont_touch of WX5530: signal is true;
	signal WX5531: std_logic; attribute dont_touch of WX5531: signal is true;
	signal WX5532: std_logic; attribute dont_touch of WX5532: signal is true;
	signal WX5533: std_logic; attribute dont_touch of WX5533: signal is true;
	signal WX5534: std_logic; attribute dont_touch of WX5534: signal is true;
	signal WX5535: std_logic; attribute dont_touch of WX5535: signal is true;
	signal WX5536: std_logic; attribute dont_touch of WX5536: signal is true;
	signal WX5537: std_logic; attribute dont_touch of WX5537: signal is true;
	signal WX5538: std_logic; attribute dont_touch of WX5538: signal is true;
	signal WX5539: std_logic; attribute dont_touch of WX5539: signal is true;
	signal WX5540: std_logic; attribute dont_touch of WX5540: signal is true;
	signal WX5541: std_logic; attribute dont_touch of WX5541: signal is true;
	signal WX5542: std_logic; attribute dont_touch of WX5542: signal is true;
	signal WX5543: std_logic; attribute dont_touch of WX5543: signal is true;
	signal WX5544: std_logic; attribute dont_touch of WX5544: signal is true;
	signal WX5545: std_logic; attribute dont_touch of WX5545: signal is true;
	signal WX5546: std_logic; attribute dont_touch of WX5546: signal is true;
	signal WX5547: std_logic; attribute dont_touch of WX5547: signal is true;
	signal WX5548: std_logic; attribute dont_touch of WX5548: signal is true;
	signal WX5549: std_logic; attribute dont_touch of WX5549: signal is true;
	signal WX5550: std_logic; attribute dont_touch of WX5550: signal is true;
	signal WX5551: std_logic; attribute dont_touch of WX5551: signal is true;
	signal WX5552: std_logic; attribute dont_touch of WX5552: signal is true;
	signal WX5553: std_logic; attribute dont_touch of WX5553: signal is true;
	signal WX5554: std_logic; attribute dont_touch of WX5554: signal is true;
	signal WX5555: std_logic; attribute dont_touch of WX5555: signal is true;
	signal WX5556: std_logic; attribute dont_touch of WX5556: signal is true;
	signal WX5557: std_logic; attribute dont_touch of WX5557: signal is true;
	signal WX5558: std_logic; attribute dont_touch of WX5558: signal is true;
	signal WX5559: std_logic; attribute dont_touch of WX5559: signal is true;
	signal WX5560: std_logic; attribute dont_touch of WX5560: signal is true;
	signal WX5561: std_logic; attribute dont_touch of WX5561: signal is true;
	signal WX5562: std_logic; attribute dont_touch of WX5562: signal is true;
	signal WX5563: std_logic; attribute dont_touch of WX5563: signal is true;
	signal WX5564: std_logic; attribute dont_touch of WX5564: signal is true;
	signal WX5565: std_logic; attribute dont_touch of WX5565: signal is true;
	signal WX5566: std_logic; attribute dont_touch of WX5566: signal is true;
	signal WX5567: std_logic; attribute dont_touch of WX5567: signal is true;
	signal WX5568: std_logic; attribute dont_touch of WX5568: signal is true;
	signal WX5569: std_logic; attribute dont_touch of WX5569: signal is true;
	signal WX5570: std_logic; attribute dont_touch of WX5570: signal is true;
	signal WX5571: std_logic; attribute dont_touch of WX5571: signal is true;
	signal WX5572: std_logic; attribute dont_touch of WX5572: signal is true;
	signal WX5573: std_logic; attribute dont_touch of WX5573: signal is true;
	signal WX5574: std_logic; attribute dont_touch of WX5574: signal is true;
	signal WX5575: std_logic; attribute dont_touch of WX5575: signal is true;
	signal WX5576: std_logic; attribute dont_touch of WX5576: signal is true;
	signal WX5577: std_logic; attribute dont_touch of WX5577: signal is true;
	signal WX5578: std_logic; attribute dont_touch of WX5578: signal is true;
	signal WX5579: std_logic; attribute dont_touch of WX5579: signal is true;
	signal WX5580: std_logic; attribute dont_touch of WX5580: signal is true;
	signal WX5581: std_logic; attribute dont_touch of WX5581: signal is true;
	signal WX5582: std_logic; attribute dont_touch of WX5582: signal is true;
	signal WX5583: std_logic; attribute dont_touch of WX5583: signal is true;
	signal WX5584: std_logic; attribute dont_touch of WX5584: signal is true;
	signal WX5585: std_logic; attribute dont_touch of WX5585: signal is true;
	signal WX5586: std_logic; attribute dont_touch of WX5586: signal is true;
	signal WX5587: std_logic; attribute dont_touch of WX5587: signal is true;
	signal WX5588: std_logic; attribute dont_touch of WX5588: signal is true;
	signal WX5589: std_logic; attribute dont_touch of WX5589: signal is true;
	signal WX5590: std_logic; attribute dont_touch of WX5590: signal is true;
	signal WX5591: std_logic; attribute dont_touch of WX5591: signal is true;
	signal WX5592: std_logic; attribute dont_touch of WX5592: signal is true;
	signal WX5593: std_logic; attribute dont_touch of WX5593: signal is true;
	signal WX5594: std_logic; attribute dont_touch of WX5594: signal is true;
	signal WX5595: std_logic; attribute dont_touch of WX5595: signal is true;
	signal WX5596: std_logic; attribute dont_touch of WX5596: signal is true;
	signal WX5597: std_logic; attribute dont_touch of WX5597: signal is true;
	signal WX5598: std_logic; attribute dont_touch of WX5598: signal is true;
	signal WX5599: std_logic; attribute dont_touch of WX5599: signal is true;
	signal WX5600: std_logic; attribute dont_touch of WX5600: signal is true;
	signal WX5601: std_logic; attribute dont_touch of WX5601: signal is true;
	signal WX5602: std_logic; attribute dont_touch of WX5602: signal is true;
	signal WX5603: std_logic; attribute dont_touch of WX5603: signal is true;
	signal WX5604: std_logic; attribute dont_touch of WX5604: signal is true;
	signal WX5605: std_logic; attribute dont_touch of WX5605: signal is true;
	signal WX5606: std_logic; attribute dont_touch of WX5606: signal is true;
	signal WX5607: std_logic; attribute dont_touch of WX5607: signal is true;
	signal WX5608: std_logic; attribute dont_touch of WX5608: signal is true;
	signal WX5609: std_logic; attribute dont_touch of WX5609: signal is true;
	signal WX5610: std_logic; attribute dont_touch of WX5610: signal is true;
	signal WX5611: std_logic; attribute dont_touch of WX5611: signal is true;
	signal WX5612: std_logic; attribute dont_touch of WX5612: signal is true;
	signal WX5613: std_logic; attribute dont_touch of WX5613: signal is true;
	signal WX5614: std_logic; attribute dont_touch of WX5614: signal is true;
	signal WX5615: std_logic; attribute dont_touch of WX5615: signal is true;
	signal WX5616: std_logic; attribute dont_touch of WX5616: signal is true;
	signal WX5617: std_logic; attribute dont_touch of WX5617: signal is true;
	signal WX5618: std_logic; attribute dont_touch of WX5618: signal is true;
	signal WX5619: std_logic; attribute dont_touch of WX5619: signal is true;
	signal WX5620: std_logic; attribute dont_touch of WX5620: signal is true;
	signal WX5621: std_logic; attribute dont_touch of WX5621: signal is true;
	signal WX5622: std_logic; attribute dont_touch of WX5622: signal is true;
	signal WX5623: std_logic; attribute dont_touch of WX5623: signal is true;
	signal WX5624: std_logic; attribute dont_touch of WX5624: signal is true;
	signal WX5625: std_logic; attribute dont_touch of WX5625: signal is true;
	signal WX5626: std_logic; attribute dont_touch of WX5626: signal is true;
	signal WX5627: std_logic; attribute dont_touch of WX5627: signal is true;
	signal WX5628: std_logic; attribute dont_touch of WX5628: signal is true;
	signal WX5629: std_logic; attribute dont_touch of WX5629: signal is true;
	signal WX5630: std_logic; attribute dont_touch of WX5630: signal is true;
	signal WX5631: std_logic; attribute dont_touch of WX5631: signal is true;
	signal WX5632: std_logic; attribute dont_touch of WX5632: signal is true;
	signal WX5633: std_logic; attribute dont_touch of WX5633: signal is true;
	signal WX5634: std_logic; attribute dont_touch of WX5634: signal is true;
	signal WX5635: std_logic; attribute dont_touch of WX5635: signal is true;
	signal WX5636: std_logic; attribute dont_touch of WX5636: signal is true;
	signal WX5637: std_logic; attribute dont_touch of WX5637: signal is true;
	signal WX5638: std_logic; attribute dont_touch of WX5638: signal is true;
	signal WX5639: std_logic; attribute dont_touch of WX5639: signal is true;
	signal WX5640: std_logic; attribute dont_touch of WX5640: signal is true;
	signal WX5641: std_logic; attribute dont_touch of WX5641: signal is true;
	signal WX5642: std_logic; attribute dont_touch of WX5642: signal is true;
	signal WX5643: std_logic; attribute dont_touch of WX5643: signal is true;
	signal WX5644: std_logic; attribute dont_touch of WX5644: signal is true;
	signal WX5645: std_logic; attribute dont_touch of WX5645: signal is true;
	signal WX5646: std_logic; attribute dont_touch of WX5646: signal is true;
	signal WX5647: std_logic; attribute dont_touch of WX5647: signal is true;
	signal WX5648: std_logic; attribute dont_touch of WX5648: signal is true;
	signal WX5649: std_logic; attribute dont_touch of WX5649: signal is true;
	signal WX5650: std_logic; attribute dont_touch of WX5650: signal is true;
	signal WX5651: std_logic; attribute dont_touch of WX5651: signal is true;
	signal WX5652: std_logic; attribute dont_touch of WX5652: signal is true;
	signal WX5653: std_logic; attribute dont_touch of WX5653: signal is true;
	signal WX5654: std_logic; attribute dont_touch of WX5654: signal is true;
	signal WX5655: std_logic; attribute dont_touch of WX5655: signal is true;
	signal WX5656: std_logic; attribute dont_touch of WX5656: signal is true;
	signal WX5657: std_logic; attribute dont_touch of WX5657: signal is true;
	signal WX5658: std_logic; attribute dont_touch of WX5658: signal is true;
	signal WX5659: std_logic; attribute dont_touch of WX5659: signal is true;
	signal WX5660: std_logic; attribute dont_touch of WX5660: signal is true;
	signal WX5661: std_logic; attribute dont_touch of WX5661: signal is true;
	signal WX5662: std_logic; attribute dont_touch of WX5662: signal is true;
	signal WX5663: std_logic; attribute dont_touch of WX5663: signal is true;
	signal WX5664: std_logic; attribute dont_touch of WX5664: signal is true;
	signal WX5665: std_logic; attribute dont_touch of WX5665: signal is true;
	signal WX5666: std_logic; attribute dont_touch of WX5666: signal is true;
	signal WX5667: std_logic; attribute dont_touch of WX5667: signal is true;
	signal WX5668: std_logic; attribute dont_touch of WX5668: signal is true;
	signal WX5669: std_logic; attribute dont_touch of WX5669: signal is true;
	signal WX5670: std_logic; attribute dont_touch of WX5670: signal is true;
	signal WX5671: std_logic; attribute dont_touch of WX5671: signal is true;
	signal WX5672: std_logic; attribute dont_touch of WX5672: signal is true;
	signal WX5673: std_logic; attribute dont_touch of WX5673: signal is true;
	signal WX5674: std_logic; attribute dont_touch of WX5674: signal is true;
	signal WX5675: std_logic; attribute dont_touch of WX5675: signal is true;
	signal WX5676: std_logic; attribute dont_touch of WX5676: signal is true;
	signal WX5677: std_logic; attribute dont_touch of WX5677: signal is true;
	signal WX5678: std_logic; attribute dont_touch of WX5678: signal is true;
	signal WX5679: std_logic; attribute dont_touch of WX5679: signal is true;
	signal WX5680: std_logic; attribute dont_touch of WX5680: signal is true;
	signal WX5681: std_logic; attribute dont_touch of WX5681: signal is true;
	signal WX5682: std_logic; attribute dont_touch of WX5682: signal is true;
	signal WX5683: std_logic; attribute dont_touch of WX5683: signal is true;
	signal WX5684: std_logic; attribute dont_touch of WX5684: signal is true;
	signal WX5685: std_logic; attribute dont_touch of WX5685: signal is true;
	signal WX5686: std_logic; attribute dont_touch of WX5686: signal is true;
	signal WX5687: std_logic; attribute dont_touch of WX5687: signal is true;
	signal WX5688: std_logic; attribute dont_touch of WX5688: signal is true;
	signal WX5689: std_logic; attribute dont_touch of WX5689: signal is true;
	signal WX5690: std_logic; attribute dont_touch of WX5690: signal is true;
	signal WX5691: std_logic; attribute dont_touch of WX5691: signal is true;
	signal WX5692: std_logic; attribute dont_touch of WX5692: signal is true;
	signal WX5693: std_logic; attribute dont_touch of WX5693: signal is true;
	signal WX5694: std_logic; attribute dont_touch of WX5694: signal is true;
	signal WX5695: std_logic; attribute dont_touch of WX5695: signal is true;
	signal WX5696: std_logic; attribute dont_touch of WX5696: signal is true;
	signal WX5697: std_logic; attribute dont_touch of WX5697: signal is true;
	signal WX5698: std_logic; attribute dont_touch of WX5698: signal is true;
	signal WX5699: std_logic; attribute dont_touch of WX5699: signal is true;
	signal WX5700: std_logic; attribute dont_touch of WX5700: signal is true;
	signal WX5701: std_logic; attribute dont_touch of WX5701: signal is true;
	signal WX5702: std_logic; attribute dont_touch of WX5702: signal is true;
	signal WX5703: std_logic; attribute dont_touch of WX5703: signal is true;
	signal WX5704: std_logic; attribute dont_touch of WX5704: signal is true;
	signal WX5705: std_logic; attribute dont_touch of WX5705: signal is true;
	signal WX5706: std_logic; attribute dont_touch of WX5706: signal is true;
	signal WX5707: std_logic; attribute dont_touch of WX5707: signal is true;
	signal WX5708: std_logic; attribute dont_touch of WX5708: signal is true;
	signal WX5709: std_logic; attribute dont_touch of WX5709: signal is true;
	signal WX5710: std_logic; attribute dont_touch of WX5710: signal is true;
	signal WX5711: std_logic; attribute dont_touch of WX5711: signal is true;
	signal WX5712: std_logic; attribute dont_touch of WX5712: signal is true;
	signal WX5713: std_logic; attribute dont_touch of WX5713: signal is true;
	signal WX5714: std_logic; attribute dont_touch of WX5714: signal is true;
	signal WX5715: std_logic; attribute dont_touch of WX5715: signal is true;
	signal WX5716: std_logic; attribute dont_touch of WX5716: signal is true;
	signal WX5717: std_logic; attribute dont_touch of WX5717: signal is true;
	signal WX5718: std_logic; attribute dont_touch of WX5718: signal is true;
	signal WX5719: std_logic; attribute dont_touch of WX5719: signal is true;
	signal WX5720: std_logic; attribute dont_touch of WX5720: signal is true;
	signal WX5721: std_logic; attribute dont_touch of WX5721: signal is true;
	signal WX5722: std_logic; attribute dont_touch of WX5722: signal is true;
	signal WX5723: std_logic; attribute dont_touch of WX5723: signal is true;
	signal WX5724: std_logic; attribute dont_touch of WX5724: signal is true;
	signal WX5725: std_logic; attribute dont_touch of WX5725: signal is true;
	signal WX5726: std_logic; attribute dont_touch of WX5726: signal is true;
	signal WX5727: std_logic; attribute dont_touch of WX5727: signal is true;
	signal WX5728: std_logic; attribute dont_touch of WX5728: signal is true;
	signal WX5729: std_logic; attribute dont_touch of WX5729: signal is true;
	signal WX5730: std_logic; attribute dont_touch of WX5730: signal is true;
	signal WX5731: std_logic; attribute dont_touch of WX5731: signal is true;
	signal WX5732: std_logic; attribute dont_touch of WX5732: signal is true;
	signal WX5733: std_logic; attribute dont_touch of WX5733: signal is true;
	signal WX5734: std_logic; attribute dont_touch of WX5734: signal is true;
	signal WX5735: std_logic; attribute dont_touch of WX5735: signal is true;
	signal WX5736: std_logic; attribute dont_touch of WX5736: signal is true;
	signal WX5737: std_logic; attribute dont_touch of WX5737: signal is true;
	signal WX5738: std_logic; attribute dont_touch of WX5738: signal is true;
	signal WX5739: std_logic; attribute dont_touch of WX5739: signal is true;
	signal WX5740: std_logic; attribute dont_touch of WX5740: signal is true;
	signal WX5741: std_logic; attribute dont_touch of WX5741: signal is true;
	signal WX5742: std_logic; attribute dont_touch of WX5742: signal is true;
	signal WX5743: std_logic; attribute dont_touch of WX5743: signal is true;
	signal WX5744: std_logic; attribute dont_touch of WX5744: signal is true;
	signal WX5745: std_logic; attribute dont_touch of WX5745: signal is true;
	signal WX5746: std_logic; attribute dont_touch of WX5746: signal is true;
	signal WX5747: std_logic; attribute dont_touch of WX5747: signal is true;
	signal WX5748: std_logic; attribute dont_touch of WX5748: signal is true;
	signal WX5749: std_logic; attribute dont_touch of WX5749: signal is true;
	signal WX5750: std_logic; attribute dont_touch of WX5750: signal is true;
	signal WX5751: std_logic; attribute dont_touch of WX5751: signal is true;
	signal WX5752: std_logic; attribute dont_touch of WX5752: signal is true;
	signal WX5753: std_logic; attribute dont_touch of WX5753: signal is true;
	signal WX5754: std_logic; attribute dont_touch of WX5754: signal is true;
	signal WX5755: std_logic; attribute dont_touch of WX5755: signal is true;
	signal WX5756: std_logic; attribute dont_touch of WX5756: signal is true;
	signal WX5757: std_logic; attribute dont_touch of WX5757: signal is true;
	signal WX5758: std_logic; attribute dont_touch of WX5758: signal is true;
	signal WX5759: std_logic; attribute dont_touch of WX5759: signal is true;
	signal WX5760: std_logic; attribute dont_touch of WX5760: signal is true;
	signal WX5761: std_logic; attribute dont_touch of WX5761: signal is true;
	signal WX5762: std_logic; attribute dont_touch of WX5762: signal is true;
	signal WX5763: std_logic; attribute dont_touch of WX5763: signal is true;
	signal WX5764: std_logic; attribute dont_touch of WX5764: signal is true;
	signal WX5765: std_logic; attribute dont_touch of WX5765: signal is true;
	signal WX5766: std_logic; attribute dont_touch of WX5766: signal is true;
	signal WX5767: std_logic; attribute dont_touch of WX5767: signal is true;
	signal WX5768: std_logic; attribute dont_touch of WX5768: signal is true;
	signal WX5769: std_logic; attribute dont_touch of WX5769: signal is true;
	signal WX5770: std_logic; attribute dont_touch of WX5770: signal is true;
	signal WX5771: std_logic; attribute dont_touch of WX5771: signal is true;
	signal WX5772: std_logic; attribute dont_touch of WX5772: signal is true;
	signal WX5773: std_logic; attribute dont_touch of WX5773: signal is true;
	signal WX5774: std_logic; attribute dont_touch of WX5774: signal is true;
	signal WX5775: std_logic; attribute dont_touch of WX5775: signal is true;
	signal WX5776: std_logic; attribute dont_touch of WX5776: signal is true;
	signal WX5777: std_logic; attribute dont_touch of WX5777: signal is true;
	signal WX5778: std_logic; attribute dont_touch of WX5778: signal is true;
	signal WX5779: std_logic; attribute dont_touch of WX5779: signal is true;
	signal WX5780: std_logic; attribute dont_touch of WX5780: signal is true;
	signal WX5781: std_logic; attribute dont_touch of WX5781: signal is true;
	signal WX5782: std_logic; attribute dont_touch of WX5782: signal is true;
	signal WX5783: std_logic; attribute dont_touch of WX5783: signal is true;
	signal WX5784: std_logic; attribute dont_touch of WX5784: signal is true;
	signal WX5785: std_logic; attribute dont_touch of WX5785: signal is true;
	signal WX5786: std_logic; attribute dont_touch of WX5786: signal is true;
	signal WX5787: std_logic; attribute dont_touch of WX5787: signal is true;
	signal WX5788: std_logic; attribute dont_touch of WX5788: signal is true;
	signal WX5789: std_logic; attribute dont_touch of WX5789: signal is true;
	signal WX5790: std_logic; attribute dont_touch of WX5790: signal is true;
	signal WX5791: std_logic; attribute dont_touch of WX5791: signal is true;
	signal WX5792: std_logic; attribute dont_touch of WX5792: signal is true;
	signal WX5793: std_logic; attribute dont_touch of WX5793: signal is true;
	signal WX5794: std_logic; attribute dont_touch of WX5794: signal is true;
	signal WX5795: std_logic; attribute dont_touch of WX5795: signal is true;
	signal WX5796: std_logic; attribute dont_touch of WX5796: signal is true;
	signal WX5797: std_logic; attribute dont_touch of WX5797: signal is true;
	signal WX5798: std_logic; attribute dont_touch of WX5798: signal is true;
	signal WX5799: std_logic; attribute dont_touch of WX5799: signal is true;
	signal WX5800: std_logic; attribute dont_touch of WX5800: signal is true;
	signal WX5801: std_logic; attribute dont_touch of WX5801: signal is true;
	signal WX5802: std_logic; attribute dont_touch of WX5802: signal is true;
	signal WX5803: std_logic; attribute dont_touch of WX5803: signal is true;
	signal WX5804: std_logic; attribute dont_touch of WX5804: signal is true;
	signal WX5805: std_logic; attribute dont_touch of WX5805: signal is true;
	signal WX5806: std_logic; attribute dont_touch of WX5806: signal is true;
	signal WX5807: std_logic; attribute dont_touch of WX5807: signal is true;
	signal WX5808: std_logic; attribute dont_touch of WX5808: signal is true;
	signal WX5809: std_logic; attribute dont_touch of WX5809: signal is true;
	signal WX5810: std_logic; attribute dont_touch of WX5810: signal is true;
	signal WX5811: std_logic; attribute dont_touch of WX5811: signal is true;
	signal WX5812: std_logic; attribute dont_touch of WX5812: signal is true;
	signal WX5813: std_logic; attribute dont_touch of WX5813: signal is true;
	signal WX5814: std_logic; attribute dont_touch of WX5814: signal is true;
	signal WX5815: std_logic; attribute dont_touch of WX5815: signal is true;
	signal WX5816: std_logic; attribute dont_touch of WX5816: signal is true;
	signal WX5817: std_logic; attribute dont_touch of WX5817: signal is true;
	signal WX5818: std_logic; attribute dont_touch of WX5818: signal is true;
	signal WX5819: std_logic; attribute dont_touch of WX5819: signal is true;
	signal WX5820: std_logic; attribute dont_touch of WX5820: signal is true;
	signal WX5821: std_logic; attribute dont_touch of WX5821: signal is true;
	signal WX5822: std_logic; attribute dont_touch of WX5822: signal is true;
	signal WX5823: std_logic; attribute dont_touch of WX5823: signal is true;
	signal WX5824: std_logic; attribute dont_touch of WX5824: signal is true;
	signal WX5825: std_logic; attribute dont_touch of WX5825: signal is true;
	signal WX5826: std_logic; attribute dont_touch of WX5826: signal is true;
	signal WX5827: std_logic; attribute dont_touch of WX5827: signal is true;
	signal WX5828: std_logic; attribute dont_touch of WX5828: signal is true;
	signal WX5829: std_logic; attribute dont_touch of WX5829: signal is true;
	signal WX5830: std_logic; attribute dont_touch of WX5830: signal is true;
	signal WX5831: std_logic; attribute dont_touch of WX5831: signal is true;
	signal WX5832: std_logic; attribute dont_touch of WX5832: signal is true;
	signal WX5833: std_logic; attribute dont_touch of WX5833: signal is true;
	signal WX5834: std_logic; attribute dont_touch of WX5834: signal is true;
	signal WX5835: std_logic; attribute dont_touch of WX5835: signal is true;
	signal WX5836: std_logic; attribute dont_touch of WX5836: signal is true;
	signal WX5837: std_logic; attribute dont_touch of WX5837: signal is true;
	signal WX5838: std_logic; attribute dont_touch of WX5838: signal is true;
	signal WX5839: std_logic; attribute dont_touch of WX5839: signal is true;
	signal WX5840: std_logic; attribute dont_touch of WX5840: signal is true;
	signal WX5841: std_logic; attribute dont_touch of WX5841: signal is true;
	signal WX5842: std_logic; attribute dont_touch of WX5842: signal is true;
	signal WX5843: std_logic; attribute dont_touch of WX5843: signal is true;
	signal WX5844: std_logic; attribute dont_touch of WX5844: signal is true;
	signal WX5845: std_logic; attribute dont_touch of WX5845: signal is true;
	signal WX5846: std_logic; attribute dont_touch of WX5846: signal is true;
	signal WX5847: std_logic; attribute dont_touch of WX5847: signal is true;
	signal WX5848: std_logic; attribute dont_touch of WX5848: signal is true;
	signal WX5849: std_logic; attribute dont_touch of WX5849: signal is true;
	signal WX5850: std_logic; attribute dont_touch of WX5850: signal is true;
	signal WX5851: std_logic; attribute dont_touch of WX5851: signal is true;
	signal WX5852: std_logic; attribute dont_touch of WX5852: signal is true;
	signal WX5853: std_logic; attribute dont_touch of WX5853: signal is true;
	signal WX5854: std_logic; attribute dont_touch of WX5854: signal is true;
	signal WX5855: std_logic; attribute dont_touch of WX5855: signal is true;
	signal WX5856: std_logic; attribute dont_touch of WX5856: signal is true;
	signal WX5857: std_logic; attribute dont_touch of WX5857: signal is true;
	signal WX5858: std_logic; attribute dont_touch of WX5858: signal is true;
	signal WX5859: std_logic; attribute dont_touch of WX5859: signal is true;
	signal WX5860: std_logic; attribute dont_touch of WX5860: signal is true;
	signal WX5861: std_logic; attribute dont_touch of WX5861: signal is true;
	signal WX5862: std_logic; attribute dont_touch of WX5862: signal is true;
	signal WX5863: std_logic; attribute dont_touch of WX5863: signal is true;
	signal WX5864: std_logic; attribute dont_touch of WX5864: signal is true;
	signal WX5865: std_logic; attribute dont_touch of WX5865: signal is true;
	signal WX5866: std_logic; attribute dont_touch of WX5866: signal is true;
	signal WX5867: std_logic; attribute dont_touch of WX5867: signal is true;
	signal WX5868: std_logic; attribute dont_touch of WX5868: signal is true;
	signal WX5869: std_logic; attribute dont_touch of WX5869: signal is true;
	signal WX5870: std_logic; attribute dont_touch of WX5870: signal is true;
	signal WX5871: std_logic; attribute dont_touch of WX5871: signal is true;
	signal WX5872: std_logic; attribute dont_touch of WX5872: signal is true;
	signal WX5873: std_logic; attribute dont_touch of WX5873: signal is true;
	signal WX5874: std_logic; attribute dont_touch of WX5874: signal is true;
	signal WX5875: std_logic; attribute dont_touch of WX5875: signal is true;
	signal WX5876: std_logic; attribute dont_touch of WX5876: signal is true;
	signal WX5877: std_logic; attribute dont_touch of WX5877: signal is true;
	signal WX5878: std_logic; attribute dont_touch of WX5878: signal is true;
	signal WX5879: std_logic; attribute dont_touch of WX5879: signal is true;
	signal WX5880: std_logic; attribute dont_touch of WX5880: signal is true;
	signal WX5881: std_logic; attribute dont_touch of WX5881: signal is true;
	signal WX5882: std_logic; attribute dont_touch of WX5882: signal is true;
	signal WX5883: std_logic; attribute dont_touch of WX5883: signal is true;
	signal WX5884: std_logic; attribute dont_touch of WX5884: signal is true;
	signal WX5885: std_logic; attribute dont_touch of WX5885: signal is true;
	signal WX5886: std_logic; attribute dont_touch of WX5886: signal is true;
	signal WX5887: std_logic; attribute dont_touch of WX5887: signal is true;
	signal WX5888: std_logic; attribute dont_touch of WX5888: signal is true;
	signal WX5889: std_logic; attribute dont_touch of WX5889: signal is true;
	signal WX5890: std_logic; attribute dont_touch of WX5890: signal is true;
	signal WX5891: std_logic; attribute dont_touch of WX5891: signal is true;
	signal WX5892: std_logic; attribute dont_touch of WX5892: signal is true;
	signal WX5893: std_logic; attribute dont_touch of WX5893: signal is true;
	signal WX5894: std_logic; attribute dont_touch of WX5894: signal is true;
	signal WX5895: std_logic; attribute dont_touch of WX5895: signal is true;
	signal WX5896: std_logic; attribute dont_touch of WX5896: signal is true;
	signal WX5897: std_logic; attribute dont_touch of WX5897: signal is true;
	signal WX5898: std_logic; attribute dont_touch of WX5898: signal is true;
	signal WX5899: std_logic; attribute dont_touch of WX5899: signal is true;
	signal WX5900: std_logic; attribute dont_touch of WX5900: signal is true;
	signal WX5901: std_logic; attribute dont_touch of WX5901: signal is true;
	signal WX5902: std_logic; attribute dont_touch of WX5902: signal is true;
	signal WX5903: std_logic; attribute dont_touch of WX5903: signal is true;
	signal WX5904: std_logic; attribute dont_touch of WX5904: signal is true;
	signal WX5905: std_logic; attribute dont_touch of WX5905: signal is true;
	signal WX5906: std_logic; attribute dont_touch of WX5906: signal is true;
	signal WX5907: std_logic; attribute dont_touch of WX5907: signal is true;
	signal WX5908: std_logic; attribute dont_touch of WX5908: signal is true;
	signal WX5909: std_logic; attribute dont_touch of WX5909: signal is true;
	signal WX5910: std_logic; attribute dont_touch of WX5910: signal is true;
	signal WX5911: std_logic; attribute dont_touch of WX5911: signal is true;
	signal WX5912: std_logic; attribute dont_touch of WX5912: signal is true;
	signal WX5913: std_logic; attribute dont_touch of WX5913: signal is true;
	signal WX5914: std_logic; attribute dont_touch of WX5914: signal is true;
	signal WX5915: std_logic; attribute dont_touch of WX5915: signal is true;
	signal WX5916: std_logic; attribute dont_touch of WX5916: signal is true;
	signal WX5917: std_logic; attribute dont_touch of WX5917: signal is true;
	signal WX5918: std_logic; attribute dont_touch of WX5918: signal is true;
	signal WX5919: std_logic; attribute dont_touch of WX5919: signal is true;
	signal WX5920: std_logic; attribute dont_touch of WX5920: signal is true;
	signal WX5921: std_logic; attribute dont_touch of WX5921: signal is true;
	signal WX5922: std_logic; attribute dont_touch of WX5922: signal is true;
	signal WX5923: std_logic; attribute dont_touch of WX5923: signal is true;
	signal WX5924: std_logic; attribute dont_touch of WX5924: signal is true;
	signal WX5925: std_logic; attribute dont_touch of WX5925: signal is true;
	signal WX5926: std_logic; attribute dont_touch of WX5926: signal is true;
	signal WX5927: std_logic; attribute dont_touch of WX5927: signal is true;
	signal WX5928: std_logic; attribute dont_touch of WX5928: signal is true;
	signal WX5929: std_logic; attribute dont_touch of WX5929: signal is true;
	signal WX5930: std_logic; attribute dont_touch of WX5930: signal is true;
	signal WX5931: std_logic; attribute dont_touch of WX5931: signal is true;
	signal WX5932: std_logic; attribute dont_touch of WX5932: signal is true;
	signal WX5933: std_logic; attribute dont_touch of WX5933: signal is true;
	signal WX5934: std_logic; attribute dont_touch of WX5934: signal is true;
	signal WX5935: std_logic; attribute dont_touch of WX5935: signal is true;
	signal WX5936: std_logic; attribute dont_touch of WX5936: signal is true;
	signal WX5937: std_logic; attribute dont_touch of WX5937: signal is true;
	signal WX5938: std_logic; attribute dont_touch of WX5938: signal is true;
	signal WX5939: std_logic; attribute dont_touch of WX5939: signal is true;
	signal WX5940: std_logic; attribute dont_touch of WX5940: signal is true;
	signal WX5941: std_logic; attribute dont_touch of WX5941: signal is true;
	signal WX5942: std_logic; attribute dont_touch of WX5942: signal is true;
	signal WX5943: std_logic; attribute dont_touch of WX5943: signal is true;
	signal WX5944: std_logic; attribute dont_touch of WX5944: signal is true;
	signal WX5945: std_logic; attribute dont_touch of WX5945: signal is true;
	signal WX5946: std_logic; attribute dont_touch of WX5946: signal is true;
	signal WX5947: std_logic; attribute dont_touch of WX5947: signal is true;
	signal WX5948: std_logic; attribute dont_touch of WX5948: signal is true;
	signal WX5949: std_logic; attribute dont_touch of WX5949: signal is true;
	signal WX5950: std_logic; attribute dont_touch of WX5950: signal is true;
	signal WX5951: std_logic; attribute dont_touch of WX5951: signal is true;
	signal WX5952: std_logic; attribute dont_touch of WX5952: signal is true;
	signal WX5953: std_logic; attribute dont_touch of WX5953: signal is true;
	signal WX5954: std_logic; attribute dont_touch of WX5954: signal is true;
	signal WX5955: std_logic; attribute dont_touch of WX5955: signal is true;
	signal WX5956: std_logic; attribute dont_touch of WX5956: signal is true;
	signal WX5957: std_logic; attribute dont_touch of WX5957: signal is true;
	signal WX5958: std_logic; attribute dont_touch of WX5958: signal is true;
	signal WX5959: std_logic; attribute dont_touch of WX5959: signal is true;
	signal WX5960: std_logic; attribute dont_touch of WX5960: signal is true;
	signal WX5961: std_logic; attribute dont_touch of WX5961: signal is true;
	signal WX5962: std_logic; attribute dont_touch of WX5962: signal is true;
	signal WX5963: std_logic; attribute dont_touch of WX5963: signal is true;
	signal WX5964: std_logic; attribute dont_touch of WX5964: signal is true;
	signal WX5965: std_logic; attribute dont_touch of WX5965: signal is true;
	signal WX5966: std_logic; attribute dont_touch of WX5966: signal is true;
	signal WX5967: std_logic; attribute dont_touch of WX5967: signal is true;
	signal WX5968: std_logic; attribute dont_touch of WX5968: signal is true;
	signal WX5969: std_logic; attribute dont_touch of WX5969: signal is true;
	signal WX5970: std_logic; attribute dont_touch of WX5970: signal is true;
	signal WX5971: std_logic; attribute dont_touch of WX5971: signal is true;
	signal WX5972: std_logic; attribute dont_touch of WX5972: signal is true;
	signal WX5973: std_logic; attribute dont_touch of WX5973: signal is true;
	signal WX5974: std_logic; attribute dont_touch of WX5974: signal is true;
	signal WX5975: std_logic; attribute dont_touch of WX5975: signal is true;
	signal WX5976: std_logic; attribute dont_touch of WX5976: signal is true;
	signal WX5977: std_logic; attribute dont_touch of WX5977: signal is true;
	signal WX5978: std_logic; attribute dont_touch of WX5978: signal is true;
	signal WX5979: std_logic; attribute dont_touch of WX5979: signal is true;
	signal WX5980: std_logic; attribute dont_touch of WX5980: signal is true;
	signal WX5981: std_logic; attribute dont_touch of WX5981: signal is true;
	signal WX5982: std_logic; attribute dont_touch of WX5982: signal is true;
	signal WX5983: std_logic; attribute dont_touch of WX5983: signal is true;
	signal WX5984: std_logic; attribute dont_touch of WX5984: signal is true;
	signal WX5985: std_logic; attribute dont_touch of WX5985: signal is true;
	signal WX5986: std_logic; attribute dont_touch of WX5986: signal is true;
	signal WX5987: std_logic; attribute dont_touch of WX5987: signal is true;
	signal WX5988: std_logic; attribute dont_touch of WX5988: signal is true;
	signal WX5989: std_logic; attribute dont_touch of WX5989: signal is true;
	signal WX5990: std_logic; attribute dont_touch of WX5990: signal is true;
	signal WX5991: std_logic; attribute dont_touch of WX5991: signal is true;
	signal WX5992: std_logic; attribute dont_touch of WX5992: signal is true;
	signal WX5993: std_logic; attribute dont_touch of WX5993: signal is true;
	signal WX5994: std_logic; attribute dont_touch of WX5994: signal is true;
	signal WX5995: std_logic; attribute dont_touch of WX5995: signal is true;
	signal WX5996: std_logic; attribute dont_touch of WX5996: signal is true;
	signal WX5997: std_logic; attribute dont_touch of WX5997: signal is true;
	signal WX5998: std_logic; attribute dont_touch of WX5998: signal is true;
	signal WX5999: std_logic; attribute dont_touch of WX5999: signal is true;
	signal WX6000: std_logic; attribute dont_touch of WX6000: signal is true;
	signal WX6001: std_logic; attribute dont_touch of WX6001: signal is true;
	signal WX6002: std_logic; attribute dont_touch of WX6002: signal is true;
	signal WX6003: std_logic; attribute dont_touch of WX6003: signal is true;
	signal WX6004: std_logic; attribute dont_touch of WX6004: signal is true;
	signal WX6005: std_logic; attribute dont_touch of WX6005: signal is true;
	signal WX6006: std_logic; attribute dont_touch of WX6006: signal is true;
	signal WX6007: std_logic; attribute dont_touch of WX6007: signal is true;
	signal WX6008: std_logic; attribute dont_touch of WX6008: signal is true;
	signal WX6009: std_logic; attribute dont_touch of WX6009: signal is true;
	signal WX6010: std_logic; attribute dont_touch of WX6010: signal is true;
	signal WX6011: std_logic; attribute dont_touch of WX6011: signal is true;
	signal WX6012: std_logic; attribute dont_touch of WX6012: signal is true;
	signal WX6013: std_logic; attribute dont_touch of WX6013: signal is true;
	signal WX6014: std_logic; attribute dont_touch of WX6014: signal is true;
	signal WX6015: std_logic; attribute dont_touch of WX6015: signal is true;
	signal WX6016: std_logic; attribute dont_touch of WX6016: signal is true;
	signal WX6017: std_logic; attribute dont_touch of WX6017: signal is true;
	signal WX6018: std_logic; attribute dont_touch of WX6018: signal is true;
	signal WX6019: std_logic; attribute dont_touch of WX6019: signal is true;
	signal WX6020: std_logic; attribute dont_touch of WX6020: signal is true;
	signal WX6021: std_logic; attribute dont_touch of WX6021: signal is true;
	signal WX6022: std_logic; attribute dont_touch of WX6022: signal is true;
	signal WX6023: std_logic; attribute dont_touch of WX6023: signal is true;
	signal WX6024: std_logic; attribute dont_touch of WX6024: signal is true;
	signal WX6025: std_logic; attribute dont_touch of WX6025: signal is true;
	signal WX6026: std_logic; attribute dont_touch of WX6026: signal is true;
	signal WX6027: std_logic; attribute dont_touch of WX6027: signal is true;
	signal WX6028: std_logic; attribute dont_touch of WX6028: signal is true;
	signal WX6029: std_logic; attribute dont_touch of WX6029: signal is true;
	signal WX6030: std_logic; attribute dont_touch of WX6030: signal is true;
	signal WX6031: std_logic; attribute dont_touch of WX6031: signal is true;
	signal WX6032: std_logic; attribute dont_touch of WX6032: signal is true;
	signal WX6033: std_logic; attribute dont_touch of WX6033: signal is true;
	signal WX6034: std_logic; attribute dont_touch of WX6034: signal is true;
	signal WX6035: std_logic; attribute dont_touch of WX6035: signal is true;
	signal WX6036: std_logic; attribute dont_touch of WX6036: signal is true;
	signal WX6037: std_logic; attribute dont_touch of WX6037: signal is true;
	signal WX6038: std_logic; attribute dont_touch of WX6038: signal is true;
	signal WX6039: std_logic; attribute dont_touch of WX6039: signal is true;
	signal WX6040: std_logic; attribute dont_touch of WX6040: signal is true;
	signal WX6041: std_logic; attribute dont_touch of WX6041: signal is true;
	signal WX6042: std_logic; attribute dont_touch of WX6042: signal is true;
	signal WX6043: std_logic; attribute dont_touch of WX6043: signal is true;
	signal WX6044: std_logic; attribute dont_touch of WX6044: signal is true;
	signal WX6045: std_logic; attribute dont_touch of WX6045: signal is true;
	signal WX6046: std_logic; attribute dont_touch of WX6046: signal is true;
	signal WX6047: std_logic; attribute dont_touch of WX6047: signal is true;
	signal WX6048: std_logic; attribute dont_touch of WX6048: signal is true;
	signal WX6049: std_logic; attribute dont_touch of WX6049: signal is true;
	signal WX6050: std_logic; attribute dont_touch of WX6050: signal is true;
	signal WX6051: std_logic; attribute dont_touch of WX6051: signal is true;
	signal WX6052: std_logic; attribute dont_touch of WX6052: signal is true;
	signal WX6053: std_logic; attribute dont_touch of WX6053: signal is true;
	signal WX6054: std_logic; attribute dont_touch of WX6054: signal is true;
	signal WX6055: std_logic; attribute dont_touch of WX6055: signal is true;
	signal WX6056: std_logic; attribute dont_touch of WX6056: signal is true;
	signal WX6057: std_logic; attribute dont_touch of WX6057: signal is true;
	signal WX6058: std_logic; attribute dont_touch of WX6058: signal is true;
	signal WX6059: std_logic; attribute dont_touch of WX6059: signal is true;
	signal WX6060: std_logic; attribute dont_touch of WX6060: signal is true;
	signal WX6061: std_logic; attribute dont_touch of WX6061: signal is true;
	signal WX6062: std_logic; attribute dont_touch of WX6062: signal is true;
	signal WX6063: std_logic; attribute dont_touch of WX6063: signal is true;
	signal WX6064: std_logic; attribute dont_touch of WX6064: signal is true;
	signal WX6065: std_logic; attribute dont_touch of WX6065: signal is true;
	signal WX6066: std_logic; attribute dont_touch of WX6066: signal is true;
	signal WX6067: std_logic; attribute dont_touch of WX6067: signal is true;
	signal WX6068: std_logic; attribute dont_touch of WX6068: signal is true;
	signal WX6069: std_logic; attribute dont_touch of WX6069: signal is true;
	signal WX6070: std_logic; attribute dont_touch of WX6070: signal is true;
	signal WX6071: std_logic; attribute dont_touch of WX6071: signal is true;
	signal WX6072: std_logic; attribute dont_touch of WX6072: signal is true;
	signal WX6073: std_logic; attribute dont_touch of WX6073: signal is true;
	signal WX6074: std_logic; attribute dont_touch of WX6074: signal is true;
	signal WX6075: std_logic; attribute dont_touch of WX6075: signal is true;
	signal WX6076: std_logic; attribute dont_touch of WX6076: signal is true;
	signal WX6077: std_logic; attribute dont_touch of WX6077: signal is true;
	signal WX6078: std_logic; attribute dont_touch of WX6078: signal is true;
	signal WX6079: std_logic; attribute dont_touch of WX6079: signal is true;
	signal WX6080: std_logic; attribute dont_touch of WX6080: signal is true;
	signal WX6081: std_logic; attribute dont_touch of WX6081: signal is true;
	signal WX6082: std_logic; attribute dont_touch of WX6082: signal is true;
	signal WX6083: std_logic; attribute dont_touch of WX6083: signal is true;
	signal WX6084: std_logic; attribute dont_touch of WX6084: signal is true;
	signal WX6085: std_logic; attribute dont_touch of WX6085: signal is true;
	signal WX6086: std_logic; attribute dont_touch of WX6086: signal is true;
	signal WX6087: std_logic; attribute dont_touch of WX6087: signal is true;
	signal WX6088: std_logic; attribute dont_touch of WX6088: signal is true;
	signal WX6089: std_logic; attribute dont_touch of WX6089: signal is true;
	signal WX6090: std_logic; attribute dont_touch of WX6090: signal is true;
	signal WX6091: std_logic; attribute dont_touch of WX6091: signal is true;
	signal WX6092: std_logic; attribute dont_touch of WX6092: signal is true;
	signal WX6093: std_logic; attribute dont_touch of WX6093: signal is true;
	signal WX6094: std_logic; attribute dont_touch of WX6094: signal is true;
	signal WX6095: std_logic; attribute dont_touch of WX6095: signal is true;
	signal WX6096: std_logic; attribute dont_touch of WX6096: signal is true;
	signal WX6097: std_logic; attribute dont_touch of WX6097: signal is true;
	signal WX6098: std_logic; attribute dont_touch of WX6098: signal is true;
	signal WX6099: std_logic; attribute dont_touch of WX6099: signal is true;
	signal WX6100: std_logic; attribute dont_touch of WX6100: signal is true;
	signal WX6101: std_logic; attribute dont_touch of WX6101: signal is true;
	signal WX6102: std_logic; attribute dont_touch of WX6102: signal is true;
	signal WX6103: std_logic; attribute dont_touch of WX6103: signal is true;
	signal WX6104: std_logic; attribute dont_touch of WX6104: signal is true;
	signal WX6105: std_logic; attribute dont_touch of WX6105: signal is true;
	signal WX6106: std_logic; attribute dont_touch of WX6106: signal is true;
	signal WX6107: std_logic; attribute dont_touch of WX6107: signal is true;
	signal WX6108: std_logic; attribute dont_touch of WX6108: signal is true;
	signal WX6109: std_logic; attribute dont_touch of WX6109: signal is true;
	signal WX6110: std_logic; attribute dont_touch of WX6110: signal is true;
	signal WX6111: std_logic; attribute dont_touch of WX6111: signal is true;
	signal WX6112: std_logic; attribute dont_touch of WX6112: signal is true;
	signal WX6113: std_logic; attribute dont_touch of WX6113: signal is true;
	signal WX6114: std_logic; attribute dont_touch of WX6114: signal is true;
	signal WX6115: std_logic; attribute dont_touch of WX6115: signal is true;
	signal WX6116: std_logic; attribute dont_touch of WX6116: signal is true;
	signal WX6117: std_logic; attribute dont_touch of WX6117: signal is true;
	signal WX6118: std_logic; attribute dont_touch of WX6118: signal is true;
	signal WX6119: std_logic; attribute dont_touch of WX6119: signal is true;
	signal WX6120: std_logic; attribute dont_touch of WX6120: signal is true;
	signal WX6121: std_logic; attribute dont_touch of WX6121: signal is true;
	signal WX6122: std_logic; attribute dont_touch of WX6122: signal is true;
	signal WX6123: std_logic; attribute dont_touch of WX6123: signal is true;
	signal WX6124: std_logic; attribute dont_touch of WX6124: signal is true;
	signal WX6125: std_logic; attribute dont_touch of WX6125: signal is true;
	signal WX6126: std_logic; attribute dont_touch of WX6126: signal is true;
	signal WX6127: std_logic; attribute dont_touch of WX6127: signal is true;
	signal WX6128: std_logic; attribute dont_touch of WX6128: signal is true;
	signal WX6129: std_logic; attribute dont_touch of WX6129: signal is true;
	signal WX6130: std_logic; attribute dont_touch of WX6130: signal is true;
	signal WX6131: std_logic; attribute dont_touch of WX6131: signal is true;
	signal WX6132: std_logic; attribute dont_touch of WX6132: signal is true;
	signal WX6133: std_logic; attribute dont_touch of WX6133: signal is true;
	signal WX6134: std_logic; attribute dont_touch of WX6134: signal is true;
	signal WX6135: std_logic; attribute dont_touch of WX6135: signal is true;
	signal WX6136: std_logic; attribute dont_touch of WX6136: signal is true;
	signal WX6137: std_logic; attribute dont_touch of WX6137: signal is true;
	signal WX6138: std_logic; attribute dont_touch of WX6138: signal is true;
	signal WX6139: std_logic; attribute dont_touch of WX6139: signal is true;
	signal WX6140: std_logic; attribute dont_touch of WX6140: signal is true;
	signal WX6141: std_logic; attribute dont_touch of WX6141: signal is true;
	signal WX6142: std_logic; attribute dont_touch of WX6142: signal is true;
	signal WX6143: std_logic; attribute dont_touch of WX6143: signal is true;
	signal WX6144: std_logic; attribute dont_touch of WX6144: signal is true;
	signal WX6145: std_logic; attribute dont_touch of WX6145: signal is true;
	signal WX6146: std_logic; attribute dont_touch of WX6146: signal is true;
	signal WX6147: std_logic; attribute dont_touch of WX6147: signal is true;
	signal WX6148: std_logic; attribute dont_touch of WX6148: signal is true;
	signal WX6149: std_logic; attribute dont_touch of WX6149: signal is true;
	signal WX6150: std_logic; attribute dont_touch of WX6150: signal is true;
	signal WX6151: std_logic; attribute dont_touch of WX6151: signal is true;
	signal WX6152: std_logic; attribute dont_touch of WX6152: signal is true;
	signal WX6153: std_logic; attribute dont_touch of WX6153: signal is true;
	signal WX6154: std_logic; attribute dont_touch of WX6154: signal is true;
	signal WX6155: std_logic; attribute dont_touch of WX6155: signal is true;
	signal WX6156: std_logic; attribute dont_touch of WX6156: signal is true;
	signal WX6157: std_logic; attribute dont_touch of WX6157: signal is true;
	signal WX6158: std_logic; attribute dont_touch of WX6158: signal is true;
	signal WX6159: std_logic; attribute dont_touch of WX6159: signal is true;
	signal WX6160: std_logic; attribute dont_touch of WX6160: signal is true;
	signal WX6161: std_logic; attribute dont_touch of WX6161: signal is true;
	signal WX6162: std_logic; attribute dont_touch of WX6162: signal is true;
	signal WX6163: std_logic; attribute dont_touch of WX6163: signal is true;
	signal WX6164: std_logic; attribute dont_touch of WX6164: signal is true;
	signal WX6165: std_logic; attribute dont_touch of WX6165: signal is true;
	signal WX6166: std_logic; attribute dont_touch of WX6166: signal is true;
	signal WX6167: std_logic; attribute dont_touch of WX6167: signal is true;
	signal WX6168: std_logic; attribute dont_touch of WX6168: signal is true;
	signal WX6169: std_logic; attribute dont_touch of WX6169: signal is true;
	signal WX6170: std_logic; attribute dont_touch of WX6170: signal is true;
	signal WX6171: std_logic; attribute dont_touch of WX6171: signal is true;
	signal WX6172: std_logic; attribute dont_touch of WX6172: signal is true;
	signal WX6173: std_logic; attribute dont_touch of WX6173: signal is true;
	signal WX6174: std_logic; attribute dont_touch of WX6174: signal is true;
	signal WX6175: std_logic; attribute dont_touch of WX6175: signal is true;
	signal WX6176: std_logic; attribute dont_touch of WX6176: signal is true;
	signal WX6177: std_logic; attribute dont_touch of WX6177: signal is true;
	signal WX6178: std_logic; attribute dont_touch of WX6178: signal is true;
	signal WX6179: std_logic; attribute dont_touch of WX6179: signal is true;
	signal WX6180: std_logic; attribute dont_touch of WX6180: signal is true;
	signal WX6181: std_logic; attribute dont_touch of WX6181: signal is true;
	signal WX6182: std_logic; attribute dont_touch of WX6182: signal is true;
	signal WX6183: std_logic; attribute dont_touch of WX6183: signal is true;
	signal WX6184: std_logic; attribute dont_touch of WX6184: signal is true;
	signal WX6185: std_logic; attribute dont_touch of WX6185: signal is true;
	signal WX6186: std_logic; attribute dont_touch of WX6186: signal is true;
	signal WX6187: std_logic; attribute dont_touch of WX6187: signal is true;
	signal WX6188: std_logic; attribute dont_touch of WX6188: signal is true;
	signal WX6189: std_logic; attribute dont_touch of WX6189: signal is true;
	signal WX6190: std_logic; attribute dont_touch of WX6190: signal is true;
	signal WX6191: std_logic; attribute dont_touch of WX6191: signal is true;
	signal WX6192: std_logic; attribute dont_touch of WX6192: signal is true;
	signal WX6193: std_logic; attribute dont_touch of WX6193: signal is true;
	signal WX6194: std_logic; attribute dont_touch of WX6194: signal is true;
	signal WX6195: std_logic; attribute dont_touch of WX6195: signal is true;
	signal WX6196: std_logic; attribute dont_touch of WX6196: signal is true;
	signal WX6197: std_logic; attribute dont_touch of WX6197: signal is true;
	signal WX6198: std_logic; attribute dont_touch of WX6198: signal is true;
	signal WX6199: std_logic; attribute dont_touch of WX6199: signal is true;
	signal WX6200: std_logic; attribute dont_touch of WX6200: signal is true;
	signal WX6201: std_logic; attribute dont_touch of WX6201: signal is true;
	signal WX6202: std_logic; attribute dont_touch of WX6202: signal is true;
	signal WX6203: std_logic; attribute dont_touch of WX6203: signal is true;
	signal WX6204: std_logic; attribute dont_touch of WX6204: signal is true;
	signal WX6205: std_logic; attribute dont_touch of WX6205: signal is true;
	signal WX6206: std_logic; attribute dont_touch of WX6206: signal is true;
	signal WX6207: std_logic; attribute dont_touch of WX6207: signal is true;
	signal WX6208: std_logic; attribute dont_touch of WX6208: signal is true;
	signal WX6209: std_logic; attribute dont_touch of WX6209: signal is true;
	signal WX6210: std_logic; attribute dont_touch of WX6210: signal is true;
	signal WX6211: std_logic; attribute dont_touch of WX6211: signal is true;
	signal WX6212: std_logic; attribute dont_touch of WX6212: signal is true;
	signal WX6213: std_logic; attribute dont_touch of WX6213: signal is true;
	signal WX6214: std_logic; attribute dont_touch of WX6214: signal is true;
	signal WX6215: std_logic; attribute dont_touch of WX6215: signal is true;
	signal WX6216: std_logic; attribute dont_touch of WX6216: signal is true;
	signal WX6217: std_logic; attribute dont_touch of WX6217: signal is true;
	signal WX6218: std_logic; attribute dont_touch of WX6218: signal is true;
	signal WX6219: std_logic; attribute dont_touch of WX6219: signal is true;
	signal WX6220: std_logic; attribute dont_touch of WX6220: signal is true;
	signal WX6221: std_logic; attribute dont_touch of WX6221: signal is true;
	signal WX6222: std_logic; attribute dont_touch of WX6222: signal is true;
	signal WX6223: std_logic; attribute dont_touch of WX6223: signal is true;
	signal WX6224: std_logic; attribute dont_touch of WX6224: signal is true;
	signal WX6225: std_logic; attribute dont_touch of WX6225: signal is true;
	signal WX6226: std_logic; attribute dont_touch of WX6226: signal is true;
	signal WX6227: std_logic; attribute dont_touch of WX6227: signal is true;
	signal WX6228: std_logic; attribute dont_touch of WX6228: signal is true;
	signal WX6229: std_logic; attribute dont_touch of WX6229: signal is true;
	signal WX6230: std_logic; attribute dont_touch of WX6230: signal is true;
	signal WX6231: std_logic; attribute dont_touch of WX6231: signal is true;
	signal WX6232: std_logic; attribute dont_touch of WX6232: signal is true;
	signal WX6233: std_logic; attribute dont_touch of WX6233: signal is true;
	signal WX6234: std_logic; attribute dont_touch of WX6234: signal is true;
	signal WX6235: std_logic; attribute dont_touch of WX6235: signal is true;
	signal WX6236: std_logic; attribute dont_touch of WX6236: signal is true;
	signal WX6237: std_logic; attribute dont_touch of WX6237: signal is true;
	signal WX6238: std_logic; attribute dont_touch of WX6238: signal is true;
	signal WX6239: std_logic; attribute dont_touch of WX6239: signal is true;
	signal WX6240: std_logic; attribute dont_touch of WX6240: signal is true;
	signal WX6241: std_logic; attribute dont_touch of WX6241: signal is true;
	signal WX6242: std_logic; attribute dont_touch of WX6242: signal is true;
	signal WX6243: std_logic; attribute dont_touch of WX6243: signal is true;
	signal WX6244: std_logic; attribute dont_touch of WX6244: signal is true;
	signal WX6245: std_logic; attribute dont_touch of WX6245: signal is true;
	signal WX6246: std_logic; attribute dont_touch of WX6246: signal is true;
	signal WX6247: std_logic; attribute dont_touch of WX6247: signal is true;
	signal WX6248: std_logic; attribute dont_touch of WX6248: signal is true;
	signal WX6249: std_logic; attribute dont_touch of WX6249: signal is true;
	signal WX6250: std_logic; attribute dont_touch of WX6250: signal is true;
	signal WX6251: std_logic; attribute dont_touch of WX6251: signal is true;
	signal WX6252: std_logic; attribute dont_touch of WX6252: signal is true;
	signal WX6253: std_logic; attribute dont_touch of WX6253: signal is true;
	signal WX6254: std_logic; attribute dont_touch of WX6254: signal is true;
	signal WX6255: std_logic; attribute dont_touch of WX6255: signal is true;
	signal WX6256: std_logic; attribute dont_touch of WX6256: signal is true;
	signal WX6257: std_logic; attribute dont_touch of WX6257: signal is true;
	signal WX6258: std_logic; attribute dont_touch of WX6258: signal is true;
	signal WX6259: std_logic; attribute dont_touch of WX6259: signal is true;
	signal WX6260: std_logic; attribute dont_touch of WX6260: signal is true;
	signal WX6261: std_logic; attribute dont_touch of WX6261: signal is true;
	signal WX6262: std_logic; attribute dont_touch of WX6262: signal is true;
	signal WX6263: std_logic; attribute dont_touch of WX6263: signal is true;
	signal WX6264: std_logic; attribute dont_touch of WX6264: signal is true;
	signal WX6265: std_logic; attribute dont_touch of WX6265: signal is true;
	signal WX6266: std_logic; attribute dont_touch of WX6266: signal is true;
	signal WX6267: std_logic; attribute dont_touch of WX6267: signal is true;
	signal WX6268: std_logic; attribute dont_touch of WX6268: signal is true;
	signal WX6269: std_logic; attribute dont_touch of WX6269: signal is true;
	signal WX6270: std_logic; attribute dont_touch of WX6270: signal is true;
	signal WX6271: std_logic; attribute dont_touch of WX6271: signal is true;
	signal WX6272: std_logic; attribute dont_touch of WX6272: signal is true;
	signal WX6273: std_logic; attribute dont_touch of WX6273: signal is true;
	signal WX6274: std_logic; attribute dont_touch of WX6274: signal is true;
	signal WX6275: std_logic; attribute dont_touch of WX6275: signal is true;
	signal WX6276: std_logic; attribute dont_touch of WX6276: signal is true;
	signal WX6277: std_logic; attribute dont_touch of WX6277: signal is true;
	signal WX6278: std_logic; attribute dont_touch of WX6278: signal is true;
	signal WX6279: std_logic; attribute dont_touch of WX6279: signal is true;
	signal WX6280: std_logic; attribute dont_touch of WX6280: signal is true;
	signal WX6281: std_logic; attribute dont_touch of WX6281: signal is true;
	signal WX6282: std_logic; attribute dont_touch of WX6282: signal is true;
	signal WX6283: std_logic; attribute dont_touch of WX6283: signal is true;
	signal WX6284: std_logic; attribute dont_touch of WX6284: signal is true;
	signal WX6285: std_logic; attribute dont_touch of WX6285: signal is true;
	signal WX6286: std_logic; attribute dont_touch of WX6286: signal is true;
	signal WX6287: std_logic; attribute dont_touch of WX6287: signal is true;
	signal WX6288: std_logic; attribute dont_touch of WX6288: signal is true;
	signal WX6289: std_logic; attribute dont_touch of WX6289: signal is true;
	signal WX6290: std_logic; attribute dont_touch of WX6290: signal is true;
	signal WX6291: std_logic; attribute dont_touch of WX6291: signal is true;
	signal WX6292: std_logic; attribute dont_touch of WX6292: signal is true;
	signal WX6293: std_logic; attribute dont_touch of WX6293: signal is true;
	signal WX6294: std_logic; attribute dont_touch of WX6294: signal is true;
	signal WX6295: std_logic; attribute dont_touch of WX6295: signal is true;
	signal WX6296: std_logic; attribute dont_touch of WX6296: signal is true;
	signal WX6297: std_logic; attribute dont_touch of WX6297: signal is true;
	signal WX6298: std_logic; attribute dont_touch of WX6298: signal is true;
	signal WX6299: std_logic; attribute dont_touch of WX6299: signal is true;
	signal WX6300: std_logic; attribute dont_touch of WX6300: signal is true;
	signal WX6301: std_logic; attribute dont_touch of WX6301: signal is true;
	signal WX6302: std_logic; attribute dont_touch of WX6302: signal is true;
	signal WX6303: std_logic; attribute dont_touch of WX6303: signal is true;
	signal WX6304: std_logic; attribute dont_touch of WX6304: signal is true;
	signal WX6305: std_logic; attribute dont_touch of WX6305: signal is true;
	signal WX6306: std_logic; attribute dont_touch of WX6306: signal is true;
	signal WX6307: std_logic; attribute dont_touch of WX6307: signal is true;
	signal WX6308: std_logic; attribute dont_touch of WX6308: signal is true;
	signal WX6309: std_logic; attribute dont_touch of WX6309: signal is true;
	signal WX6310: std_logic; attribute dont_touch of WX6310: signal is true;
	signal WX6311: std_logic; attribute dont_touch of WX6311: signal is true;
	signal WX6312: std_logic; attribute dont_touch of WX6312: signal is true;
	signal WX6313: std_logic; attribute dont_touch of WX6313: signal is true;
	signal WX6314: std_logic; attribute dont_touch of WX6314: signal is true;
	signal WX6315: std_logic; attribute dont_touch of WX6315: signal is true;
	signal WX6316: std_logic; attribute dont_touch of WX6316: signal is true;
	signal WX6317: std_logic; attribute dont_touch of WX6317: signal is true;
	signal WX6318: std_logic; attribute dont_touch of WX6318: signal is true;
	signal WX6319: std_logic; attribute dont_touch of WX6319: signal is true;
	signal WX6320: std_logic; attribute dont_touch of WX6320: signal is true;
	signal WX6321: std_logic; attribute dont_touch of WX6321: signal is true;
	signal WX6322: std_logic; attribute dont_touch of WX6322: signal is true;
	signal WX6323: std_logic; attribute dont_touch of WX6323: signal is true;
	signal WX6324: std_logic; attribute dont_touch of WX6324: signal is true;
	signal WX6325: std_logic; attribute dont_touch of WX6325: signal is true;
	signal WX6326: std_logic; attribute dont_touch of WX6326: signal is true;
	signal WX6327: std_logic; attribute dont_touch of WX6327: signal is true;
	signal WX6328: std_logic; attribute dont_touch of WX6328: signal is true;
	signal WX6329: std_logic; attribute dont_touch of WX6329: signal is true;
	signal WX6330: std_logic; attribute dont_touch of WX6330: signal is true;
	signal WX6331: std_logic; attribute dont_touch of WX6331: signal is true;
	signal WX6332: std_logic; attribute dont_touch of WX6332: signal is true;
	signal WX6333: std_logic; attribute dont_touch of WX6333: signal is true;
	signal WX6334: std_logic; attribute dont_touch of WX6334: signal is true;
	signal WX6335: std_logic; attribute dont_touch of WX6335: signal is true;
	signal WX6336: std_logic; attribute dont_touch of WX6336: signal is true;
	signal WX6337: std_logic; attribute dont_touch of WX6337: signal is true;
	signal WX6338: std_logic; attribute dont_touch of WX6338: signal is true;
	signal WX6339: std_logic; attribute dont_touch of WX6339: signal is true;
	signal WX6340: std_logic; attribute dont_touch of WX6340: signal is true;
	signal WX6341: std_logic; attribute dont_touch of WX6341: signal is true;
	signal WX6342: std_logic; attribute dont_touch of WX6342: signal is true;
	signal WX6343: std_logic; attribute dont_touch of WX6343: signal is true;
	signal WX6344: std_logic; attribute dont_touch of WX6344: signal is true;
	signal WX6345: std_logic; attribute dont_touch of WX6345: signal is true;
	signal WX6346: std_logic; attribute dont_touch of WX6346: signal is true;
	signal WX6347: std_logic; attribute dont_touch of WX6347: signal is true;
	signal WX6348: std_logic; attribute dont_touch of WX6348: signal is true;
	signal WX6349: std_logic; attribute dont_touch of WX6349: signal is true;
	signal WX6350: std_logic; attribute dont_touch of WX6350: signal is true;
	signal WX6351: std_logic; attribute dont_touch of WX6351: signal is true;
	signal WX6352: std_logic; attribute dont_touch of WX6352: signal is true;
	signal WX6353: std_logic; attribute dont_touch of WX6353: signal is true;
	signal WX6354: std_logic; attribute dont_touch of WX6354: signal is true;
	signal WX6355: std_logic; attribute dont_touch of WX6355: signal is true;
	signal WX6356: std_logic; attribute dont_touch of WX6356: signal is true;
	signal WX6357: std_logic; attribute dont_touch of WX6357: signal is true;
	signal WX6358: std_logic; attribute dont_touch of WX6358: signal is true;
	signal WX6359: std_logic; attribute dont_touch of WX6359: signal is true;
	signal WX6360: std_logic; attribute dont_touch of WX6360: signal is true;
	signal WX6361: std_logic; attribute dont_touch of WX6361: signal is true;
	signal WX6362: std_logic; attribute dont_touch of WX6362: signal is true;
	signal WX6363: std_logic; attribute dont_touch of WX6363: signal is true;
	signal WX6364: std_logic; attribute dont_touch of WX6364: signal is true;
	signal WX6365: std_logic; attribute dont_touch of WX6365: signal is true;
	signal WX6366: std_logic; attribute dont_touch of WX6366: signal is true;
	signal WX6367: std_logic; attribute dont_touch of WX6367: signal is true;
	signal WX6368: std_logic; attribute dont_touch of WX6368: signal is true;
	signal WX6369: std_logic; attribute dont_touch of WX6369: signal is true;
	signal WX6370: std_logic; attribute dont_touch of WX6370: signal is true;
	signal WX6371: std_logic; attribute dont_touch of WX6371: signal is true;
	signal WX6372: std_logic; attribute dont_touch of WX6372: signal is true;
	signal WX6373: std_logic; attribute dont_touch of WX6373: signal is true;
	signal WX6374: std_logic; attribute dont_touch of WX6374: signal is true;
	signal WX6375: std_logic; attribute dont_touch of WX6375: signal is true;
	signal WX6376: std_logic; attribute dont_touch of WX6376: signal is true;
	signal WX6377: std_logic; attribute dont_touch of WX6377: signal is true;
	signal WX6378: std_logic; attribute dont_touch of WX6378: signal is true;
	signal WX6379: std_logic; attribute dont_touch of WX6379: signal is true;
	signal WX6380: std_logic; attribute dont_touch of WX6380: signal is true;
	signal WX6381: std_logic; attribute dont_touch of WX6381: signal is true;
	signal WX6382: std_logic; attribute dont_touch of WX6382: signal is true;
	signal WX6383: std_logic; attribute dont_touch of WX6383: signal is true;
	signal WX6384: std_logic; attribute dont_touch of WX6384: signal is true;
	signal WX6385: std_logic; attribute dont_touch of WX6385: signal is true;
	signal WX6386: std_logic; attribute dont_touch of WX6386: signal is true;
	signal WX6387: std_logic; attribute dont_touch of WX6387: signal is true;
	signal WX6388: std_logic; attribute dont_touch of WX6388: signal is true;
	signal WX6389: std_logic; attribute dont_touch of WX6389: signal is true;
	signal WX6390: std_logic; attribute dont_touch of WX6390: signal is true;
	signal WX6391: std_logic; attribute dont_touch of WX6391: signal is true;
	signal WX6392: std_logic; attribute dont_touch of WX6392: signal is true;
	signal WX6393: std_logic; attribute dont_touch of WX6393: signal is true;
	signal WX6394: std_logic; attribute dont_touch of WX6394: signal is true;
	signal WX6395: std_logic; attribute dont_touch of WX6395: signal is true;
	signal WX6396: std_logic; attribute dont_touch of WX6396: signal is true;
	signal WX6397: std_logic; attribute dont_touch of WX6397: signal is true;
	signal WX6398: std_logic; attribute dont_touch of WX6398: signal is true;
	signal WX6399: std_logic; attribute dont_touch of WX6399: signal is true;
	signal WX6400: std_logic; attribute dont_touch of WX6400: signal is true;
	signal WX6401: std_logic; attribute dont_touch of WX6401: signal is true;
	signal WX6402: std_logic; attribute dont_touch of WX6402: signal is true;
	signal WX6403: std_logic; attribute dont_touch of WX6403: signal is true;
	signal WX6404: std_logic; attribute dont_touch of WX6404: signal is true;
	signal WX6405: std_logic; attribute dont_touch of WX6405: signal is true;
	signal WX6406: std_logic; attribute dont_touch of WX6406: signal is true;
	signal WX6407: std_logic; attribute dont_touch of WX6407: signal is true;
	signal WX6408: std_logic; attribute dont_touch of WX6408: signal is true;
	signal WX6409: std_logic; attribute dont_touch of WX6409: signal is true;
	signal WX6410: std_logic; attribute dont_touch of WX6410: signal is true;
	signal WX6411: std_logic; attribute dont_touch of WX6411: signal is true;
	signal WX6412: std_logic; attribute dont_touch of WX6412: signal is true;
	signal WX6413: std_logic; attribute dont_touch of WX6413: signal is true;
	signal WX6414: std_logic; attribute dont_touch of WX6414: signal is true;
	signal WX6415: std_logic; attribute dont_touch of WX6415: signal is true;
	signal WX6416: std_logic; attribute dont_touch of WX6416: signal is true;
	signal WX6417: std_logic; attribute dont_touch of WX6417: signal is true;
	signal WX6418: std_logic; attribute dont_touch of WX6418: signal is true;
	signal WX6419: std_logic; attribute dont_touch of WX6419: signal is true;
	signal WX6420: std_logic; attribute dont_touch of WX6420: signal is true;
	signal WX6421: std_logic; attribute dont_touch of WX6421: signal is true;
	signal WX6422: std_logic; attribute dont_touch of WX6422: signal is true;
	signal WX6423: std_logic; attribute dont_touch of WX6423: signal is true;
	signal WX6424: std_logic; attribute dont_touch of WX6424: signal is true;
	signal WX6425: std_logic; attribute dont_touch of WX6425: signal is true;
	signal WX6426: std_logic; attribute dont_touch of WX6426: signal is true;
	signal WX6427: std_logic; attribute dont_touch of WX6427: signal is true;
	signal WX6428: std_logic; attribute dont_touch of WX6428: signal is true;
	signal WX6429: std_logic; attribute dont_touch of WX6429: signal is true;
	signal WX6430: std_logic; attribute dont_touch of WX6430: signal is true;
	signal WX6431: std_logic; attribute dont_touch of WX6431: signal is true;
	signal WX6432: std_logic; attribute dont_touch of WX6432: signal is true;
	signal WX6433: std_logic; attribute dont_touch of WX6433: signal is true;
	signal WX6434: std_logic; attribute dont_touch of WX6434: signal is true;
	signal WX6435: std_logic; attribute dont_touch of WX6435: signal is true;
	signal WX6436: std_logic; attribute dont_touch of WX6436: signal is true;
	signal WX6438: std_logic; attribute dont_touch of WX6438: signal is true;
	signal WX6440: std_logic; attribute dont_touch of WX6440: signal is true;
	signal WX6442: std_logic; attribute dont_touch of WX6442: signal is true;
	signal WX6444: std_logic; attribute dont_touch of WX6444: signal is true;
	signal WX6446: std_logic; attribute dont_touch of WX6446: signal is true;
	signal WX6448: std_logic; attribute dont_touch of WX6448: signal is true;
	signal WX6450: std_logic; attribute dont_touch of WX6450: signal is true;
	signal WX6452: std_logic; attribute dont_touch of WX6452: signal is true;
	signal WX6454: std_logic; attribute dont_touch of WX6454: signal is true;
	signal WX6456: std_logic; attribute dont_touch of WX6456: signal is true;
	signal WX6458: std_logic; attribute dont_touch of WX6458: signal is true;
	signal WX6460: std_logic; attribute dont_touch of WX6460: signal is true;
	signal WX6462: std_logic; attribute dont_touch of WX6462: signal is true;
	signal WX6464: std_logic; attribute dont_touch of WX6464: signal is true;
	signal WX6466: std_logic; attribute dont_touch of WX6466: signal is true;
	signal WX6468: std_logic; attribute dont_touch of WX6468: signal is true;
	signal WX6470: std_logic; attribute dont_touch of WX6470: signal is true;
	signal WX6472: std_logic; attribute dont_touch of WX6472: signal is true;
	signal WX6474: std_logic; attribute dont_touch of WX6474: signal is true;
	signal WX6476: std_logic; attribute dont_touch of WX6476: signal is true;
	signal WX6478: std_logic; attribute dont_touch of WX6478: signal is true;
	signal WX6480: std_logic; attribute dont_touch of WX6480: signal is true;
	signal WX6482: std_logic; attribute dont_touch of WX6482: signal is true;
	signal WX6484: std_logic; attribute dont_touch of WX6484: signal is true;
	signal WX6486: std_logic; attribute dont_touch of WX6486: signal is true;
	signal WX6488: std_logic; attribute dont_touch of WX6488: signal is true;
	signal WX6490: std_logic; attribute dont_touch of WX6490: signal is true;
	signal WX6492: std_logic; attribute dont_touch of WX6492: signal is true;
	signal WX6494: std_logic; attribute dont_touch of WX6494: signal is true;
	signal WX6496: std_logic; attribute dont_touch of WX6496: signal is true;
	signal WX6498: std_logic; attribute dont_touch of WX6498: signal is true;
	signal WX6500: std_logic; attribute dont_touch of WX6500: signal is true;
	signal WX6501: std_logic; attribute dont_touch of WX6501: signal is true;
	signal WX6502: std_logic; attribute dont_touch of WX6502: signal is true;
	signal WX6503: std_logic; attribute dont_touch of WX6503: signal is true;
	signal WX6504: std_logic; attribute dont_touch of WX6504: signal is true;
	signal WX6505: std_logic; attribute dont_touch of WX6505: signal is true;
	signal WX6506: std_logic; attribute dont_touch of WX6506: signal is true;
	signal WX6507: std_logic; attribute dont_touch of WX6507: signal is true;
	signal WX6508: std_logic; attribute dont_touch of WX6508: signal is true;
	signal WX6509: std_logic; attribute dont_touch of WX6509: signal is true;
	signal WX6510: std_logic; attribute dont_touch of WX6510: signal is true;
	signal WX6511: std_logic; attribute dont_touch of WX6511: signal is true;
	signal WX6512: std_logic; attribute dont_touch of WX6512: signal is true;
	signal WX6513: std_logic; attribute dont_touch of WX6513: signal is true;
	signal WX6514: std_logic; attribute dont_touch of WX6514: signal is true;
	signal WX6515: std_logic; attribute dont_touch of WX6515: signal is true;
	signal WX6516: std_logic; attribute dont_touch of WX6516: signal is true;
	signal WX6517: std_logic; attribute dont_touch of WX6517: signal is true;
	signal WX6518: std_logic; attribute dont_touch of WX6518: signal is true;
	signal WX6519: std_logic; attribute dont_touch of WX6519: signal is true;
	signal WX6520: std_logic; attribute dont_touch of WX6520: signal is true;
	signal WX6521: std_logic; attribute dont_touch of WX6521: signal is true;
	signal WX6522: std_logic; attribute dont_touch of WX6522: signal is true;
	signal WX6523: std_logic; attribute dont_touch of WX6523: signal is true;
	signal WX6524: std_logic; attribute dont_touch of WX6524: signal is true;
	signal WX6525: std_logic; attribute dont_touch of WX6525: signal is true;
	signal WX6526: std_logic; attribute dont_touch of WX6526: signal is true;
	signal WX6527: std_logic; attribute dont_touch of WX6527: signal is true;
	signal WX6528: std_logic; attribute dont_touch of WX6528: signal is true;
	signal WX6529: std_logic; attribute dont_touch of WX6529: signal is true;
	signal WX6530: std_logic; attribute dont_touch of WX6530: signal is true;
	signal WX6531: std_logic; attribute dont_touch of WX6531: signal is true;
	signal WX6532: std_logic; attribute dont_touch of WX6532: signal is true;
	signal WX6533: std_logic; attribute dont_touch of WX6533: signal is true;
	signal WX6534: std_logic; attribute dont_touch of WX6534: signal is true;
	signal WX6535: std_logic; attribute dont_touch of WX6535: signal is true;
	signal WX6536: std_logic; attribute dont_touch of WX6536: signal is true;
	signal WX6537: std_logic; attribute dont_touch of WX6537: signal is true;
	signal WX6538: std_logic; attribute dont_touch of WX6538: signal is true;
	signal WX6539: std_logic; attribute dont_touch of WX6539: signal is true;
	signal WX6540: std_logic; attribute dont_touch of WX6540: signal is true;
	signal WX6541: std_logic; attribute dont_touch of WX6541: signal is true;
	signal WX6542: std_logic; attribute dont_touch of WX6542: signal is true;
	signal WX6543: std_logic; attribute dont_touch of WX6543: signal is true;
	signal WX6544: std_logic; attribute dont_touch of WX6544: signal is true;
	signal WX6545: std_logic; attribute dont_touch of WX6545: signal is true;
	signal WX6546: std_logic; attribute dont_touch of WX6546: signal is true;
	signal WX6547: std_logic; attribute dont_touch of WX6547: signal is true;
	signal WX6548: std_logic; attribute dont_touch of WX6548: signal is true;
	signal WX6549: std_logic; attribute dont_touch of WX6549: signal is true;
	signal WX6550: std_logic; attribute dont_touch of WX6550: signal is true;
	signal WX6551: std_logic; attribute dont_touch of WX6551: signal is true;
	signal WX6552: std_logic; attribute dont_touch of WX6552: signal is true;
	signal WX6553: std_logic; attribute dont_touch of WX6553: signal is true;
	signal WX6554: std_logic; attribute dont_touch of WX6554: signal is true;
	signal WX6555: std_logic; attribute dont_touch of WX6555: signal is true;
	signal WX6556: std_logic; attribute dont_touch of WX6556: signal is true;
	signal WX6557: std_logic; attribute dont_touch of WX6557: signal is true;
	signal WX6558: std_logic; attribute dont_touch of WX6558: signal is true;
	signal WX6559: std_logic; attribute dont_touch of WX6559: signal is true;
	signal WX6560: std_logic; attribute dont_touch of WX6560: signal is true;
	signal WX6561: std_logic; attribute dont_touch of WX6561: signal is true;
	signal WX6562: std_logic; attribute dont_touch of WX6562: signal is true;
	signal WX6563: std_logic; attribute dont_touch of WX6563: signal is true;
	signal WX6564: std_logic; attribute dont_touch of WX6564: signal is true;
	signal WX6565: std_logic; attribute dont_touch of WX6565: signal is true;
	signal WX6566: std_logic; attribute dont_touch of WX6566: signal is true;
	signal WX6567: std_logic; attribute dont_touch of WX6567: signal is true;
	signal WX6568: std_logic; attribute dont_touch of WX6568: signal is true;
	signal WX6569: std_logic; attribute dont_touch of WX6569: signal is true;
	signal WX6570: std_logic; attribute dont_touch of WX6570: signal is true;
	signal WX6571: std_logic; attribute dont_touch of WX6571: signal is true;
	signal WX6572: std_logic; attribute dont_touch of WX6572: signal is true;
	signal WX6573: std_logic; attribute dont_touch of WX6573: signal is true;
	signal WX6574: std_logic; attribute dont_touch of WX6574: signal is true;
	signal WX6575: std_logic; attribute dont_touch of WX6575: signal is true;
	signal WX6576: std_logic; attribute dont_touch of WX6576: signal is true;
	signal WX6577: std_logic; attribute dont_touch of WX6577: signal is true;
	signal WX6578: std_logic; attribute dont_touch of WX6578: signal is true;
	signal WX6579: std_logic; attribute dont_touch of WX6579: signal is true;
	signal WX6580: std_logic; attribute dont_touch of WX6580: signal is true;
	signal WX6581: std_logic; attribute dont_touch of WX6581: signal is true;
	signal WX6582: std_logic; attribute dont_touch of WX6582: signal is true;
	signal WX6583: std_logic; attribute dont_touch of WX6583: signal is true;
	signal WX6584: std_logic; attribute dont_touch of WX6584: signal is true;
	signal WX6585: std_logic; attribute dont_touch of WX6585: signal is true;
	signal WX6586: std_logic; attribute dont_touch of WX6586: signal is true;
	signal WX6587: std_logic; attribute dont_touch of WX6587: signal is true;
	signal WX6588: std_logic; attribute dont_touch of WX6588: signal is true;
	signal WX6589: std_logic; attribute dont_touch of WX6589: signal is true;
	signal WX6590: std_logic; attribute dont_touch of WX6590: signal is true;
	signal WX6591: std_logic; attribute dont_touch of WX6591: signal is true;
	signal WX6592: std_logic; attribute dont_touch of WX6592: signal is true;
	signal WX6593: std_logic; attribute dont_touch of WX6593: signal is true;
	signal WX6594: std_logic; attribute dont_touch of WX6594: signal is true;
	signal WX6595: std_logic; attribute dont_touch of WX6595: signal is true;
	signal WX6596: std_logic; attribute dont_touch of WX6596: signal is true;
	signal WX6597: std_logic; attribute dont_touch of WX6597: signal is true;
	signal WX6598: std_logic; attribute dont_touch of WX6598: signal is true;
	signal WX6599: std_logic; attribute dont_touch of WX6599: signal is true;
	signal WX6600: std_logic; attribute dont_touch of WX6600: signal is true;
	signal WX6601: std_logic; attribute dont_touch of WX6601: signal is true;
	signal WX6602: std_logic; attribute dont_touch of WX6602: signal is true;
	signal WX6603: std_logic; attribute dont_touch of WX6603: signal is true;
	signal WX6604: std_logic; attribute dont_touch of WX6604: signal is true;
	signal WX6605: std_logic; attribute dont_touch of WX6605: signal is true;
	signal WX6606: std_logic; attribute dont_touch of WX6606: signal is true;
	signal WX6607: std_logic; attribute dont_touch of WX6607: signal is true;
	signal WX6608: std_logic; attribute dont_touch of WX6608: signal is true;
	signal WX6609: std_logic; attribute dont_touch of WX6609: signal is true;
	signal WX6610: std_logic; attribute dont_touch of WX6610: signal is true;
	signal WX6611: std_logic; attribute dont_touch of WX6611: signal is true;
	signal WX6612: std_logic; attribute dont_touch of WX6612: signal is true;
	signal WX6613: std_logic; attribute dont_touch of WX6613: signal is true;
	signal WX6614: std_logic; attribute dont_touch of WX6614: signal is true;
	signal WX6615: std_logic; attribute dont_touch of WX6615: signal is true;
	signal WX6616: std_logic; attribute dont_touch of WX6616: signal is true;
	signal WX6617: std_logic; attribute dont_touch of WX6617: signal is true;
	signal WX6618: std_logic; attribute dont_touch of WX6618: signal is true;
	signal WX6619: std_logic; attribute dont_touch of WX6619: signal is true;
	signal WX6620: std_logic; attribute dont_touch of WX6620: signal is true;
	signal WX6621: std_logic; attribute dont_touch of WX6621: signal is true;
	signal WX6622: std_logic; attribute dont_touch of WX6622: signal is true;
	signal WX6623: std_logic; attribute dont_touch of WX6623: signal is true;
	signal WX6624: std_logic; attribute dont_touch of WX6624: signal is true;
	signal WX6625: std_logic; attribute dont_touch of WX6625: signal is true;
	signal WX6626: std_logic; attribute dont_touch of WX6626: signal is true;
	signal WX6627: std_logic; attribute dont_touch of WX6627: signal is true;
	signal WX6628: std_logic; attribute dont_touch of WX6628: signal is true;
	signal WX6629: std_logic; attribute dont_touch of WX6629: signal is true;
	signal WX6630: std_logic; attribute dont_touch of WX6630: signal is true;
	signal WX6631: std_logic; attribute dont_touch of WX6631: signal is true;
	signal WX6632: std_logic; attribute dont_touch of WX6632: signal is true;
	signal WX6633: std_logic; attribute dont_touch of WX6633: signal is true;
	signal WX6634: std_logic; attribute dont_touch of WX6634: signal is true;
	signal WX6635: std_logic; attribute dont_touch of WX6635: signal is true;
	signal WX6636: std_logic; attribute dont_touch of WX6636: signal is true;
	signal WX6637: std_logic; attribute dont_touch of WX6637: signal is true;
	signal WX6638: std_logic; attribute dont_touch of WX6638: signal is true;
	signal WX6639: std_logic; attribute dont_touch of WX6639: signal is true;
	signal WX6640: std_logic; attribute dont_touch of WX6640: signal is true;
	signal WX6641: std_logic; attribute dont_touch of WX6641: signal is true;
	signal WX6642: std_logic; attribute dont_touch of WX6642: signal is true;
	signal WX6643: std_logic; attribute dont_touch of WX6643: signal is true;
	signal WX6644: std_logic; attribute dont_touch of WX6644: signal is true;
	signal WX6645: std_logic; attribute dont_touch of WX6645: signal is true;
	signal WX6646: std_logic; attribute dont_touch of WX6646: signal is true;
	signal WX6647: std_logic; attribute dont_touch of WX6647: signal is true;
	signal WX6648: std_logic; attribute dont_touch of WX6648: signal is true;
	signal WX6649: std_logic; attribute dont_touch of WX6649: signal is true;
	signal WX6650: std_logic; attribute dont_touch of WX6650: signal is true;
	signal WX6651: std_logic; attribute dont_touch of WX6651: signal is true;
	signal WX6652: std_logic; attribute dont_touch of WX6652: signal is true;
	signal WX6653: std_logic; attribute dont_touch of WX6653: signal is true;
	signal WX6654: std_logic; attribute dont_touch of WX6654: signal is true;
	signal WX6655: std_logic; attribute dont_touch of WX6655: signal is true;
	signal WX6656: std_logic; attribute dont_touch of WX6656: signal is true;
	signal WX6657: std_logic; attribute dont_touch of WX6657: signal is true;
	signal WX6658: std_logic; attribute dont_touch of WX6658: signal is true;
	signal WX6659: std_logic; attribute dont_touch of WX6659: signal is true;
	signal WX6660: std_logic; attribute dont_touch of WX6660: signal is true;
	signal WX6661: std_logic; attribute dont_touch of WX6661: signal is true;
	signal WX6662: std_logic; attribute dont_touch of WX6662: signal is true;
	signal WX6663: std_logic; attribute dont_touch of WX6663: signal is true;
	signal WX6664: std_logic; attribute dont_touch of WX6664: signal is true;
	signal WX6665: std_logic; attribute dont_touch of WX6665: signal is true;
	signal WX6666: std_logic; attribute dont_touch of WX6666: signal is true;
	signal WX6667: std_logic; attribute dont_touch of WX6667: signal is true;
	signal WX6668: std_logic; attribute dont_touch of WX6668: signal is true;
	signal WX6669: std_logic; attribute dont_touch of WX6669: signal is true;
	signal WX6670: std_logic; attribute dont_touch of WX6670: signal is true;
	signal WX6671: std_logic; attribute dont_touch of WX6671: signal is true;
	signal WX6672: std_logic; attribute dont_touch of WX6672: signal is true;
	signal WX6673: std_logic; attribute dont_touch of WX6673: signal is true;
	signal WX6674: std_logic; attribute dont_touch of WX6674: signal is true;
	signal WX6675: std_logic; attribute dont_touch of WX6675: signal is true;
	signal WX6676: std_logic; attribute dont_touch of WX6676: signal is true;
	signal WX6677: std_logic; attribute dont_touch of WX6677: signal is true;
	signal WX6678: std_logic; attribute dont_touch of WX6678: signal is true;
	signal WX6679: std_logic; attribute dont_touch of WX6679: signal is true;
	signal WX6680: std_logic; attribute dont_touch of WX6680: signal is true;
	signal WX6681: std_logic; attribute dont_touch of WX6681: signal is true;
	signal WX6682: std_logic; attribute dont_touch of WX6682: signal is true;
	signal WX6683: std_logic; attribute dont_touch of WX6683: signal is true;
	signal WX6684: std_logic; attribute dont_touch of WX6684: signal is true;
	signal WX6685: std_logic; attribute dont_touch of WX6685: signal is true;
	signal WX6686: std_logic; attribute dont_touch of WX6686: signal is true;
	signal WX6687: std_logic; attribute dont_touch of WX6687: signal is true;
	signal WX6688: std_logic; attribute dont_touch of WX6688: signal is true;
	signal WX6689: std_logic; attribute dont_touch of WX6689: signal is true;
	signal WX6690: std_logic; attribute dont_touch of WX6690: signal is true;
	signal WX6691: std_logic; attribute dont_touch of WX6691: signal is true;
	signal WX6692: std_logic; attribute dont_touch of WX6692: signal is true;
	signal WX6693: std_logic; attribute dont_touch of WX6693: signal is true;
	signal WX6694: std_logic; attribute dont_touch of WX6694: signal is true;
	signal WX6695: std_logic; attribute dont_touch of WX6695: signal is true;
	signal WX6696: std_logic; attribute dont_touch of WX6696: signal is true;
	signal WX6697: std_logic; attribute dont_touch of WX6697: signal is true;
	signal WX6698: std_logic; attribute dont_touch of WX6698: signal is true;
	signal WX6699: std_logic; attribute dont_touch of WX6699: signal is true;
	signal WX6700: std_logic; attribute dont_touch of WX6700: signal is true;
	signal WX6701: std_logic; attribute dont_touch of WX6701: signal is true;
	signal WX6702: std_logic; attribute dont_touch of WX6702: signal is true;
	signal WX6703: std_logic; attribute dont_touch of WX6703: signal is true;
	signal WX6704: std_logic; attribute dont_touch of WX6704: signal is true;
	signal WX6705: std_logic; attribute dont_touch of WX6705: signal is true;
	signal WX6706: std_logic; attribute dont_touch of WX6706: signal is true;
	signal WX6707: std_logic; attribute dont_touch of WX6707: signal is true;
	signal WX6708: std_logic; attribute dont_touch of WX6708: signal is true;
	signal WX6709: std_logic; attribute dont_touch of WX6709: signal is true;
	signal WX6710: std_logic; attribute dont_touch of WX6710: signal is true;
	signal WX6711: std_logic; attribute dont_touch of WX6711: signal is true;
	signal WX6712: std_logic; attribute dont_touch of WX6712: signal is true;
	signal WX6713: std_logic; attribute dont_touch of WX6713: signal is true;
	signal WX6714: std_logic; attribute dont_touch of WX6714: signal is true;
	signal WX6715: std_logic; attribute dont_touch of WX6715: signal is true;
	signal WX6716: std_logic; attribute dont_touch of WX6716: signal is true;
	signal WX6717: std_logic; attribute dont_touch of WX6717: signal is true;
	signal WX6718: std_logic; attribute dont_touch of WX6718: signal is true;
	signal WX6719: std_logic; attribute dont_touch of WX6719: signal is true;
	signal WX6720: std_logic; attribute dont_touch of WX6720: signal is true;
	signal WX6721: std_logic; attribute dont_touch of WX6721: signal is true;
	signal WX6722: std_logic; attribute dont_touch of WX6722: signal is true;
	signal WX6723: std_logic; attribute dont_touch of WX6723: signal is true;
	signal WX6724: std_logic; attribute dont_touch of WX6724: signal is true;
	signal WX6725: std_logic; attribute dont_touch of WX6725: signal is true;
	signal WX6726: std_logic; attribute dont_touch of WX6726: signal is true;
	signal WX6727: std_logic; attribute dont_touch of WX6727: signal is true;
	signal WX6728: std_logic; attribute dont_touch of WX6728: signal is true;
	signal WX6729: std_logic; attribute dont_touch of WX6729: signal is true;
	signal WX6730: std_logic; attribute dont_touch of WX6730: signal is true;
	signal WX6731: std_logic; attribute dont_touch of WX6731: signal is true;
	signal WX6732: std_logic; attribute dont_touch of WX6732: signal is true;
	signal WX6733: std_logic; attribute dont_touch of WX6733: signal is true;
	signal WX6734: std_logic; attribute dont_touch of WX6734: signal is true;
	signal WX6735: std_logic; attribute dont_touch of WX6735: signal is true;
	signal WX6736: std_logic; attribute dont_touch of WX6736: signal is true;
	signal WX6737: std_logic; attribute dont_touch of WX6737: signal is true;
	signal WX6738: std_logic; attribute dont_touch of WX6738: signal is true;
	signal WX6739: std_logic; attribute dont_touch of WX6739: signal is true;
	signal WX6740: std_logic; attribute dont_touch of WX6740: signal is true;
	signal WX6741: std_logic; attribute dont_touch of WX6741: signal is true;
	signal WX6742: std_logic; attribute dont_touch of WX6742: signal is true;
	signal WX6743: std_logic; attribute dont_touch of WX6743: signal is true;
	signal WX6744: std_logic; attribute dont_touch of WX6744: signal is true;
	signal WX6745: std_logic; attribute dont_touch of WX6745: signal is true;
	signal WX6746: std_logic; attribute dont_touch of WX6746: signal is true;
	signal WX6747: std_logic; attribute dont_touch of WX6747: signal is true;
	signal WX6748: std_logic; attribute dont_touch of WX6748: signal is true;
	signal WX6749: std_logic; attribute dont_touch of WX6749: signal is true;
	signal WX6750: std_logic; attribute dont_touch of WX6750: signal is true;
	signal WX6751: std_logic; attribute dont_touch of WX6751: signal is true;
	signal WX6752: std_logic; attribute dont_touch of WX6752: signal is true;
	signal WX6753: std_logic; attribute dont_touch of WX6753: signal is true;
	signal WX6754: std_logic; attribute dont_touch of WX6754: signal is true;
	signal WX6755: std_logic; attribute dont_touch of WX6755: signal is true;
	signal WX6756: std_logic; attribute dont_touch of WX6756: signal is true;
	signal WX6757: std_logic; attribute dont_touch of WX6757: signal is true;
	signal WX6758: std_logic; attribute dont_touch of WX6758: signal is true;
	signal WX6759: std_logic; attribute dont_touch of WX6759: signal is true;
	signal WX6760: std_logic; attribute dont_touch of WX6760: signal is true;
	signal WX6761: std_logic; attribute dont_touch of WX6761: signal is true;
	signal WX6762: std_logic; attribute dont_touch of WX6762: signal is true;
	signal WX6763: std_logic; attribute dont_touch of WX6763: signal is true;
	signal WX6764: std_logic; attribute dont_touch of WX6764: signal is true;
	signal WX6765: std_logic; attribute dont_touch of WX6765: signal is true;
	signal WX6766: std_logic; attribute dont_touch of WX6766: signal is true;
	signal WX6767: std_logic; attribute dont_touch of WX6767: signal is true;
	signal WX6768: std_logic; attribute dont_touch of WX6768: signal is true;
	signal WX6769: std_logic; attribute dont_touch of WX6769: signal is true;
	signal WX6770: std_logic; attribute dont_touch of WX6770: signal is true;
	signal WX6771: std_logic; attribute dont_touch of WX6771: signal is true;
	signal WX6772: std_logic; attribute dont_touch of WX6772: signal is true;
	signal WX6773: std_logic; attribute dont_touch of WX6773: signal is true;
	signal WX6774: std_logic; attribute dont_touch of WX6774: signal is true;
	signal WX6775: std_logic; attribute dont_touch of WX6775: signal is true;
	signal WX6776: std_logic; attribute dont_touch of WX6776: signal is true;
	signal WX6777: std_logic; attribute dont_touch of WX6777: signal is true;
	signal WX6778: std_logic; attribute dont_touch of WX6778: signal is true;
	signal WX6779: std_logic; attribute dont_touch of WX6779: signal is true;
	signal WX6780: std_logic; attribute dont_touch of WX6780: signal is true;
	signal WX6781: std_logic; attribute dont_touch of WX6781: signal is true;
	signal WX6782: std_logic; attribute dont_touch of WX6782: signal is true;
	signal WX6783: std_logic; attribute dont_touch of WX6783: signal is true;
	signal WX6784: std_logic; attribute dont_touch of WX6784: signal is true;
	signal WX6785: std_logic; attribute dont_touch of WX6785: signal is true;
	signal WX6786: std_logic; attribute dont_touch of WX6786: signal is true;
	signal WX6787: std_logic; attribute dont_touch of WX6787: signal is true;
	signal WX6788: std_logic; attribute dont_touch of WX6788: signal is true;
	signal WX6789: std_logic; attribute dont_touch of WX6789: signal is true;
	signal WX6790: std_logic; attribute dont_touch of WX6790: signal is true;
	signal WX6791: std_logic; attribute dont_touch of WX6791: signal is true;
	signal WX6792: std_logic; attribute dont_touch of WX6792: signal is true;
	signal WX6793: std_logic; attribute dont_touch of WX6793: signal is true;
	signal WX6794: std_logic; attribute dont_touch of WX6794: signal is true;
	signal WX6795: std_logic; attribute dont_touch of WX6795: signal is true;
	signal WX6796: std_logic; attribute dont_touch of WX6796: signal is true;
	signal WX6797: std_logic; attribute dont_touch of WX6797: signal is true;
	signal WX6798: std_logic; attribute dont_touch of WX6798: signal is true;
	signal WX6799: std_logic; attribute dont_touch of WX6799: signal is true;
	signal WX6800: std_logic; attribute dont_touch of WX6800: signal is true;
	signal WX6801: std_logic; attribute dont_touch of WX6801: signal is true;
	signal WX6802: std_logic; attribute dont_touch of WX6802: signal is true;
	signal WX6803: std_logic; attribute dont_touch of WX6803: signal is true;
	signal WX6804: std_logic; attribute dont_touch of WX6804: signal is true;
	signal WX6805: std_logic; attribute dont_touch of WX6805: signal is true;
	signal WX6806: std_logic; attribute dont_touch of WX6806: signal is true;
	signal WX6807: std_logic; attribute dont_touch of WX6807: signal is true;
	signal WX6808: std_logic; attribute dont_touch of WX6808: signal is true;
	signal WX6809: std_logic; attribute dont_touch of WX6809: signal is true;
	signal WX6810: std_logic; attribute dont_touch of WX6810: signal is true;
	signal WX6811: std_logic; attribute dont_touch of WX6811: signal is true;
	signal WX6812: std_logic; attribute dont_touch of WX6812: signal is true;
	signal WX6813: std_logic; attribute dont_touch of WX6813: signal is true;
	signal WX6814: std_logic; attribute dont_touch of WX6814: signal is true;
	signal WX6815: std_logic; attribute dont_touch of WX6815: signal is true;
	signal WX6816: std_logic; attribute dont_touch of WX6816: signal is true;
	signal WX6817: std_logic; attribute dont_touch of WX6817: signal is true;
	signal WX6818: std_logic; attribute dont_touch of WX6818: signal is true;
	signal WX6819: std_logic; attribute dont_touch of WX6819: signal is true;
	signal WX6820: std_logic; attribute dont_touch of WX6820: signal is true;
	signal WX6821: std_logic; attribute dont_touch of WX6821: signal is true;
	signal WX6822: std_logic; attribute dont_touch of WX6822: signal is true;
	signal WX6823: std_logic; attribute dont_touch of WX6823: signal is true;
	signal WX6824: std_logic; attribute dont_touch of WX6824: signal is true;
	signal WX6825: std_logic; attribute dont_touch of WX6825: signal is true;
	signal WX6826: std_logic; attribute dont_touch of WX6826: signal is true;
	signal WX6827: std_logic; attribute dont_touch of WX6827: signal is true;
	signal WX6828: std_logic; attribute dont_touch of WX6828: signal is true;
	signal WX6829: std_logic; attribute dont_touch of WX6829: signal is true;
	signal WX6830: std_logic; attribute dont_touch of WX6830: signal is true;
	signal WX6831: std_logic; attribute dont_touch of WX6831: signal is true;
	signal WX6832: std_logic; attribute dont_touch of WX6832: signal is true;
	signal WX6833: std_logic; attribute dont_touch of WX6833: signal is true;
	signal WX6834: std_logic; attribute dont_touch of WX6834: signal is true;
	signal WX6835: std_logic; attribute dont_touch of WX6835: signal is true;
	signal WX6836: std_logic; attribute dont_touch of WX6836: signal is true;
	signal WX6837: std_logic; attribute dont_touch of WX6837: signal is true;
	signal WX6838: std_logic; attribute dont_touch of WX6838: signal is true;
	signal WX6839: std_logic; attribute dont_touch of WX6839: signal is true;
	signal WX6840: std_logic; attribute dont_touch of WX6840: signal is true;
	signal WX6841: std_logic; attribute dont_touch of WX6841: signal is true;
	signal WX6842: std_logic; attribute dont_touch of WX6842: signal is true;
	signal WX6843: std_logic; attribute dont_touch of WX6843: signal is true;
	signal WX6844: std_logic; attribute dont_touch of WX6844: signal is true;
	signal WX6845: std_logic; attribute dont_touch of WX6845: signal is true;
	signal WX6846: std_logic; attribute dont_touch of WX6846: signal is true;
	signal WX6847: std_logic; attribute dont_touch of WX6847: signal is true;
	signal WX6848: std_logic; attribute dont_touch of WX6848: signal is true;
	signal WX6849: std_logic; attribute dont_touch of WX6849: signal is true;
	signal WX6850: std_logic; attribute dont_touch of WX6850: signal is true;
	signal WX6851: std_logic; attribute dont_touch of WX6851: signal is true;
	signal WX6852: std_logic; attribute dont_touch of WX6852: signal is true;
	signal WX6853: std_logic; attribute dont_touch of WX6853: signal is true;
	signal WX6854: std_logic; attribute dont_touch of WX6854: signal is true;
	signal WX6855: std_logic; attribute dont_touch of WX6855: signal is true;
	signal WX6856: std_logic; attribute dont_touch of WX6856: signal is true;
	signal WX6857: std_logic; attribute dont_touch of WX6857: signal is true;
	signal WX6858: std_logic; attribute dont_touch of WX6858: signal is true;
	signal WX6859: std_logic; attribute dont_touch of WX6859: signal is true;
	signal WX6860: std_logic; attribute dont_touch of WX6860: signal is true;
	signal WX6861: std_logic; attribute dont_touch of WX6861: signal is true;
	signal WX6862: std_logic; attribute dont_touch of WX6862: signal is true;
	signal WX6863: std_logic; attribute dont_touch of WX6863: signal is true;
	signal WX6864: std_logic; attribute dont_touch of WX6864: signal is true;
	signal WX6865: std_logic; attribute dont_touch of WX6865: signal is true;
	signal WX6866: std_logic; attribute dont_touch of WX6866: signal is true;
	signal WX6867: std_logic; attribute dont_touch of WX6867: signal is true;
	signal WX6868: std_logic; attribute dont_touch of WX6868: signal is true;
	signal WX6869: std_logic; attribute dont_touch of WX6869: signal is true;
	signal WX6870: std_logic; attribute dont_touch of WX6870: signal is true;
	signal WX6871: std_logic; attribute dont_touch of WX6871: signal is true;
	signal WX6872: std_logic; attribute dont_touch of WX6872: signal is true;
	signal WX6873: std_logic; attribute dont_touch of WX6873: signal is true;
	signal WX6874: std_logic; attribute dont_touch of WX6874: signal is true;
	signal WX6875: std_logic; attribute dont_touch of WX6875: signal is true;
	signal WX6876: std_logic; attribute dont_touch of WX6876: signal is true;
	signal WX6877: std_logic; attribute dont_touch of WX6877: signal is true;
	signal WX6878: std_logic; attribute dont_touch of WX6878: signal is true;
	signal WX6879: std_logic; attribute dont_touch of WX6879: signal is true;
	signal WX6880: std_logic; attribute dont_touch of WX6880: signal is true;
	signal WX6881: std_logic; attribute dont_touch of WX6881: signal is true;
	signal WX6882: std_logic; attribute dont_touch of WX6882: signal is true;
	signal WX6883: std_logic; attribute dont_touch of WX6883: signal is true;
	signal WX6884: std_logic; attribute dont_touch of WX6884: signal is true;
	signal WX6885: std_logic; attribute dont_touch of WX6885: signal is true;
	signal WX6886: std_logic; attribute dont_touch of WX6886: signal is true;
	signal WX6887: std_logic; attribute dont_touch of WX6887: signal is true;
	signal WX6888: std_logic; attribute dont_touch of WX6888: signal is true;
	signal WX6889: std_logic; attribute dont_touch of WX6889: signal is true;
	signal WX6890: std_logic; attribute dont_touch of WX6890: signal is true;
	signal WX6891: std_logic; attribute dont_touch of WX6891: signal is true;
	signal WX6892: std_logic; attribute dont_touch of WX6892: signal is true;
	signal WX6893: std_logic; attribute dont_touch of WX6893: signal is true;
	signal WX6894: std_logic; attribute dont_touch of WX6894: signal is true;
	signal WX6895: std_logic; attribute dont_touch of WX6895: signal is true;
	signal WX6896: std_logic; attribute dont_touch of WX6896: signal is true;
	signal WX6897: std_logic; attribute dont_touch of WX6897: signal is true;
	signal WX6898: std_logic; attribute dont_touch of WX6898: signal is true;
	signal WX6899: std_logic; attribute dont_touch of WX6899: signal is true;
	signal WX6900: std_logic; attribute dont_touch of WX6900: signal is true;
	signal WX6901: std_logic; attribute dont_touch of WX6901: signal is true;
	signal WX6902: std_logic; attribute dont_touch of WX6902: signal is true;
	signal WX6903: std_logic; attribute dont_touch of WX6903: signal is true;
	signal WX6904: std_logic; attribute dont_touch of WX6904: signal is true;
	signal WX6905: std_logic; attribute dont_touch of WX6905: signal is true;
	signal WX6906: std_logic; attribute dont_touch of WX6906: signal is true;
	signal WX6907: std_logic; attribute dont_touch of WX6907: signal is true;
	signal WX6908: std_logic; attribute dont_touch of WX6908: signal is true;
	signal WX6909: std_logic; attribute dont_touch of WX6909: signal is true;
	signal WX6910: std_logic; attribute dont_touch of WX6910: signal is true;
	signal WX6911: std_logic; attribute dont_touch of WX6911: signal is true;
	signal WX6912: std_logic; attribute dont_touch of WX6912: signal is true;
	signal WX6913: std_logic; attribute dont_touch of WX6913: signal is true;
	signal WX6914: std_logic; attribute dont_touch of WX6914: signal is true;
	signal WX6915: std_logic; attribute dont_touch of WX6915: signal is true;
	signal WX6916: std_logic; attribute dont_touch of WX6916: signal is true;
	signal WX6917: std_logic; attribute dont_touch of WX6917: signal is true;
	signal WX6918: std_logic; attribute dont_touch of WX6918: signal is true;
	signal WX6919: std_logic; attribute dont_touch of WX6919: signal is true;
	signal WX6920: std_logic; attribute dont_touch of WX6920: signal is true;
	signal WX6921: std_logic; attribute dont_touch of WX6921: signal is true;
	signal WX6922: std_logic; attribute dont_touch of WX6922: signal is true;
	signal WX6923: std_logic; attribute dont_touch of WX6923: signal is true;
	signal WX6924: std_logic; attribute dont_touch of WX6924: signal is true;
	signal WX6925: std_logic; attribute dont_touch of WX6925: signal is true;
	signal WX6926: std_logic; attribute dont_touch of WX6926: signal is true;
	signal WX6927: std_logic; attribute dont_touch of WX6927: signal is true;
	signal WX6928: std_logic; attribute dont_touch of WX6928: signal is true;
	signal WX6929: std_logic; attribute dont_touch of WX6929: signal is true;
	signal WX6930: std_logic; attribute dont_touch of WX6930: signal is true;
	signal WX6931: std_logic; attribute dont_touch of WX6931: signal is true;
	signal WX6932: std_logic; attribute dont_touch of WX6932: signal is true;
	signal WX6933: std_logic; attribute dont_touch of WX6933: signal is true;
	signal WX6934: std_logic; attribute dont_touch of WX6934: signal is true;
	signal WX6935: std_logic; attribute dont_touch of WX6935: signal is true;
	signal WX6936: std_logic; attribute dont_touch of WX6936: signal is true;
	signal WX6937: std_logic; attribute dont_touch of WX6937: signal is true;
	signal WX6938: std_logic; attribute dont_touch of WX6938: signal is true;
	signal WX6939: std_logic; attribute dont_touch of WX6939: signal is true;
	signal WX6940: std_logic; attribute dont_touch of WX6940: signal is true;
	signal WX6941: std_logic; attribute dont_touch of WX6941: signal is true;
	signal WX6942: std_logic; attribute dont_touch of WX6942: signal is true;
	signal WX6943: std_logic; attribute dont_touch of WX6943: signal is true;
	signal WX6944: std_logic; attribute dont_touch of WX6944: signal is true;
	signal WX6945: std_logic; attribute dont_touch of WX6945: signal is true;
	signal WX6946: std_logic; attribute dont_touch of WX6946: signal is true;
	signal WX6947: std_logic; attribute dont_touch of WX6947: signal is true;
	signal WX6948: std_logic; attribute dont_touch of WX6948: signal is true;
	signal WX6949: std_logic; attribute dont_touch of WX6949: signal is true;
	signal WX6950: std_logic; attribute dont_touch of WX6950: signal is true;
	signal WX6951: std_logic; attribute dont_touch of WX6951: signal is true;
	signal WX6952: std_logic; attribute dont_touch of WX6952: signal is true;
	signal WX6953: std_logic; attribute dont_touch of WX6953: signal is true;
	signal WX6954: std_logic; attribute dont_touch of WX6954: signal is true;
	signal WX6955: std_logic; attribute dont_touch of WX6955: signal is true;
	signal WX6956: std_logic; attribute dont_touch of WX6956: signal is true;
	signal WX6957: std_logic; attribute dont_touch of WX6957: signal is true;
	signal WX6958: std_logic; attribute dont_touch of WX6958: signal is true;
	signal WX6959: std_logic; attribute dont_touch of WX6959: signal is true;
	signal WX6960: std_logic; attribute dont_touch of WX6960: signal is true;
	signal WX6961: std_logic; attribute dont_touch of WX6961: signal is true;
	signal WX6962: std_logic; attribute dont_touch of WX6962: signal is true;
	signal WX6963: std_logic; attribute dont_touch of WX6963: signal is true;
	signal WX6964: std_logic; attribute dont_touch of WX6964: signal is true;
	signal WX6965: std_logic; attribute dont_touch of WX6965: signal is true;
	signal WX6966: std_logic; attribute dont_touch of WX6966: signal is true;
	signal WX6967: std_logic; attribute dont_touch of WX6967: signal is true;
	signal WX6968: std_logic; attribute dont_touch of WX6968: signal is true;
	signal WX6969: std_logic; attribute dont_touch of WX6969: signal is true;
	signal WX6970: std_logic; attribute dont_touch of WX6970: signal is true;
	signal WX6971: std_logic; attribute dont_touch of WX6971: signal is true;
	signal WX6972: std_logic; attribute dont_touch of WX6972: signal is true;
	signal WX6973: std_logic; attribute dont_touch of WX6973: signal is true;
	signal WX6974: std_logic; attribute dont_touch of WX6974: signal is true;
	signal WX6975: std_logic; attribute dont_touch of WX6975: signal is true;
	signal WX6976: std_logic; attribute dont_touch of WX6976: signal is true;
	signal WX6977: std_logic; attribute dont_touch of WX6977: signal is true;
	signal WX6978: std_logic; attribute dont_touch of WX6978: signal is true;
	signal WX6979: std_logic; attribute dont_touch of WX6979: signal is true;
	signal WX6980: std_logic; attribute dont_touch of WX6980: signal is true;
	signal WX6981: std_logic; attribute dont_touch of WX6981: signal is true;
	signal WX6982: std_logic; attribute dont_touch of WX6982: signal is true;
	signal WX6983: std_logic; attribute dont_touch of WX6983: signal is true;
	signal WX6984: std_logic; attribute dont_touch of WX6984: signal is true;
	signal WX6985: std_logic; attribute dont_touch of WX6985: signal is true;
	signal WX6986: std_logic; attribute dont_touch of WX6986: signal is true;
	signal WX6987: std_logic; attribute dont_touch of WX6987: signal is true;
	signal WX6988: std_logic; attribute dont_touch of WX6988: signal is true;
	signal WX6989: std_logic; attribute dont_touch of WX6989: signal is true;
	signal WX6990: std_logic; attribute dont_touch of WX6990: signal is true;
	signal WX6991: std_logic; attribute dont_touch of WX6991: signal is true;
	signal WX6992: std_logic; attribute dont_touch of WX6992: signal is true;
	signal WX6993: std_logic; attribute dont_touch of WX6993: signal is true;
	signal WX6994: std_logic; attribute dont_touch of WX6994: signal is true;
	signal WX6995: std_logic; attribute dont_touch of WX6995: signal is true;
	signal WX6996: std_logic; attribute dont_touch of WX6996: signal is true;
	signal WX6997: std_logic; attribute dont_touch of WX6997: signal is true;
	signal WX6998: std_logic; attribute dont_touch of WX6998: signal is true;
	signal WX6999: std_logic; attribute dont_touch of WX6999: signal is true;
	signal WX7000: std_logic; attribute dont_touch of WX7000: signal is true;
	signal WX7001: std_logic; attribute dont_touch of WX7001: signal is true;
	signal WX7002: std_logic; attribute dont_touch of WX7002: signal is true;
	signal WX7003: std_logic; attribute dont_touch of WX7003: signal is true;
	signal WX7004: std_logic; attribute dont_touch of WX7004: signal is true;
	signal WX7005: std_logic; attribute dont_touch of WX7005: signal is true;
	signal WX7006: std_logic; attribute dont_touch of WX7006: signal is true;
	signal WX7007: std_logic; attribute dont_touch of WX7007: signal is true;
	signal WX7008: std_logic; attribute dont_touch of WX7008: signal is true;
	signal WX7009: std_logic; attribute dont_touch of WX7009: signal is true;
	signal WX7010: std_logic; attribute dont_touch of WX7010: signal is true;
	signal WX7011: std_logic; attribute dont_touch of WX7011: signal is true;
	signal WX7012: std_logic; attribute dont_touch of WX7012: signal is true;
	signal WX7013: std_logic; attribute dont_touch of WX7013: signal is true;
	signal WX7014: std_logic; attribute dont_touch of WX7014: signal is true;
	signal WX7015: std_logic; attribute dont_touch of WX7015: signal is true;
	signal WX7016: std_logic; attribute dont_touch of WX7016: signal is true;
	signal WX7017: std_logic; attribute dont_touch of WX7017: signal is true;
	signal WX7018: std_logic; attribute dont_touch of WX7018: signal is true;
	signal WX7019: std_logic; attribute dont_touch of WX7019: signal is true;
	signal WX7020: std_logic; attribute dont_touch of WX7020: signal is true;
	signal WX7021: std_logic; attribute dont_touch of WX7021: signal is true;
	signal WX7022: std_logic; attribute dont_touch of WX7022: signal is true;
	signal WX7023: std_logic; attribute dont_touch of WX7023: signal is true;
	signal WX7024: std_logic; attribute dont_touch of WX7024: signal is true;
	signal WX7025: std_logic; attribute dont_touch of WX7025: signal is true;
	signal WX7026: std_logic; attribute dont_touch of WX7026: signal is true;
	signal WX7027: std_logic; attribute dont_touch of WX7027: signal is true;
	signal WX7028: std_logic; attribute dont_touch of WX7028: signal is true;
	signal WX7029: std_logic; attribute dont_touch of WX7029: signal is true;
	signal WX7030: std_logic; attribute dont_touch of WX7030: signal is true;
	signal WX7031: std_logic; attribute dont_touch of WX7031: signal is true;
	signal WX7032: std_logic; attribute dont_touch of WX7032: signal is true;
	signal WX7033: std_logic; attribute dont_touch of WX7033: signal is true;
	signal WX7034: std_logic; attribute dont_touch of WX7034: signal is true;
	signal WX7035: std_logic; attribute dont_touch of WX7035: signal is true;
	signal WX7036: std_logic; attribute dont_touch of WX7036: signal is true;
	signal WX7037: std_logic; attribute dont_touch of WX7037: signal is true;
	signal WX7038: std_logic; attribute dont_touch of WX7038: signal is true;
	signal WX7039: std_logic; attribute dont_touch of WX7039: signal is true;
	signal WX7040: std_logic; attribute dont_touch of WX7040: signal is true;
	signal WX7041: std_logic; attribute dont_touch of WX7041: signal is true;
	signal WX7042: std_logic; attribute dont_touch of WX7042: signal is true;
	signal WX7043: std_logic; attribute dont_touch of WX7043: signal is true;
	signal WX7044: std_logic; attribute dont_touch of WX7044: signal is true;
	signal WX7045: std_logic; attribute dont_touch of WX7045: signal is true;
	signal WX7046: std_logic; attribute dont_touch of WX7046: signal is true;
	signal WX7047: std_logic; attribute dont_touch of WX7047: signal is true;
	signal WX7048: std_logic; attribute dont_touch of WX7048: signal is true;
	signal WX7049: std_logic; attribute dont_touch of WX7049: signal is true;
	signal WX7050: std_logic; attribute dont_touch of WX7050: signal is true;
	signal WX7051: std_logic; attribute dont_touch of WX7051: signal is true;
	signal WX7052: std_logic; attribute dont_touch of WX7052: signal is true;
	signal WX7053: std_logic; attribute dont_touch of WX7053: signal is true;
	signal WX7054: std_logic; attribute dont_touch of WX7054: signal is true;
	signal WX7055: std_logic; attribute dont_touch of WX7055: signal is true;
	signal WX7056: std_logic; attribute dont_touch of WX7056: signal is true;
	signal WX7057: std_logic; attribute dont_touch of WX7057: signal is true;
	signal WX7058: std_logic; attribute dont_touch of WX7058: signal is true;
	signal WX7059: std_logic; attribute dont_touch of WX7059: signal is true;
	signal WX7060: std_logic; attribute dont_touch of WX7060: signal is true;
	signal WX7061: std_logic; attribute dont_touch of WX7061: signal is true;
	signal WX7062: std_logic; attribute dont_touch of WX7062: signal is true;
	signal WX7063: std_logic; attribute dont_touch of WX7063: signal is true;
	signal WX7064: std_logic; attribute dont_touch of WX7064: signal is true;
	signal WX7065: std_logic; attribute dont_touch of WX7065: signal is true;
	signal WX7066: std_logic; attribute dont_touch of WX7066: signal is true;
	signal WX7067: std_logic; attribute dont_touch of WX7067: signal is true;
	signal WX7068: std_logic; attribute dont_touch of WX7068: signal is true;
	signal WX7069: std_logic; attribute dont_touch of WX7069: signal is true;
	signal WX7070: std_logic; attribute dont_touch of WX7070: signal is true;
	signal WX7071: std_logic; attribute dont_touch of WX7071: signal is true;
	signal WX7072: std_logic; attribute dont_touch of WX7072: signal is true;
	signal WX7073: std_logic; attribute dont_touch of WX7073: signal is true;
	signal WX7074: std_logic; attribute dont_touch of WX7074: signal is true;
	signal WX7075: std_logic; attribute dont_touch of WX7075: signal is true;
	signal WX7076: std_logic; attribute dont_touch of WX7076: signal is true;
	signal WX7077: std_logic; attribute dont_touch of WX7077: signal is true;
	signal WX7078: std_logic; attribute dont_touch of WX7078: signal is true;
	signal WX7079: std_logic; attribute dont_touch of WX7079: signal is true;
	signal WX7080: std_logic; attribute dont_touch of WX7080: signal is true;
	signal WX7081: std_logic; attribute dont_touch of WX7081: signal is true;
	signal WX7082: std_logic; attribute dont_touch of WX7082: signal is true;
	signal WX7083: std_logic; attribute dont_touch of WX7083: signal is true;
	signal WX7084: std_logic; attribute dont_touch of WX7084: signal is true;
	signal WX7085: std_logic; attribute dont_touch of WX7085: signal is true;
	signal WX7086: std_logic; attribute dont_touch of WX7086: signal is true;
	signal WX7087: std_logic; attribute dont_touch of WX7087: signal is true;
	signal WX7088: std_logic; attribute dont_touch of WX7088: signal is true;
	signal WX7089: std_logic; attribute dont_touch of WX7089: signal is true;
	signal WX7090: std_logic; attribute dont_touch of WX7090: signal is true;
	signal WX7091: std_logic; attribute dont_touch of WX7091: signal is true;
	signal WX7092: std_logic; attribute dont_touch of WX7092: signal is true;
	signal WX7093: std_logic; attribute dont_touch of WX7093: signal is true;
	signal WX7094: std_logic; attribute dont_touch of WX7094: signal is true;
	signal WX7095: std_logic; attribute dont_touch of WX7095: signal is true;
	signal WX7096: std_logic; attribute dont_touch of WX7096: signal is true;
	signal WX7097: std_logic; attribute dont_touch of WX7097: signal is true;
	signal WX7098: std_logic; attribute dont_touch of WX7098: signal is true;
	signal WX7099: std_logic; attribute dont_touch of WX7099: signal is true;
	signal WX7100: std_logic; attribute dont_touch of WX7100: signal is true;
	signal WX7101: std_logic; attribute dont_touch of WX7101: signal is true;
	signal WX7102: std_logic; attribute dont_touch of WX7102: signal is true;
	signal WX7103: std_logic; attribute dont_touch of WX7103: signal is true;
	signal WX7104: std_logic; attribute dont_touch of WX7104: signal is true;
	signal WX7105: std_logic; attribute dont_touch of WX7105: signal is true;
	signal WX7106: std_logic; attribute dont_touch of WX7106: signal is true;
	signal WX7107: std_logic; attribute dont_touch of WX7107: signal is true;
	signal WX7108: std_logic; attribute dont_touch of WX7108: signal is true;
	signal WX7109: std_logic; attribute dont_touch of WX7109: signal is true;
	signal WX7110: std_logic; attribute dont_touch of WX7110: signal is true;
	signal WX7111: std_logic; attribute dont_touch of WX7111: signal is true;
	signal WX7112: std_logic; attribute dont_touch of WX7112: signal is true;
	signal WX7113: std_logic; attribute dont_touch of WX7113: signal is true;
	signal WX7114: std_logic; attribute dont_touch of WX7114: signal is true;
	signal WX7115: std_logic; attribute dont_touch of WX7115: signal is true;
	signal WX7116: std_logic; attribute dont_touch of WX7116: signal is true;
	signal WX7117: std_logic; attribute dont_touch of WX7117: signal is true;
	signal WX7118: std_logic; attribute dont_touch of WX7118: signal is true;
	signal WX7119: std_logic; attribute dont_touch of WX7119: signal is true;
	signal WX7120: std_logic; attribute dont_touch of WX7120: signal is true;
	signal WX7121: std_logic; attribute dont_touch of WX7121: signal is true;
	signal WX7122: std_logic; attribute dont_touch of WX7122: signal is true;
	signal WX7123: std_logic; attribute dont_touch of WX7123: signal is true;
	signal WX7124: std_logic; attribute dont_touch of WX7124: signal is true;
	signal WX7125: std_logic; attribute dont_touch of WX7125: signal is true;
	signal WX7126: std_logic; attribute dont_touch of WX7126: signal is true;
	signal WX7127: std_logic; attribute dont_touch of WX7127: signal is true;
	signal WX7128: std_logic; attribute dont_touch of WX7128: signal is true;
	signal WX7129: std_logic; attribute dont_touch of WX7129: signal is true;
	signal WX7130: std_logic; attribute dont_touch of WX7130: signal is true;
	signal WX7131: std_logic; attribute dont_touch of WX7131: signal is true;
	signal WX7132: std_logic; attribute dont_touch of WX7132: signal is true;
	signal WX7133: std_logic; attribute dont_touch of WX7133: signal is true;
	signal WX7134: std_logic; attribute dont_touch of WX7134: signal is true;
	signal WX7135: std_logic; attribute dont_touch of WX7135: signal is true;
	signal WX7136: std_logic; attribute dont_touch of WX7136: signal is true;
	signal WX7137: std_logic; attribute dont_touch of WX7137: signal is true;
	signal WX7138: std_logic; attribute dont_touch of WX7138: signal is true;
	signal WX7139: std_logic; attribute dont_touch of WX7139: signal is true;
	signal WX7140: std_logic; attribute dont_touch of WX7140: signal is true;
	signal WX7141: std_logic; attribute dont_touch of WX7141: signal is true;
	signal WX7142: std_logic; attribute dont_touch of WX7142: signal is true;
	signal WX7143: std_logic; attribute dont_touch of WX7143: signal is true;
	signal WX7144: std_logic; attribute dont_touch of WX7144: signal is true;
	signal WX7145: std_logic; attribute dont_touch of WX7145: signal is true;
	signal WX7146: std_logic; attribute dont_touch of WX7146: signal is true;
	signal WX7147: std_logic; attribute dont_touch of WX7147: signal is true;
	signal WX7148: std_logic; attribute dont_touch of WX7148: signal is true;
	signal WX7149: std_logic; attribute dont_touch of WX7149: signal is true;
	signal WX7150: std_logic; attribute dont_touch of WX7150: signal is true;
	signal WX7151: std_logic; attribute dont_touch of WX7151: signal is true;
	signal WX7152: std_logic; attribute dont_touch of WX7152: signal is true;
	signal WX7153: std_logic; attribute dont_touch of WX7153: signal is true;
	signal WX7154: std_logic; attribute dont_touch of WX7154: signal is true;
	signal WX7155: std_logic; attribute dont_touch of WX7155: signal is true;
	signal WX7156: std_logic; attribute dont_touch of WX7156: signal is true;
	signal WX7157: std_logic; attribute dont_touch of WX7157: signal is true;
	signal WX7158: std_logic; attribute dont_touch of WX7158: signal is true;
	signal WX7159: std_logic; attribute dont_touch of WX7159: signal is true;
	signal WX7160: std_logic; attribute dont_touch of WX7160: signal is true;
	signal WX7161: std_logic; attribute dont_touch of WX7161: signal is true;
	signal WX7162: std_logic; attribute dont_touch of WX7162: signal is true;
	signal WX7163: std_logic; attribute dont_touch of WX7163: signal is true;
	signal WX7164: std_logic; attribute dont_touch of WX7164: signal is true;
	signal WX7165: std_logic; attribute dont_touch of WX7165: signal is true;
	signal WX7166: std_logic; attribute dont_touch of WX7166: signal is true;
	signal WX7167: std_logic; attribute dont_touch of WX7167: signal is true;
	signal WX7168: std_logic; attribute dont_touch of WX7168: signal is true;
	signal WX7169: std_logic; attribute dont_touch of WX7169: signal is true;
	signal WX7170: std_logic; attribute dont_touch of WX7170: signal is true;
	signal WX7171: std_logic; attribute dont_touch of WX7171: signal is true;
	signal WX7172: std_logic; attribute dont_touch of WX7172: signal is true;
	signal WX7173: std_logic; attribute dont_touch of WX7173: signal is true;
	signal WX7174: std_logic; attribute dont_touch of WX7174: signal is true;
	signal WX7175: std_logic; attribute dont_touch of WX7175: signal is true;
	signal WX7176: std_logic; attribute dont_touch of WX7176: signal is true;
	signal WX7177: std_logic; attribute dont_touch of WX7177: signal is true;
	signal WX7178: std_logic; attribute dont_touch of WX7178: signal is true;
	signal WX7179: std_logic; attribute dont_touch of WX7179: signal is true;
	signal WX7180: std_logic; attribute dont_touch of WX7180: signal is true;
	signal WX7181: std_logic; attribute dont_touch of WX7181: signal is true;
	signal WX7182: std_logic; attribute dont_touch of WX7182: signal is true;
	signal WX7183: std_logic; attribute dont_touch of WX7183: signal is true;
	signal WX7184: std_logic; attribute dont_touch of WX7184: signal is true;
	signal WX7185: std_logic; attribute dont_touch of WX7185: signal is true;
	signal WX7186: std_logic; attribute dont_touch of WX7186: signal is true;
	signal WX7187: std_logic; attribute dont_touch of WX7187: signal is true;
	signal WX7188: std_logic; attribute dont_touch of WX7188: signal is true;
	signal WX7189: std_logic; attribute dont_touch of WX7189: signal is true;
	signal WX7190: std_logic; attribute dont_touch of WX7190: signal is true;
	signal WX7191: std_logic; attribute dont_touch of WX7191: signal is true;
	signal WX7192: std_logic; attribute dont_touch of WX7192: signal is true;
	signal WX7193: std_logic; attribute dont_touch of WX7193: signal is true;
	signal WX7194: std_logic; attribute dont_touch of WX7194: signal is true;
	signal WX7195: std_logic; attribute dont_touch of WX7195: signal is true;
	signal WX7196: std_logic; attribute dont_touch of WX7196: signal is true;
	signal WX7197: std_logic; attribute dont_touch of WX7197: signal is true;
	signal WX7198: std_logic; attribute dont_touch of WX7198: signal is true;
	signal WX7199: std_logic; attribute dont_touch of WX7199: signal is true;
	signal WX7200: std_logic; attribute dont_touch of WX7200: signal is true;
	signal WX7201: std_logic; attribute dont_touch of WX7201: signal is true;
	signal WX7202: std_logic; attribute dont_touch of WX7202: signal is true;
	signal WX7203: std_logic; attribute dont_touch of WX7203: signal is true;
	signal WX7204: std_logic; attribute dont_touch of WX7204: signal is true;
	signal WX7205: std_logic; attribute dont_touch of WX7205: signal is true;
	signal WX7206: std_logic; attribute dont_touch of WX7206: signal is true;
	signal WX7207: std_logic; attribute dont_touch of WX7207: signal is true;
	signal WX7208: std_logic; attribute dont_touch of WX7208: signal is true;
	signal WX7209: std_logic; attribute dont_touch of WX7209: signal is true;
	signal WX7210: std_logic; attribute dont_touch of WX7210: signal is true;
	signal WX7211: std_logic; attribute dont_touch of WX7211: signal is true;
	signal WX7212: std_logic; attribute dont_touch of WX7212: signal is true;
	signal WX7213: std_logic; attribute dont_touch of WX7213: signal is true;
	signal WX7214: std_logic; attribute dont_touch of WX7214: signal is true;
	signal WX7215: std_logic; attribute dont_touch of WX7215: signal is true;
	signal WX7216: std_logic; attribute dont_touch of WX7216: signal is true;
	signal WX7217: std_logic; attribute dont_touch of WX7217: signal is true;
	signal WX7218: std_logic; attribute dont_touch of WX7218: signal is true;
	signal WX7219: std_logic; attribute dont_touch of WX7219: signal is true;
	signal WX7220: std_logic; attribute dont_touch of WX7220: signal is true;
	signal WX7221: std_logic; attribute dont_touch of WX7221: signal is true;
	signal WX7222: std_logic; attribute dont_touch of WX7222: signal is true;
	signal WX7223: std_logic; attribute dont_touch of WX7223: signal is true;
	signal WX7224: std_logic; attribute dont_touch of WX7224: signal is true;
	signal WX7225: std_logic; attribute dont_touch of WX7225: signal is true;
	signal WX7226: std_logic; attribute dont_touch of WX7226: signal is true;
	signal WX7227: std_logic; attribute dont_touch of WX7227: signal is true;
	signal WX7228: std_logic; attribute dont_touch of WX7228: signal is true;
	signal WX7229: std_logic; attribute dont_touch of WX7229: signal is true;
	signal WX7230: std_logic; attribute dont_touch of WX7230: signal is true;
	signal WX7231: std_logic; attribute dont_touch of WX7231: signal is true;
	signal WX7232: std_logic; attribute dont_touch of WX7232: signal is true;
	signal WX7233: std_logic; attribute dont_touch of WX7233: signal is true;
	signal WX7234: std_logic; attribute dont_touch of WX7234: signal is true;
	signal WX7235: std_logic; attribute dont_touch of WX7235: signal is true;
	signal WX7236: std_logic; attribute dont_touch of WX7236: signal is true;
	signal WX7237: std_logic; attribute dont_touch of WX7237: signal is true;
	signal WX7238: std_logic; attribute dont_touch of WX7238: signal is true;
	signal WX7239: std_logic; attribute dont_touch of WX7239: signal is true;
	signal WX7240: std_logic; attribute dont_touch of WX7240: signal is true;
	signal WX7241: std_logic; attribute dont_touch of WX7241: signal is true;
	signal WX7242: std_logic; attribute dont_touch of WX7242: signal is true;
	signal WX7243: std_logic; attribute dont_touch of WX7243: signal is true;
	signal WX7244: std_logic; attribute dont_touch of WX7244: signal is true;
	signal WX7245: std_logic; attribute dont_touch of WX7245: signal is true;
	signal WX7246: std_logic; attribute dont_touch of WX7246: signal is true;
	signal WX7247: std_logic; attribute dont_touch of WX7247: signal is true;
	signal WX7248: std_logic; attribute dont_touch of WX7248: signal is true;
	signal WX7249: std_logic; attribute dont_touch of WX7249: signal is true;
	signal WX7250: std_logic; attribute dont_touch of WX7250: signal is true;
	signal WX7251: std_logic; attribute dont_touch of WX7251: signal is true;
	signal WX7252: std_logic; attribute dont_touch of WX7252: signal is true;
	signal WX7253: std_logic; attribute dont_touch of WX7253: signal is true;
	signal WX7254: std_logic; attribute dont_touch of WX7254: signal is true;
	signal WX7255: std_logic; attribute dont_touch of WX7255: signal is true;
	signal WX7256: std_logic; attribute dont_touch of WX7256: signal is true;
	signal WX7257: std_logic; attribute dont_touch of WX7257: signal is true;
	signal WX7258: std_logic; attribute dont_touch of WX7258: signal is true;
	signal WX7259: std_logic; attribute dont_touch of WX7259: signal is true;
	signal WX7260: std_logic; attribute dont_touch of WX7260: signal is true;
	signal WX7261: std_logic; attribute dont_touch of WX7261: signal is true;
	signal WX7262: std_logic; attribute dont_touch of WX7262: signal is true;
	signal WX7263: std_logic; attribute dont_touch of WX7263: signal is true;
	signal WX7264: std_logic; attribute dont_touch of WX7264: signal is true;
	signal WX7265: std_logic; attribute dont_touch of WX7265: signal is true;
	signal WX7266: std_logic; attribute dont_touch of WX7266: signal is true;
	signal WX7267: std_logic; attribute dont_touch of WX7267: signal is true;
	signal WX7268: std_logic; attribute dont_touch of WX7268: signal is true;
	signal WX7269: std_logic; attribute dont_touch of WX7269: signal is true;
	signal WX7270: std_logic; attribute dont_touch of WX7270: signal is true;
	signal WX7271: std_logic; attribute dont_touch of WX7271: signal is true;
	signal WX7272: std_logic; attribute dont_touch of WX7272: signal is true;
	signal WX7273: std_logic; attribute dont_touch of WX7273: signal is true;
	signal WX7274: std_logic; attribute dont_touch of WX7274: signal is true;
	signal WX7275: std_logic; attribute dont_touch of WX7275: signal is true;
	signal WX7276: std_logic; attribute dont_touch of WX7276: signal is true;
	signal WX7277: std_logic; attribute dont_touch of WX7277: signal is true;
	signal WX7278: std_logic; attribute dont_touch of WX7278: signal is true;
	signal WX7279: std_logic; attribute dont_touch of WX7279: signal is true;
	signal WX7280: std_logic; attribute dont_touch of WX7280: signal is true;
	signal WX7281: std_logic; attribute dont_touch of WX7281: signal is true;
	signal WX7282: std_logic; attribute dont_touch of WX7282: signal is true;
	signal WX7283: std_logic; attribute dont_touch of WX7283: signal is true;
	signal WX7284: std_logic; attribute dont_touch of WX7284: signal is true;
	signal WX7285: std_logic; attribute dont_touch of WX7285: signal is true;
	signal WX7286: std_logic; attribute dont_touch of WX7286: signal is true;
	signal WX7287: std_logic; attribute dont_touch of WX7287: signal is true;
	signal WX7288: std_logic; attribute dont_touch of WX7288: signal is true;
	signal WX7289: std_logic; attribute dont_touch of WX7289: signal is true;
	signal WX7290: std_logic; attribute dont_touch of WX7290: signal is true;
	signal WX7291: std_logic; attribute dont_touch of WX7291: signal is true;
	signal WX7292: std_logic; attribute dont_touch of WX7292: signal is true;
	signal WX7293: std_logic; attribute dont_touch of WX7293: signal is true;
	signal WX7294: std_logic; attribute dont_touch of WX7294: signal is true;
	signal WX7295: std_logic; attribute dont_touch of WX7295: signal is true;
	signal WX7296: std_logic; attribute dont_touch of WX7296: signal is true;
	signal WX7297: std_logic; attribute dont_touch of WX7297: signal is true;
	signal WX7298: std_logic; attribute dont_touch of WX7298: signal is true;
	signal WX7299: std_logic; attribute dont_touch of WX7299: signal is true;
	signal WX7300: std_logic; attribute dont_touch of WX7300: signal is true;
	signal WX7301: std_logic; attribute dont_touch of WX7301: signal is true;
	signal WX7302: std_logic; attribute dont_touch of WX7302: signal is true;
	signal WX7303: std_logic; attribute dont_touch of WX7303: signal is true;
	signal WX7304: std_logic; attribute dont_touch of WX7304: signal is true;
	signal WX7305: std_logic; attribute dont_touch of WX7305: signal is true;
	signal WX7306: std_logic; attribute dont_touch of WX7306: signal is true;
	signal WX7307: std_logic; attribute dont_touch of WX7307: signal is true;
	signal WX7308: std_logic; attribute dont_touch of WX7308: signal is true;
	signal WX7309: std_logic; attribute dont_touch of WX7309: signal is true;
	signal WX7310: std_logic; attribute dont_touch of WX7310: signal is true;
	signal WX7311: std_logic; attribute dont_touch of WX7311: signal is true;
	signal WX7312: std_logic; attribute dont_touch of WX7312: signal is true;
	signal WX7313: std_logic; attribute dont_touch of WX7313: signal is true;
	signal WX7314: std_logic; attribute dont_touch of WX7314: signal is true;
	signal WX7315: std_logic; attribute dont_touch of WX7315: signal is true;
	signal WX7316: std_logic; attribute dont_touch of WX7316: signal is true;
	signal WX7317: std_logic; attribute dont_touch of WX7317: signal is true;
	signal WX7318: std_logic; attribute dont_touch of WX7318: signal is true;
	signal WX7319: std_logic; attribute dont_touch of WX7319: signal is true;
	signal WX7320: std_logic; attribute dont_touch of WX7320: signal is true;
	signal WX7321: std_logic; attribute dont_touch of WX7321: signal is true;
	signal WX7322: std_logic; attribute dont_touch of WX7322: signal is true;
	signal WX7323: std_logic; attribute dont_touch of WX7323: signal is true;
	signal WX7324: std_logic; attribute dont_touch of WX7324: signal is true;
	signal WX7325: std_logic; attribute dont_touch of WX7325: signal is true;
	signal WX7326: std_logic; attribute dont_touch of WX7326: signal is true;
	signal WX7327: std_logic; attribute dont_touch of WX7327: signal is true;
	signal WX7328: std_logic; attribute dont_touch of WX7328: signal is true;
	signal WX7329: std_logic; attribute dont_touch of WX7329: signal is true;
	signal WX7330: std_logic; attribute dont_touch of WX7330: signal is true;
	signal WX7331: std_logic; attribute dont_touch of WX7331: signal is true;
	signal WX7332: std_logic; attribute dont_touch of WX7332: signal is true;
	signal WX7333: std_logic; attribute dont_touch of WX7333: signal is true;
	signal WX7334: std_logic; attribute dont_touch of WX7334: signal is true;
	signal WX7335: std_logic; attribute dont_touch of WX7335: signal is true;
	signal WX7336: std_logic; attribute dont_touch of WX7336: signal is true;
	signal WX7337: std_logic; attribute dont_touch of WX7337: signal is true;
	signal WX7338: std_logic; attribute dont_touch of WX7338: signal is true;
	signal WX7339: std_logic; attribute dont_touch of WX7339: signal is true;
	signal WX7340: std_logic; attribute dont_touch of WX7340: signal is true;
	signal WX7341: std_logic; attribute dont_touch of WX7341: signal is true;
	signal WX7342: std_logic; attribute dont_touch of WX7342: signal is true;
	signal WX7343: std_logic; attribute dont_touch of WX7343: signal is true;
	signal WX7344: std_logic; attribute dont_touch of WX7344: signal is true;
	signal WX7345: std_logic; attribute dont_touch of WX7345: signal is true;
	signal WX7346: std_logic; attribute dont_touch of WX7346: signal is true;
	signal WX7347: std_logic; attribute dont_touch of WX7347: signal is true;
	signal WX7348: std_logic; attribute dont_touch of WX7348: signal is true;
	signal WX7349: std_logic; attribute dont_touch of WX7349: signal is true;
	signal WX7350: std_logic; attribute dont_touch of WX7350: signal is true;
	signal WX7351: std_logic; attribute dont_touch of WX7351: signal is true;
	signal WX7352: std_logic; attribute dont_touch of WX7352: signal is true;
	signal WX7353: std_logic; attribute dont_touch of WX7353: signal is true;
	signal WX7354: std_logic; attribute dont_touch of WX7354: signal is true;
	signal WX7355: std_logic; attribute dont_touch of WX7355: signal is true;
	signal WX7356: std_logic; attribute dont_touch of WX7356: signal is true;
	signal WX7357: std_logic; attribute dont_touch of WX7357: signal is true;
	signal WX7358: std_logic; attribute dont_touch of WX7358: signal is true;
	signal WX7359: std_logic; attribute dont_touch of WX7359: signal is true;
	signal WX7360: std_logic; attribute dont_touch of WX7360: signal is true;
	signal WX7361: std_logic; attribute dont_touch of WX7361: signal is true;
	signal WX7362: std_logic; attribute dont_touch of WX7362: signal is true;
	signal WX7363: std_logic; attribute dont_touch of WX7363: signal is true;
	signal WX7364: std_logic; attribute dont_touch of WX7364: signal is true;
	signal WX7365: std_logic; attribute dont_touch of WX7365: signal is true;
	signal WX7366: std_logic; attribute dont_touch of WX7366: signal is true;
	signal WX7367: std_logic; attribute dont_touch of WX7367: signal is true;
	signal WX7368: std_logic; attribute dont_touch of WX7368: signal is true;
	signal WX7369: std_logic; attribute dont_touch of WX7369: signal is true;
	signal WX7370: std_logic; attribute dont_touch of WX7370: signal is true;
	signal WX7371: std_logic; attribute dont_touch of WX7371: signal is true;
	signal WX7372: std_logic; attribute dont_touch of WX7372: signal is true;
	signal WX7373: std_logic; attribute dont_touch of WX7373: signal is true;
	signal WX7374: std_logic; attribute dont_touch of WX7374: signal is true;
	signal WX7375: std_logic; attribute dont_touch of WX7375: signal is true;
	signal WX7376: std_logic; attribute dont_touch of WX7376: signal is true;
	signal WX7377: std_logic; attribute dont_touch of WX7377: signal is true;
	signal WX7378: std_logic; attribute dont_touch of WX7378: signal is true;
	signal WX7379: std_logic; attribute dont_touch of WX7379: signal is true;
	signal WX7380: std_logic; attribute dont_touch of WX7380: signal is true;
	signal WX7381: std_logic; attribute dont_touch of WX7381: signal is true;
	signal WX7382: std_logic; attribute dont_touch of WX7382: signal is true;
	signal WX7383: std_logic; attribute dont_touch of WX7383: signal is true;
	signal WX7384: std_logic; attribute dont_touch of WX7384: signal is true;
	signal WX7385: std_logic; attribute dont_touch of WX7385: signal is true;
	signal WX7386: std_logic; attribute dont_touch of WX7386: signal is true;
	signal WX7387: std_logic; attribute dont_touch of WX7387: signal is true;
	signal WX7388: std_logic; attribute dont_touch of WX7388: signal is true;
	signal WX7389: std_logic; attribute dont_touch of WX7389: signal is true;
	signal WX7390: std_logic; attribute dont_touch of WX7390: signal is true;
	signal WX7391: std_logic; attribute dont_touch of WX7391: signal is true;
	signal WX7392: std_logic; attribute dont_touch of WX7392: signal is true;
	signal WX7393: std_logic; attribute dont_touch of WX7393: signal is true;
	signal WX7394: std_logic; attribute dont_touch of WX7394: signal is true;
	signal WX7395: std_logic; attribute dont_touch of WX7395: signal is true;
	signal WX7396: std_logic; attribute dont_touch of WX7396: signal is true;
	signal WX7397: std_logic; attribute dont_touch of WX7397: signal is true;
	signal WX7398: std_logic; attribute dont_touch of WX7398: signal is true;
	signal WX7399: std_logic; attribute dont_touch of WX7399: signal is true;
	signal WX7400: std_logic; attribute dont_touch of WX7400: signal is true;
	signal WX7401: std_logic; attribute dont_touch of WX7401: signal is true;
	signal WX7402: std_logic; attribute dont_touch of WX7402: signal is true;
	signal WX7403: std_logic; attribute dont_touch of WX7403: signal is true;
	signal WX7404: std_logic; attribute dont_touch of WX7404: signal is true;
	signal WX7405: std_logic; attribute dont_touch of WX7405: signal is true;
	signal WX7406: std_logic; attribute dont_touch of WX7406: signal is true;
	signal WX7407: std_logic; attribute dont_touch of WX7407: signal is true;
	signal WX7408: std_logic; attribute dont_touch of WX7408: signal is true;
	signal WX7409: std_logic; attribute dont_touch of WX7409: signal is true;
	signal WX7410: std_logic; attribute dont_touch of WX7410: signal is true;
	signal WX7411: std_logic; attribute dont_touch of WX7411: signal is true;
	signal WX7412: std_logic; attribute dont_touch of WX7412: signal is true;
	signal WX7413: std_logic; attribute dont_touch of WX7413: signal is true;
	signal WX7414: std_logic; attribute dont_touch of WX7414: signal is true;
	signal WX7415: std_logic; attribute dont_touch of WX7415: signal is true;
	signal WX7416: std_logic; attribute dont_touch of WX7416: signal is true;
	signal WX7417: std_logic; attribute dont_touch of WX7417: signal is true;
	signal WX7418: std_logic; attribute dont_touch of WX7418: signal is true;
	signal WX7419: std_logic; attribute dont_touch of WX7419: signal is true;
	signal WX7420: std_logic; attribute dont_touch of WX7420: signal is true;
	signal WX7421: std_logic; attribute dont_touch of WX7421: signal is true;
	signal WX7422: std_logic; attribute dont_touch of WX7422: signal is true;
	signal WX7423: std_logic; attribute dont_touch of WX7423: signal is true;
	signal WX7424: std_logic; attribute dont_touch of WX7424: signal is true;
	signal WX7425: std_logic; attribute dont_touch of WX7425: signal is true;
	signal WX7426: std_logic; attribute dont_touch of WX7426: signal is true;
	signal WX7427: std_logic; attribute dont_touch of WX7427: signal is true;
	signal WX7428: std_logic; attribute dont_touch of WX7428: signal is true;
	signal WX7429: std_logic; attribute dont_touch of WX7429: signal is true;
	signal WX7430: std_logic; attribute dont_touch of WX7430: signal is true;
	signal WX7431: std_logic; attribute dont_touch of WX7431: signal is true;
	signal WX7432: std_logic; attribute dont_touch of WX7432: signal is true;
	signal WX7433: std_logic; attribute dont_touch of WX7433: signal is true;
	signal WX7434: std_logic; attribute dont_touch of WX7434: signal is true;
	signal WX7435: std_logic; attribute dont_touch of WX7435: signal is true;
	signal WX7436: std_logic; attribute dont_touch of WX7436: signal is true;
	signal WX7437: std_logic; attribute dont_touch of WX7437: signal is true;
	signal WX7438: std_logic; attribute dont_touch of WX7438: signal is true;
	signal WX7439: std_logic; attribute dont_touch of WX7439: signal is true;
	signal WX7440: std_logic; attribute dont_touch of WX7440: signal is true;
	signal WX7441: std_logic; attribute dont_touch of WX7441: signal is true;
	signal WX7442: std_logic; attribute dont_touch of WX7442: signal is true;
	signal WX7443: std_logic; attribute dont_touch of WX7443: signal is true;
	signal WX7444: std_logic; attribute dont_touch of WX7444: signal is true;
	signal WX7445: std_logic; attribute dont_touch of WX7445: signal is true;
	signal WX7446: std_logic; attribute dont_touch of WX7446: signal is true;
	signal WX7447: std_logic; attribute dont_touch of WX7447: signal is true;
	signal WX7448: std_logic; attribute dont_touch of WX7448: signal is true;
	signal WX7449: std_logic; attribute dont_touch of WX7449: signal is true;
	signal WX7450: std_logic; attribute dont_touch of WX7450: signal is true;
	signal WX7451: std_logic; attribute dont_touch of WX7451: signal is true;
	signal WX7452: std_logic; attribute dont_touch of WX7452: signal is true;
	signal WX7453: std_logic; attribute dont_touch of WX7453: signal is true;
	signal WX7454: std_logic; attribute dont_touch of WX7454: signal is true;
	signal WX7455: std_logic; attribute dont_touch of WX7455: signal is true;
	signal WX7456: std_logic; attribute dont_touch of WX7456: signal is true;
	signal WX7457: std_logic; attribute dont_touch of WX7457: signal is true;
	signal WX7458: std_logic; attribute dont_touch of WX7458: signal is true;
	signal WX7459: std_logic; attribute dont_touch of WX7459: signal is true;
	signal WX7460: std_logic; attribute dont_touch of WX7460: signal is true;
	signal WX7461: std_logic; attribute dont_touch of WX7461: signal is true;
	signal WX7462: std_logic; attribute dont_touch of WX7462: signal is true;
	signal WX7463: std_logic; attribute dont_touch of WX7463: signal is true;
	signal WX7464: std_logic; attribute dont_touch of WX7464: signal is true;
	signal WX7465: std_logic; attribute dont_touch of WX7465: signal is true;
	signal WX7466: std_logic; attribute dont_touch of WX7466: signal is true;
	signal WX7467: std_logic; attribute dont_touch of WX7467: signal is true;
	signal WX7468: std_logic; attribute dont_touch of WX7468: signal is true;
	signal WX7469: std_logic; attribute dont_touch of WX7469: signal is true;
	signal WX7470: std_logic; attribute dont_touch of WX7470: signal is true;
	signal WX7471: std_logic; attribute dont_touch of WX7471: signal is true;
	signal WX7472: std_logic; attribute dont_touch of WX7472: signal is true;
	signal WX7473: std_logic; attribute dont_touch of WX7473: signal is true;
	signal WX7474: std_logic; attribute dont_touch of WX7474: signal is true;
	signal WX7475: std_logic; attribute dont_touch of WX7475: signal is true;
	signal WX7476: std_logic; attribute dont_touch of WX7476: signal is true;
	signal WX7477: std_logic; attribute dont_touch of WX7477: signal is true;
	signal WX7478: std_logic; attribute dont_touch of WX7478: signal is true;
	signal WX7479: std_logic; attribute dont_touch of WX7479: signal is true;
	signal WX7480: std_logic; attribute dont_touch of WX7480: signal is true;
	signal WX7481: std_logic; attribute dont_touch of WX7481: signal is true;
	signal WX7482: std_logic; attribute dont_touch of WX7482: signal is true;
	signal WX7483: std_logic; attribute dont_touch of WX7483: signal is true;
	signal WX7484: std_logic; attribute dont_touch of WX7484: signal is true;
	signal WX7485: std_logic; attribute dont_touch of WX7485: signal is true;
	signal WX7486: std_logic; attribute dont_touch of WX7486: signal is true;
	signal WX7487: std_logic; attribute dont_touch of WX7487: signal is true;
	signal WX7488: std_logic; attribute dont_touch of WX7488: signal is true;
	signal WX7489: std_logic; attribute dont_touch of WX7489: signal is true;
	signal WX7490: std_logic; attribute dont_touch of WX7490: signal is true;
	signal WX7491: std_logic; attribute dont_touch of WX7491: signal is true;
	signal WX7492: std_logic; attribute dont_touch of WX7492: signal is true;
	signal WX7493: std_logic; attribute dont_touch of WX7493: signal is true;
	signal WX7494: std_logic; attribute dont_touch of WX7494: signal is true;
	signal WX7495: std_logic; attribute dont_touch of WX7495: signal is true;
	signal WX7496: std_logic; attribute dont_touch of WX7496: signal is true;
	signal WX7497: std_logic; attribute dont_touch of WX7497: signal is true;
	signal WX7498: std_logic; attribute dont_touch of WX7498: signal is true;
	signal WX7499: std_logic; attribute dont_touch of WX7499: signal is true;
	signal WX7500: std_logic; attribute dont_touch of WX7500: signal is true;
	signal WX7501: std_logic; attribute dont_touch of WX7501: signal is true;
	signal WX7502: std_logic; attribute dont_touch of WX7502: signal is true;
	signal WX7503: std_logic; attribute dont_touch of WX7503: signal is true;
	signal WX7504: std_logic; attribute dont_touch of WX7504: signal is true;
	signal WX7505: std_logic; attribute dont_touch of WX7505: signal is true;
	signal WX7506: std_logic; attribute dont_touch of WX7506: signal is true;
	signal WX7507: std_logic; attribute dont_touch of WX7507: signal is true;
	signal WX7508: std_logic; attribute dont_touch of WX7508: signal is true;
	signal WX7509: std_logic; attribute dont_touch of WX7509: signal is true;
	signal WX7510: std_logic; attribute dont_touch of WX7510: signal is true;
	signal WX7511: std_logic; attribute dont_touch of WX7511: signal is true;
	signal WX7512: std_logic; attribute dont_touch of WX7512: signal is true;
	signal WX7513: std_logic; attribute dont_touch of WX7513: signal is true;
	signal WX7514: std_logic; attribute dont_touch of WX7514: signal is true;
	signal WX7515: std_logic; attribute dont_touch of WX7515: signal is true;
	signal WX7516: std_logic; attribute dont_touch of WX7516: signal is true;
	signal WX7517: std_logic; attribute dont_touch of WX7517: signal is true;
	signal WX7518: std_logic; attribute dont_touch of WX7518: signal is true;
	signal WX7519: std_logic; attribute dont_touch of WX7519: signal is true;
	signal WX7520: std_logic; attribute dont_touch of WX7520: signal is true;
	signal WX7521: std_logic; attribute dont_touch of WX7521: signal is true;
	signal WX7522: std_logic; attribute dont_touch of WX7522: signal is true;
	signal WX7523: std_logic; attribute dont_touch of WX7523: signal is true;
	signal WX7524: std_logic; attribute dont_touch of WX7524: signal is true;
	signal WX7525: std_logic; attribute dont_touch of WX7525: signal is true;
	signal WX7526: std_logic; attribute dont_touch of WX7526: signal is true;
	signal WX7527: std_logic; attribute dont_touch of WX7527: signal is true;
	signal WX7528: std_logic; attribute dont_touch of WX7528: signal is true;
	signal WX7529: std_logic; attribute dont_touch of WX7529: signal is true;
	signal WX7530: std_logic; attribute dont_touch of WX7530: signal is true;
	signal WX7531: std_logic; attribute dont_touch of WX7531: signal is true;
	signal WX7532: std_logic; attribute dont_touch of WX7532: signal is true;
	signal WX7533: std_logic; attribute dont_touch of WX7533: signal is true;
	signal WX7534: std_logic; attribute dont_touch of WX7534: signal is true;
	signal WX7535: std_logic; attribute dont_touch of WX7535: signal is true;
	signal WX7536: std_logic; attribute dont_touch of WX7536: signal is true;
	signal WX7537: std_logic; attribute dont_touch of WX7537: signal is true;
	signal WX7538: std_logic; attribute dont_touch of WX7538: signal is true;
	signal WX7539: std_logic; attribute dont_touch of WX7539: signal is true;
	signal WX7540: std_logic; attribute dont_touch of WX7540: signal is true;
	signal WX7541: std_logic; attribute dont_touch of WX7541: signal is true;
	signal WX7542: std_logic; attribute dont_touch of WX7542: signal is true;
	signal WX7543: std_logic; attribute dont_touch of WX7543: signal is true;
	signal WX7544: std_logic; attribute dont_touch of WX7544: signal is true;
	signal WX7545: std_logic; attribute dont_touch of WX7545: signal is true;
	signal WX7546: std_logic; attribute dont_touch of WX7546: signal is true;
	signal WX7547: std_logic; attribute dont_touch of WX7547: signal is true;
	signal WX7548: std_logic; attribute dont_touch of WX7548: signal is true;
	signal WX7549: std_logic; attribute dont_touch of WX7549: signal is true;
	signal WX7550: std_logic; attribute dont_touch of WX7550: signal is true;
	signal WX7551: std_logic; attribute dont_touch of WX7551: signal is true;
	signal WX7552: std_logic; attribute dont_touch of WX7552: signal is true;
	signal WX7553: std_logic; attribute dont_touch of WX7553: signal is true;
	signal WX7554: std_logic; attribute dont_touch of WX7554: signal is true;
	signal WX7555: std_logic; attribute dont_touch of WX7555: signal is true;
	signal WX7556: std_logic; attribute dont_touch of WX7556: signal is true;
	signal WX7557: std_logic; attribute dont_touch of WX7557: signal is true;
	signal WX7558: std_logic; attribute dont_touch of WX7558: signal is true;
	signal WX7559: std_logic; attribute dont_touch of WX7559: signal is true;
	signal WX7560: std_logic; attribute dont_touch of WX7560: signal is true;
	signal WX7561: std_logic; attribute dont_touch of WX7561: signal is true;
	signal WX7562: std_logic; attribute dont_touch of WX7562: signal is true;
	signal WX7563: std_logic; attribute dont_touch of WX7563: signal is true;
	signal WX7564: std_logic; attribute dont_touch of WX7564: signal is true;
	signal WX7565: std_logic; attribute dont_touch of WX7565: signal is true;
	signal WX7566: std_logic; attribute dont_touch of WX7566: signal is true;
	signal WX7567: std_logic; attribute dont_touch of WX7567: signal is true;
	signal WX7568: std_logic; attribute dont_touch of WX7568: signal is true;
	signal WX7569: std_logic; attribute dont_touch of WX7569: signal is true;
	signal WX7570: std_logic; attribute dont_touch of WX7570: signal is true;
	signal WX7571: std_logic; attribute dont_touch of WX7571: signal is true;
	signal WX7572: std_logic; attribute dont_touch of WX7572: signal is true;
	signal WX7573: std_logic; attribute dont_touch of WX7573: signal is true;
	signal WX7574: std_logic; attribute dont_touch of WX7574: signal is true;
	signal WX7575: std_logic; attribute dont_touch of WX7575: signal is true;
	signal WX7576: std_logic; attribute dont_touch of WX7576: signal is true;
	signal WX7577: std_logic; attribute dont_touch of WX7577: signal is true;
	signal WX7578: std_logic; attribute dont_touch of WX7578: signal is true;
	signal WX7579: std_logic; attribute dont_touch of WX7579: signal is true;
	signal WX7580: std_logic; attribute dont_touch of WX7580: signal is true;
	signal WX7581: std_logic; attribute dont_touch of WX7581: signal is true;
	signal WX7582: std_logic; attribute dont_touch of WX7582: signal is true;
	signal WX7583: std_logic; attribute dont_touch of WX7583: signal is true;
	signal WX7584: std_logic; attribute dont_touch of WX7584: signal is true;
	signal WX7585: std_logic; attribute dont_touch of WX7585: signal is true;
	signal WX7586: std_logic; attribute dont_touch of WX7586: signal is true;
	signal WX7587: std_logic; attribute dont_touch of WX7587: signal is true;
	signal WX7588: std_logic; attribute dont_touch of WX7588: signal is true;
	signal WX7589: std_logic; attribute dont_touch of WX7589: signal is true;
	signal WX7590: std_logic; attribute dont_touch of WX7590: signal is true;
	signal WX7591: std_logic; attribute dont_touch of WX7591: signal is true;
	signal WX7592: std_logic; attribute dont_touch of WX7592: signal is true;
	signal WX7593: std_logic; attribute dont_touch of WX7593: signal is true;
	signal WX7594: std_logic; attribute dont_touch of WX7594: signal is true;
	signal WX7595: std_logic; attribute dont_touch of WX7595: signal is true;
	signal WX7596: std_logic; attribute dont_touch of WX7596: signal is true;
	signal WX7597: std_logic; attribute dont_touch of WX7597: signal is true;
	signal WX7598: std_logic; attribute dont_touch of WX7598: signal is true;
	signal WX7599: std_logic; attribute dont_touch of WX7599: signal is true;
	signal WX7600: std_logic; attribute dont_touch of WX7600: signal is true;
	signal WX7601: std_logic; attribute dont_touch of WX7601: signal is true;
	signal WX7602: std_logic; attribute dont_touch of WX7602: signal is true;
	signal WX7603: std_logic; attribute dont_touch of WX7603: signal is true;
	signal WX7604: std_logic; attribute dont_touch of WX7604: signal is true;
	signal WX7605: std_logic; attribute dont_touch of WX7605: signal is true;
	signal WX7606: std_logic; attribute dont_touch of WX7606: signal is true;
	signal WX7607: std_logic; attribute dont_touch of WX7607: signal is true;
	signal WX7608: std_logic; attribute dont_touch of WX7608: signal is true;
	signal WX7609: std_logic; attribute dont_touch of WX7609: signal is true;
	signal WX7610: std_logic; attribute dont_touch of WX7610: signal is true;
	signal WX7611: std_logic; attribute dont_touch of WX7611: signal is true;
	signal WX7612: std_logic; attribute dont_touch of WX7612: signal is true;
	signal WX7613: std_logic; attribute dont_touch of WX7613: signal is true;
	signal WX7614: std_logic; attribute dont_touch of WX7614: signal is true;
	signal WX7615: std_logic; attribute dont_touch of WX7615: signal is true;
	signal WX7616: std_logic; attribute dont_touch of WX7616: signal is true;
	signal WX7617: std_logic; attribute dont_touch of WX7617: signal is true;
	signal WX7618: std_logic; attribute dont_touch of WX7618: signal is true;
	signal WX7619: std_logic; attribute dont_touch of WX7619: signal is true;
	signal WX7620: std_logic; attribute dont_touch of WX7620: signal is true;
	signal WX7621: std_logic; attribute dont_touch of WX7621: signal is true;
	signal WX7622: std_logic; attribute dont_touch of WX7622: signal is true;
	signal WX7623: std_logic; attribute dont_touch of WX7623: signal is true;
	signal WX7624: std_logic; attribute dont_touch of WX7624: signal is true;
	signal WX7625: std_logic; attribute dont_touch of WX7625: signal is true;
	signal WX7626: std_logic; attribute dont_touch of WX7626: signal is true;
	signal WX7627: std_logic; attribute dont_touch of WX7627: signal is true;
	signal WX7628: std_logic; attribute dont_touch of WX7628: signal is true;
	signal WX7629: std_logic; attribute dont_touch of WX7629: signal is true;
	signal WX7630: std_logic; attribute dont_touch of WX7630: signal is true;
	signal WX7631: std_logic; attribute dont_touch of WX7631: signal is true;
	signal WX7632: std_logic; attribute dont_touch of WX7632: signal is true;
	signal WX7633: std_logic; attribute dont_touch of WX7633: signal is true;
	signal WX7634: std_logic; attribute dont_touch of WX7634: signal is true;
	signal WX7635: std_logic; attribute dont_touch of WX7635: signal is true;
	signal WX7636: std_logic; attribute dont_touch of WX7636: signal is true;
	signal WX7637: std_logic; attribute dont_touch of WX7637: signal is true;
	signal WX7638: std_logic; attribute dont_touch of WX7638: signal is true;
	signal WX7639: std_logic; attribute dont_touch of WX7639: signal is true;
	signal WX7640: std_logic; attribute dont_touch of WX7640: signal is true;
	signal WX7641: std_logic; attribute dont_touch of WX7641: signal is true;
	signal WX7642: std_logic; attribute dont_touch of WX7642: signal is true;
	signal WX7643: std_logic; attribute dont_touch of WX7643: signal is true;
	signal WX7644: std_logic; attribute dont_touch of WX7644: signal is true;
	signal WX7645: std_logic; attribute dont_touch of WX7645: signal is true;
	signal WX7646: std_logic; attribute dont_touch of WX7646: signal is true;
	signal WX7647: std_logic; attribute dont_touch of WX7647: signal is true;
	signal WX7648: std_logic; attribute dont_touch of WX7648: signal is true;
	signal WX7649: std_logic; attribute dont_touch of WX7649: signal is true;
	signal WX7650: std_logic; attribute dont_touch of WX7650: signal is true;
	signal WX7651: std_logic; attribute dont_touch of WX7651: signal is true;
	signal WX7652: std_logic; attribute dont_touch of WX7652: signal is true;
	signal WX7653: std_logic; attribute dont_touch of WX7653: signal is true;
	signal WX7654: std_logic; attribute dont_touch of WX7654: signal is true;
	signal WX7655: std_logic; attribute dont_touch of WX7655: signal is true;
	signal WX7656: std_logic; attribute dont_touch of WX7656: signal is true;
	signal WX7657: std_logic; attribute dont_touch of WX7657: signal is true;
	signal WX7658: std_logic; attribute dont_touch of WX7658: signal is true;
	signal WX7659: std_logic; attribute dont_touch of WX7659: signal is true;
	signal WX7660: std_logic; attribute dont_touch of WX7660: signal is true;
	signal WX7661: std_logic; attribute dont_touch of WX7661: signal is true;
	signal WX7662: std_logic; attribute dont_touch of WX7662: signal is true;
	signal WX7663: std_logic; attribute dont_touch of WX7663: signal is true;
	signal WX7664: std_logic; attribute dont_touch of WX7664: signal is true;
	signal WX7665: std_logic; attribute dont_touch of WX7665: signal is true;
	signal WX7666: std_logic; attribute dont_touch of WX7666: signal is true;
	signal WX7667: std_logic; attribute dont_touch of WX7667: signal is true;
	signal WX7668: std_logic; attribute dont_touch of WX7668: signal is true;
	signal WX7669: std_logic; attribute dont_touch of WX7669: signal is true;
	signal WX7670: std_logic; attribute dont_touch of WX7670: signal is true;
	signal WX7671: std_logic; attribute dont_touch of WX7671: signal is true;
	signal WX7672: std_logic; attribute dont_touch of WX7672: signal is true;
	signal WX7673: std_logic; attribute dont_touch of WX7673: signal is true;
	signal WX7674: std_logic; attribute dont_touch of WX7674: signal is true;
	signal WX7675: std_logic; attribute dont_touch of WX7675: signal is true;
	signal WX7676: std_logic; attribute dont_touch of WX7676: signal is true;
	signal WX7677: std_logic; attribute dont_touch of WX7677: signal is true;
	signal WX7678: std_logic; attribute dont_touch of WX7678: signal is true;
	signal WX7679: std_logic; attribute dont_touch of WX7679: signal is true;
	signal WX7680: std_logic; attribute dont_touch of WX7680: signal is true;
	signal WX7681: std_logic; attribute dont_touch of WX7681: signal is true;
	signal WX7682: std_logic; attribute dont_touch of WX7682: signal is true;
	signal WX7683: std_logic; attribute dont_touch of WX7683: signal is true;
	signal WX7684: std_logic; attribute dont_touch of WX7684: signal is true;
	signal WX7685: std_logic; attribute dont_touch of WX7685: signal is true;
	signal WX7686: std_logic; attribute dont_touch of WX7686: signal is true;
	signal WX7687: std_logic; attribute dont_touch of WX7687: signal is true;
	signal WX7688: std_logic; attribute dont_touch of WX7688: signal is true;
	signal WX7689: std_logic; attribute dont_touch of WX7689: signal is true;
	signal WX7690: std_logic; attribute dont_touch of WX7690: signal is true;
	signal WX7691: std_logic; attribute dont_touch of WX7691: signal is true;
	signal WX7692: std_logic; attribute dont_touch of WX7692: signal is true;
	signal WX7693: std_logic; attribute dont_touch of WX7693: signal is true;
	signal WX7694: std_logic; attribute dont_touch of WX7694: signal is true;
	signal WX7695: std_logic; attribute dont_touch of WX7695: signal is true;
	signal WX7696: std_logic; attribute dont_touch of WX7696: signal is true;
	signal WX7697: std_logic; attribute dont_touch of WX7697: signal is true;
	signal WX7698: std_logic; attribute dont_touch of WX7698: signal is true;
	signal WX7699: std_logic; attribute dont_touch of WX7699: signal is true;
	signal WX7700: std_logic; attribute dont_touch of WX7700: signal is true;
	signal WX7701: std_logic; attribute dont_touch of WX7701: signal is true;
	signal WX7702: std_logic; attribute dont_touch of WX7702: signal is true;
	signal WX7703: std_logic; attribute dont_touch of WX7703: signal is true;
	signal WX7704: std_logic; attribute dont_touch of WX7704: signal is true;
	signal WX7705: std_logic; attribute dont_touch of WX7705: signal is true;
	signal WX7706: std_logic; attribute dont_touch of WX7706: signal is true;
	signal WX7707: std_logic; attribute dont_touch of WX7707: signal is true;
	signal WX7708: std_logic; attribute dont_touch of WX7708: signal is true;
	signal WX7709: std_logic; attribute dont_touch of WX7709: signal is true;
	signal WX7710: std_logic; attribute dont_touch of WX7710: signal is true;
	signal WX7711: std_logic; attribute dont_touch of WX7711: signal is true;
	signal WX7712: std_logic; attribute dont_touch of WX7712: signal is true;
	signal WX7713: std_logic; attribute dont_touch of WX7713: signal is true;
	signal WX7714: std_logic; attribute dont_touch of WX7714: signal is true;
	signal WX7715: std_logic; attribute dont_touch of WX7715: signal is true;
	signal WX7716: std_logic; attribute dont_touch of WX7716: signal is true;
	signal WX7717: std_logic; attribute dont_touch of WX7717: signal is true;
	signal WX7718: std_logic; attribute dont_touch of WX7718: signal is true;
	signal WX7719: std_logic; attribute dont_touch of WX7719: signal is true;
	signal WX7720: std_logic; attribute dont_touch of WX7720: signal is true;
	signal WX7721: std_logic; attribute dont_touch of WX7721: signal is true;
	signal WX7722: std_logic; attribute dont_touch of WX7722: signal is true;
	signal WX7723: std_logic; attribute dont_touch of WX7723: signal is true;
	signal WX7724: std_logic; attribute dont_touch of WX7724: signal is true;
	signal WX7725: std_logic; attribute dont_touch of WX7725: signal is true;
	signal WX7726: std_logic; attribute dont_touch of WX7726: signal is true;
	signal WX7727: std_logic; attribute dont_touch of WX7727: signal is true;
	signal WX7728: std_logic; attribute dont_touch of WX7728: signal is true;
	signal WX7729: std_logic; attribute dont_touch of WX7729: signal is true;
	signal WX7731: std_logic; attribute dont_touch of WX7731: signal is true;
	signal WX7733: std_logic; attribute dont_touch of WX7733: signal is true;
	signal WX7735: std_logic; attribute dont_touch of WX7735: signal is true;
	signal WX7737: std_logic; attribute dont_touch of WX7737: signal is true;
	signal WX7739: std_logic; attribute dont_touch of WX7739: signal is true;
	signal WX7741: std_logic; attribute dont_touch of WX7741: signal is true;
	signal WX7743: std_logic; attribute dont_touch of WX7743: signal is true;
	signal WX7745: std_logic; attribute dont_touch of WX7745: signal is true;
	signal WX7747: std_logic; attribute dont_touch of WX7747: signal is true;
	signal WX7749: std_logic; attribute dont_touch of WX7749: signal is true;
	signal WX7751: std_logic; attribute dont_touch of WX7751: signal is true;
	signal WX7753: std_logic; attribute dont_touch of WX7753: signal is true;
	signal WX7755: std_logic; attribute dont_touch of WX7755: signal is true;
	signal WX7757: std_logic; attribute dont_touch of WX7757: signal is true;
	signal WX7759: std_logic; attribute dont_touch of WX7759: signal is true;
	signal WX7761: std_logic; attribute dont_touch of WX7761: signal is true;
	signal WX7763: std_logic; attribute dont_touch of WX7763: signal is true;
	signal WX7765: std_logic; attribute dont_touch of WX7765: signal is true;
	signal WX7767: std_logic; attribute dont_touch of WX7767: signal is true;
	signal WX7769: std_logic; attribute dont_touch of WX7769: signal is true;
	signal WX7771: std_logic; attribute dont_touch of WX7771: signal is true;
	signal WX7773: std_logic; attribute dont_touch of WX7773: signal is true;
	signal WX7775: std_logic; attribute dont_touch of WX7775: signal is true;
	signal WX7777: std_logic; attribute dont_touch of WX7777: signal is true;
	signal WX7779: std_logic; attribute dont_touch of WX7779: signal is true;
	signal WX7781: std_logic; attribute dont_touch of WX7781: signal is true;
	signal WX7783: std_logic; attribute dont_touch of WX7783: signal is true;
	signal WX7785: std_logic; attribute dont_touch of WX7785: signal is true;
	signal WX7787: std_logic; attribute dont_touch of WX7787: signal is true;
	signal WX7789: std_logic; attribute dont_touch of WX7789: signal is true;
	signal WX7791: std_logic; attribute dont_touch of WX7791: signal is true;
	signal WX7793: std_logic; attribute dont_touch of WX7793: signal is true;
	signal WX7794: std_logic; attribute dont_touch of WX7794: signal is true;
	signal WX7795: std_logic; attribute dont_touch of WX7795: signal is true;
	signal WX7796: std_logic; attribute dont_touch of WX7796: signal is true;
	signal WX7797: std_logic; attribute dont_touch of WX7797: signal is true;
	signal WX7798: std_logic; attribute dont_touch of WX7798: signal is true;
	signal WX7799: std_logic; attribute dont_touch of WX7799: signal is true;
	signal WX7800: std_logic; attribute dont_touch of WX7800: signal is true;
	signal WX7801: std_logic; attribute dont_touch of WX7801: signal is true;
	signal WX7802: std_logic; attribute dont_touch of WX7802: signal is true;
	signal WX7803: std_logic; attribute dont_touch of WX7803: signal is true;
	signal WX7804: std_logic; attribute dont_touch of WX7804: signal is true;
	signal WX7805: std_logic; attribute dont_touch of WX7805: signal is true;
	signal WX7806: std_logic; attribute dont_touch of WX7806: signal is true;
	signal WX7807: std_logic; attribute dont_touch of WX7807: signal is true;
	signal WX7808: std_logic; attribute dont_touch of WX7808: signal is true;
	signal WX7809: std_logic; attribute dont_touch of WX7809: signal is true;
	signal WX7810: std_logic; attribute dont_touch of WX7810: signal is true;
	signal WX7811: std_logic; attribute dont_touch of WX7811: signal is true;
	signal WX7812: std_logic; attribute dont_touch of WX7812: signal is true;
	signal WX7813: std_logic; attribute dont_touch of WX7813: signal is true;
	signal WX7814: std_logic; attribute dont_touch of WX7814: signal is true;
	signal WX7815: std_logic; attribute dont_touch of WX7815: signal is true;
	signal WX7816: std_logic; attribute dont_touch of WX7816: signal is true;
	signal WX7817: std_logic; attribute dont_touch of WX7817: signal is true;
	signal WX7818: std_logic; attribute dont_touch of WX7818: signal is true;
	signal WX7819: std_logic; attribute dont_touch of WX7819: signal is true;
	signal WX7820: std_logic; attribute dont_touch of WX7820: signal is true;
	signal WX7821: std_logic; attribute dont_touch of WX7821: signal is true;
	signal WX7822: std_logic; attribute dont_touch of WX7822: signal is true;
	signal WX7823: std_logic; attribute dont_touch of WX7823: signal is true;
	signal WX7824: std_logic; attribute dont_touch of WX7824: signal is true;
	signal WX7825: std_logic; attribute dont_touch of WX7825: signal is true;
	signal WX7826: std_logic; attribute dont_touch of WX7826: signal is true;
	signal WX7827: std_logic; attribute dont_touch of WX7827: signal is true;
	signal WX7828: std_logic; attribute dont_touch of WX7828: signal is true;
	signal WX7829: std_logic; attribute dont_touch of WX7829: signal is true;
	signal WX7830: std_logic; attribute dont_touch of WX7830: signal is true;
	signal WX7831: std_logic; attribute dont_touch of WX7831: signal is true;
	signal WX7832: std_logic; attribute dont_touch of WX7832: signal is true;
	signal WX7833: std_logic; attribute dont_touch of WX7833: signal is true;
	signal WX7834: std_logic; attribute dont_touch of WX7834: signal is true;
	signal WX7835: std_logic; attribute dont_touch of WX7835: signal is true;
	signal WX7836: std_logic; attribute dont_touch of WX7836: signal is true;
	signal WX7837: std_logic; attribute dont_touch of WX7837: signal is true;
	signal WX7838: std_logic; attribute dont_touch of WX7838: signal is true;
	signal WX7839: std_logic; attribute dont_touch of WX7839: signal is true;
	signal WX7840: std_logic; attribute dont_touch of WX7840: signal is true;
	signal WX7841: std_logic; attribute dont_touch of WX7841: signal is true;
	signal WX7842: std_logic; attribute dont_touch of WX7842: signal is true;
	signal WX7843: std_logic; attribute dont_touch of WX7843: signal is true;
	signal WX7844: std_logic; attribute dont_touch of WX7844: signal is true;
	signal WX7845: std_logic; attribute dont_touch of WX7845: signal is true;
	signal WX7846: std_logic; attribute dont_touch of WX7846: signal is true;
	signal WX7847: std_logic; attribute dont_touch of WX7847: signal is true;
	signal WX7848: std_logic; attribute dont_touch of WX7848: signal is true;
	signal WX7849: std_logic; attribute dont_touch of WX7849: signal is true;
	signal WX7850: std_logic; attribute dont_touch of WX7850: signal is true;
	signal WX7851: std_logic; attribute dont_touch of WX7851: signal is true;
	signal WX7852: std_logic; attribute dont_touch of WX7852: signal is true;
	signal WX7853: std_logic; attribute dont_touch of WX7853: signal is true;
	signal WX7854: std_logic; attribute dont_touch of WX7854: signal is true;
	signal WX7855: std_logic; attribute dont_touch of WX7855: signal is true;
	signal WX7856: std_logic; attribute dont_touch of WX7856: signal is true;
	signal WX7857: std_logic; attribute dont_touch of WX7857: signal is true;
	signal WX7858: std_logic; attribute dont_touch of WX7858: signal is true;
	signal WX7859: std_logic; attribute dont_touch of WX7859: signal is true;
	signal WX7860: std_logic; attribute dont_touch of WX7860: signal is true;
	signal WX7861: std_logic; attribute dont_touch of WX7861: signal is true;
	signal WX7862: std_logic; attribute dont_touch of WX7862: signal is true;
	signal WX7863: std_logic; attribute dont_touch of WX7863: signal is true;
	signal WX7864: std_logic; attribute dont_touch of WX7864: signal is true;
	signal WX7865: std_logic; attribute dont_touch of WX7865: signal is true;
	signal WX7866: std_logic; attribute dont_touch of WX7866: signal is true;
	signal WX7867: std_logic; attribute dont_touch of WX7867: signal is true;
	signal WX7868: std_logic; attribute dont_touch of WX7868: signal is true;
	signal WX7869: std_logic; attribute dont_touch of WX7869: signal is true;
	signal WX7870: std_logic; attribute dont_touch of WX7870: signal is true;
	signal WX7871: std_logic; attribute dont_touch of WX7871: signal is true;
	signal WX7872: std_logic; attribute dont_touch of WX7872: signal is true;
	signal WX7873: std_logic; attribute dont_touch of WX7873: signal is true;
	signal WX7874: std_logic; attribute dont_touch of WX7874: signal is true;
	signal WX7875: std_logic; attribute dont_touch of WX7875: signal is true;
	signal WX7876: std_logic; attribute dont_touch of WX7876: signal is true;
	signal WX7877: std_logic; attribute dont_touch of WX7877: signal is true;
	signal WX7878: std_logic; attribute dont_touch of WX7878: signal is true;
	signal WX7879: std_logic; attribute dont_touch of WX7879: signal is true;
	signal WX7880: std_logic; attribute dont_touch of WX7880: signal is true;
	signal WX7881: std_logic; attribute dont_touch of WX7881: signal is true;
	signal WX7882: std_logic; attribute dont_touch of WX7882: signal is true;
	signal WX7883: std_logic; attribute dont_touch of WX7883: signal is true;
	signal WX7884: std_logic; attribute dont_touch of WX7884: signal is true;
	signal WX7885: std_logic; attribute dont_touch of WX7885: signal is true;
	signal WX7886: std_logic; attribute dont_touch of WX7886: signal is true;
	signal WX7887: std_logic; attribute dont_touch of WX7887: signal is true;
	signal WX7888: std_logic; attribute dont_touch of WX7888: signal is true;
	signal WX7889: std_logic; attribute dont_touch of WX7889: signal is true;
	signal WX7890: std_logic; attribute dont_touch of WX7890: signal is true;
	signal WX7891: std_logic; attribute dont_touch of WX7891: signal is true;
	signal WX7892: std_logic; attribute dont_touch of WX7892: signal is true;
	signal WX7893: std_logic; attribute dont_touch of WX7893: signal is true;
	signal WX7894: std_logic; attribute dont_touch of WX7894: signal is true;
	signal WX7895: std_logic; attribute dont_touch of WX7895: signal is true;
	signal WX7896: std_logic; attribute dont_touch of WX7896: signal is true;
	signal WX7897: std_logic; attribute dont_touch of WX7897: signal is true;
	signal WX7898: std_logic; attribute dont_touch of WX7898: signal is true;
	signal WX7899: std_logic; attribute dont_touch of WX7899: signal is true;
	signal WX7900: std_logic; attribute dont_touch of WX7900: signal is true;
	signal WX7901: std_logic; attribute dont_touch of WX7901: signal is true;
	signal WX7902: std_logic; attribute dont_touch of WX7902: signal is true;
	signal WX7903: std_logic; attribute dont_touch of WX7903: signal is true;
	signal WX7904: std_logic; attribute dont_touch of WX7904: signal is true;
	signal WX7905: std_logic; attribute dont_touch of WX7905: signal is true;
	signal WX7906: std_logic; attribute dont_touch of WX7906: signal is true;
	signal WX7907: std_logic; attribute dont_touch of WX7907: signal is true;
	signal WX7908: std_logic; attribute dont_touch of WX7908: signal is true;
	signal WX7909: std_logic; attribute dont_touch of WX7909: signal is true;
	signal WX7910: std_logic; attribute dont_touch of WX7910: signal is true;
	signal WX7911: std_logic; attribute dont_touch of WX7911: signal is true;
	signal WX7912: std_logic; attribute dont_touch of WX7912: signal is true;
	signal WX7913: std_logic; attribute dont_touch of WX7913: signal is true;
	signal WX7914: std_logic; attribute dont_touch of WX7914: signal is true;
	signal WX7915: std_logic; attribute dont_touch of WX7915: signal is true;
	signal WX7916: std_logic; attribute dont_touch of WX7916: signal is true;
	signal WX7917: std_logic; attribute dont_touch of WX7917: signal is true;
	signal WX7918: std_logic; attribute dont_touch of WX7918: signal is true;
	signal WX7919: std_logic; attribute dont_touch of WX7919: signal is true;
	signal WX7920: std_logic; attribute dont_touch of WX7920: signal is true;
	signal WX7921: std_logic; attribute dont_touch of WX7921: signal is true;
	signal WX7922: std_logic; attribute dont_touch of WX7922: signal is true;
	signal WX7923: std_logic; attribute dont_touch of WX7923: signal is true;
	signal WX7924: std_logic; attribute dont_touch of WX7924: signal is true;
	signal WX7925: std_logic; attribute dont_touch of WX7925: signal is true;
	signal WX7926: std_logic; attribute dont_touch of WX7926: signal is true;
	signal WX7927: std_logic; attribute dont_touch of WX7927: signal is true;
	signal WX7928: std_logic; attribute dont_touch of WX7928: signal is true;
	signal WX7929: std_logic; attribute dont_touch of WX7929: signal is true;
	signal WX7930: std_logic; attribute dont_touch of WX7930: signal is true;
	signal WX7931: std_logic; attribute dont_touch of WX7931: signal is true;
	signal WX7932: std_logic; attribute dont_touch of WX7932: signal is true;
	signal WX7933: std_logic; attribute dont_touch of WX7933: signal is true;
	signal WX7934: std_logic; attribute dont_touch of WX7934: signal is true;
	signal WX7935: std_logic; attribute dont_touch of WX7935: signal is true;
	signal WX7936: std_logic; attribute dont_touch of WX7936: signal is true;
	signal WX7937: std_logic; attribute dont_touch of WX7937: signal is true;
	signal WX7938: std_logic; attribute dont_touch of WX7938: signal is true;
	signal WX7939: std_logic; attribute dont_touch of WX7939: signal is true;
	signal WX7940: std_logic; attribute dont_touch of WX7940: signal is true;
	signal WX7941: std_logic; attribute dont_touch of WX7941: signal is true;
	signal WX7942: std_logic; attribute dont_touch of WX7942: signal is true;
	signal WX7943: std_logic; attribute dont_touch of WX7943: signal is true;
	signal WX7944: std_logic; attribute dont_touch of WX7944: signal is true;
	signal WX7945: std_logic; attribute dont_touch of WX7945: signal is true;
	signal WX7946: std_logic; attribute dont_touch of WX7946: signal is true;
	signal WX7947: std_logic; attribute dont_touch of WX7947: signal is true;
	signal WX7948: std_logic; attribute dont_touch of WX7948: signal is true;
	signal WX7949: std_logic; attribute dont_touch of WX7949: signal is true;
	signal WX7950: std_logic; attribute dont_touch of WX7950: signal is true;
	signal WX7951: std_logic; attribute dont_touch of WX7951: signal is true;
	signal WX7952: std_logic; attribute dont_touch of WX7952: signal is true;
	signal WX7953: std_logic; attribute dont_touch of WX7953: signal is true;
	signal WX7954: std_logic; attribute dont_touch of WX7954: signal is true;
	signal WX7955: std_logic; attribute dont_touch of WX7955: signal is true;
	signal WX7956: std_logic; attribute dont_touch of WX7956: signal is true;
	signal WX7957: std_logic; attribute dont_touch of WX7957: signal is true;
	signal WX7958: std_logic; attribute dont_touch of WX7958: signal is true;
	signal WX7959: std_logic; attribute dont_touch of WX7959: signal is true;
	signal WX7960: std_logic; attribute dont_touch of WX7960: signal is true;
	signal WX7961: std_logic; attribute dont_touch of WX7961: signal is true;
	signal WX7962: std_logic; attribute dont_touch of WX7962: signal is true;
	signal WX7963: std_logic; attribute dont_touch of WX7963: signal is true;
	signal WX7964: std_logic; attribute dont_touch of WX7964: signal is true;
	signal WX7965: std_logic; attribute dont_touch of WX7965: signal is true;
	signal WX7966: std_logic; attribute dont_touch of WX7966: signal is true;
	signal WX7967: std_logic; attribute dont_touch of WX7967: signal is true;
	signal WX7968: std_logic; attribute dont_touch of WX7968: signal is true;
	signal WX7969: std_logic; attribute dont_touch of WX7969: signal is true;
	signal WX7970: std_logic; attribute dont_touch of WX7970: signal is true;
	signal WX7971: std_logic; attribute dont_touch of WX7971: signal is true;
	signal WX7972: std_logic; attribute dont_touch of WX7972: signal is true;
	signal WX7973: std_logic; attribute dont_touch of WX7973: signal is true;
	signal WX7974: std_logic; attribute dont_touch of WX7974: signal is true;
	signal WX7975: std_logic; attribute dont_touch of WX7975: signal is true;
	signal WX7976: std_logic; attribute dont_touch of WX7976: signal is true;
	signal WX7977: std_logic; attribute dont_touch of WX7977: signal is true;
	signal WX7978: std_logic; attribute dont_touch of WX7978: signal is true;
	signal WX7979: std_logic; attribute dont_touch of WX7979: signal is true;
	signal WX7980: std_logic; attribute dont_touch of WX7980: signal is true;
	signal WX7981: std_logic; attribute dont_touch of WX7981: signal is true;
	signal WX7982: std_logic; attribute dont_touch of WX7982: signal is true;
	signal WX7983: std_logic; attribute dont_touch of WX7983: signal is true;
	signal WX7984: std_logic; attribute dont_touch of WX7984: signal is true;
	signal WX7985: std_logic; attribute dont_touch of WX7985: signal is true;
	signal WX7986: std_logic; attribute dont_touch of WX7986: signal is true;
	signal WX7987: std_logic; attribute dont_touch of WX7987: signal is true;
	signal WX7988: std_logic; attribute dont_touch of WX7988: signal is true;
	signal WX7989: std_logic; attribute dont_touch of WX7989: signal is true;
	signal WX7990: std_logic; attribute dont_touch of WX7990: signal is true;
	signal WX7991: std_logic; attribute dont_touch of WX7991: signal is true;
	signal WX7992: std_logic; attribute dont_touch of WX7992: signal is true;
	signal WX7993: std_logic; attribute dont_touch of WX7993: signal is true;
	signal WX7994: std_logic; attribute dont_touch of WX7994: signal is true;
	signal WX7995: std_logic; attribute dont_touch of WX7995: signal is true;
	signal WX7996: std_logic; attribute dont_touch of WX7996: signal is true;
	signal WX7997: std_logic; attribute dont_touch of WX7997: signal is true;
	signal WX7998: std_logic; attribute dont_touch of WX7998: signal is true;
	signal WX7999: std_logic; attribute dont_touch of WX7999: signal is true;
	signal WX8000: std_logic; attribute dont_touch of WX8000: signal is true;
	signal WX8001: std_logic; attribute dont_touch of WX8001: signal is true;
	signal WX8002: std_logic; attribute dont_touch of WX8002: signal is true;
	signal WX8003: std_logic; attribute dont_touch of WX8003: signal is true;
	signal WX8004: std_logic; attribute dont_touch of WX8004: signal is true;
	signal WX8005: std_logic; attribute dont_touch of WX8005: signal is true;
	signal WX8006: std_logic; attribute dont_touch of WX8006: signal is true;
	signal WX8007: std_logic; attribute dont_touch of WX8007: signal is true;
	signal WX8008: std_logic; attribute dont_touch of WX8008: signal is true;
	signal WX8009: std_logic; attribute dont_touch of WX8009: signal is true;
	signal WX8010: std_logic; attribute dont_touch of WX8010: signal is true;
	signal WX8011: std_logic; attribute dont_touch of WX8011: signal is true;
	signal WX8012: std_logic; attribute dont_touch of WX8012: signal is true;
	signal WX8013: std_logic; attribute dont_touch of WX8013: signal is true;
	signal WX8014: std_logic; attribute dont_touch of WX8014: signal is true;
	signal WX8015: std_logic; attribute dont_touch of WX8015: signal is true;
	signal WX8016: std_logic; attribute dont_touch of WX8016: signal is true;
	signal WX8017: std_logic; attribute dont_touch of WX8017: signal is true;
	signal WX8018: std_logic; attribute dont_touch of WX8018: signal is true;
	signal WX8019: std_logic; attribute dont_touch of WX8019: signal is true;
	signal WX8020: std_logic; attribute dont_touch of WX8020: signal is true;
	signal WX8021: std_logic; attribute dont_touch of WX8021: signal is true;
	signal WX8022: std_logic; attribute dont_touch of WX8022: signal is true;
	signal WX8023: std_logic; attribute dont_touch of WX8023: signal is true;
	signal WX8024: std_logic; attribute dont_touch of WX8024: signal is true;
	signal WX8025: std_logic; attribute dont_touch of WX8025: signal is true;
	signal WX8026: std_logic; attribute dont_touch of WX8026: signal is true;
	signal WX8027: std_logic; attribute dont_touch of WX8027: signal is true;
	signal WX8028: std_logic; attribute dont_touch of WX8028: signal is true;
	signal WX8029: std_logic; attribute dont_touch of WX8029: signal is true;
	signal WX8030: std_logic; attribute dont_touch of WX8030: signal is true;
	signal WX8031: std_logic; attribute dont_touch of WX8031: signal is true;
	signal WX8032: std_logic; attribute dont_touch of WX8032: signal is true;
	signal WX8033: std_logic; attribute dont_touch of WX8033: signal is true;
	signal WX8034: std_logic; attribute dont_touch of WX8034: signal is true;
	signal WX8035: std_logic; attribute dont_touch of WX8035: signal is true;
	signal WX8036: std_logic; attribute dont_touch of WX8036: signal is true;
	signal WX8037: std_logic; attribute dont_touch of WX8037: signal is true;
	signal WX8038: std_logic; attribute dont_touch of WX8038: signal is true;
	signal WX8039: std_logic; attribute dont_touch of WX8039: signal is true;
	signal WX8040: std_logic; attribute dont_touch of WX8040: signal is true;
	signal WX8041: std_logic; attribute dont_touch of WX8041: signal is true;
	signal WX8042: std_logic; attribute dont_touch of WX8042: signal is true;
	signal WX8043: std_logic; attribute dont_touch of WX8043: signal is true;
	signal WX8044: std_logic; attribute dont_touch of WX8044: signal is true;
	signal WX8045: std_logic; attribute dont_touch of WX8045: signal is true;
	signal WX8046: std_logic; attribute dont_touch of WX8046: signal is true;
	signal WX8047: std_logic; attribute dont_touch of WX8047: signal is true;
	signal WX8048: std_logic; attribute dont_touch of WX8048: signal is true;
	signal WX8049: std_logic; attribute dont_touch of WX8049: signal is true;
	signal WX8050: std_logic; attribute dont_touch of WX8050: signal is true;
	signal WX8051: std_logic; attribute dont_touch of WX8051: signal is true;
	signal WX8052: std_logic; attribute dont_touch of WX8052: signal is true;
	signal WX8053: std_logic; attribute dont_touch of WX8053: signal is true;
	signal WX8054: std_logic; attribute dont_touch of WX8054: signal is true;
	signal WX8055: std_logic; attribute dont_touch of WX8055: signal is true;
	signal WX8056: std_logic; attribute dont_touch of WX8056: signal is true;
	signal WX8057: std_logic; attribute dont_touch of WX8057: signal is true;
	signal WX8058: std_logic; attribute dont_touch of WX8058: signal is true;
	signal WX8059: std_logic; attribute dont_touch of WX8059: signal is true;
	signal WX8060: std_logic; attribute dont_touch of WX8060: signal is true;
	signal WX8061: std_logic; attribute dont_touch of WX8061: signal is true;
	signal WX8062: std_logic; attribute dont_touch of WX8062: signal is true;
	signal WX8063: std_logic; attribute dont_touch of WX8063: signal is true;
	signal WX8064: std_logic; attribute dont_touch of WX8064: signal is true;
	signal WX8065: std_logic; attribute dont_touch of WX8065: signal is true;
	signal WX8066: std_logic; attribute dont_touch of WX8066: signal is true;
	signal WX8067: std_logic; attribute dont_touch of WX8067: signal is true;
	signal WX8068: std_logic; attribute dont_touch of WX8068: signal is true;
	signal WX8069: std_logic; attribute dont_touch of WX8069: signal is true;
	signal WX8070: std_logic; attribute dont_touch of WX8070: signal is true;
	signal WX8071: std_logic; attribute dont_touch of WX8071: signal is true;
	signal WX8072: std_logic; attribute dont_touch of WX8072: signal is true;
	signal WX8073: std_logic; attribute dont_touch of WX8073: signal is true;
	signal WX8074: std_logic; attribute dont_touch of WX8074: signal is true;
	signal WX8075: std_logic; attribute dont_touch of WX8075: signal is true;
	signal WX8076: std_logic; attribute dont_touch of WX8076: signal is true;
	signal WX8077: std_logic; attribute dont_touch of WX8077: signal is true;
	signal WX8078: std_logic; attribute dont_touch of WX8078: signal is true;
	signal WX8079: std_logic; attribute dont_touch of WX8079: signal is true;
	signal WX8080: std_logic; attribute dont_touch of WX8080: signal is true;
	signal WX8081: std_logic; attribute dont_touch of WX8081: signal is true;
	signal WX8082: std_logic; attribute dont_touch of WX8082: signal is true;
	signal WX8083: std_logic; attribute dont_touch of WX8083: signal is true;
	signal WX8084: std_logic; attribute dont_touch of WX8084: signal is true;
	signal WX8085: std_logic; attribute dont_touch of WX8085: signal is true;
	signal WX8086: std_logic; attribute dont_touch of WX8086: signal is true;
	signal WX8087: std_logic; attribute dont_touch of WX8087: signal is true;
	signal WX8088: std_logic; attribute dont_touch of WX8088: signal is true;
	signal WX8089: std_logic; attribute dont_touch of WX8089: signal is true;
	signal WX8090: std_logic; attribute dont_touch of WX8090: signal is true;
	signal WX8091: std_logic; attribute dont_touch of WX8091: signal is true;
	signal WX8092: std_logic; attribute dont_touch of WX8092: signal is true;
	signal WX8093: std_logic; attribute dont_touch of WX8093: signal is true;
	signal WX8094: std_logic; attribute dont_touch of WX8094: signal is true;
	signal WX8095: std_logic; attribute dont_touch of WX8095: signal is true;
	signal WX8096: std_logic; attribute dont_touch of WX8096: signal is true;
	signal WX8097: std_logic; attribute dont_touch of WX8097: signal is true;
	signal WX8098: std_logic; attribute dont_touch of WX8098: signal is true;
	signal WX8099: std_logic; attribute dont_touch of WX8099: signal is true;
	signal WX8100: std_logic; attribute dont_touch of WX8100: signal is true;
	signal WX8101: std_logic; attribute dont_touch of WX8101: signal is true;
	signal WX8102: std_logic; attribute dont_touch of WX8102: signal is true;
	signal WX8103: std_logic; attribute dont_touch of WX8103: signal is true;
	signal WX8104: std_logic; attribute dont_touch of WX8104: signal is true;
	signal WX8105: std_logic; attribute dont_touch of WX8105: signal is true;
	signal WX8106: std_logic; attribute dont_touch of WX8106: signal is true;
	signal WX8107: std_logic; attribute dont_touch of WX8107: signal is true;
	signal WX8108: std_logic; attribute dont_touch of WX8108: signal is true;
	signal WX8109: std_logic; attribute dont_touch of WX8109: signal is true;
	signal WX8110: std_logic; attribute dont_touch of WX8110: signal is true;
	signal WX8111: std_logic; attribute dont_touch of WX8111: signal is true;
	signal WX8112: std_logic; attribute dont_touch of WX8112: signal is true;
	signal WX8113: std_logic; attribute dont_touch of WX8113: signal is true;
	signal WX8114: std_logic; attribute dont_touch of WX8114: signal is true;
	signal WX8115: std_logic; attribute dont_touch of WX8115: signal is true;
	signal WX8116: std_logic; attribute dont_touch of WX8116: signal is true;
	signal WX8117: std_logic; attribute dont_touch of WX8117: signal is true;
	signal WX8118: std_logic; attribute dont_touch of WX8118: signal is true;
	signal WX8119: std_logic; attribute dont_touch of WX8119: signal is true;
	signal WX8120: std_logic; attribute dont_touch of WX8120: signal is true;
	signal WX8121: std_logic; attribute dont_touch of WX8121: signal is true;
	signal WX8122: std_logic; attribute dont_touch of WX8122: signal is true;
	signal WX8123: std_logic; attribute dont_touch of WX8123: signal is true;
	signal WX8124: std_logic; attribute dont_touch of WX8124: signal is true;
	signal WX8125: std_logic; attribute dont_touch of WX8125: signal is true;
	signal WX8126: std_logic; attribute dont_touch of WX8126: signal is true;
	signal WX8127: std_logic; attribute dont_touch of WX8127: signal is true;
	signal WX8128: std_logic; attribute dont_touch of WX8128: signal is true;
	signal WX8129: std_logic; attribute dont_touch of WX8129: signal is true;
	signal WX8130: std_logic; attribute dont_touch of WX8130: signal is true;
	signal WX8131: std_logic; attribute dont_touch of WX8131: signal is true;
	signal WX8132: std_logic; attribute dont_touch of WX8132: signal is true;
	signal WX8133: std_logic; attribute dont_touch of WX8133: signal is true;
	signal WX8134: std_logic; attribute dont_touch of WX8134: signal is true;
	signal WX8135: std_logic; attribute dont_touch of WX8135: signal is true;
	signal WX8136: std_logic; attribute dont_touch of WX8136: signal is true;
	signal WX8137: std_logic; attribute dont_touch of WX8137: signal is true;
	signal WX8138: std_logic; attribute dont_touch of WX8138: signal is true;
	signal WX8139: std_logic; attribute dont_touch of WX8139: signal is true;
	signal WX8140: std_logic; attribute dont_touch of WX8140: signal is true;
	signal WX8141: std_logic; attribute dont_touch of WX8141: signal is true;
	signal WX8142: std_logic; attribute dont_touch of WX8142: signal is true;
	signal WX8143: std_logic; attribute dont_touch of WX8143: signal is true;
	signal WX8144: std_logic; attribute dont_touch of WX8144: signal is true;
	signal WX8145: std_logic; attribute dont_touch of WX8145: signal is true;
	signal WX8146: std_logic; attribute dont_touch of WX8146: signal is true;
	signal WX8147: std_logic; attribute dont_touch of WX8147: signal is true;
	signal WX8148: std_logic; attribute dont_touch of WX8148: signal is true;
	signal WX8149: std_logic; attribute dont_touch of WX8149: signal is true;
	signal WX8150: std_logic; attribute dont_touch of WX8150: signal is true;
	signal WX8151: std_logic; attribute dont_touch of WX8151: signal is true;
	signal WX8152: std_logic; attribute dont_touch of WX8152: signal is true;
	signal WX8153: std_logic; attribute dont_touch of WX8153: signal is true;
	signal WX8154: std_logic; attribute dont_touch of WX8154: signal is true;
	signal WX8155: std_logic; attribute dont_touch of WX8155: signal is true;
	signal WX8156: std_logic; attribute dont_touch of WX8156: signal is true;
	signal WX8157: std_logic; attribute dont_touch of WX8157: signal is true;
	signal WX8158: std_logic; attribute dont_touch of WX8158: signal is true;
	signal WX8159: std_logic; attribute dont_touch of WX8159: signal is true;
	signal WX8160: std_logic; attribute dont_touch of WX8160: signal is true;
	signal WX8161: std_logic; attribute dont_touch of WX8161: signal is true;
	signal WX8162: std_logic; attribute dont_touch of WX8162: signal is true;
	signal WX8163: std_logic; attribute dont_touch of WX8163: signal is true;
	signal WX8164: std_logic; attribute dont_touch of WX8164: signal is true;
	signal WX8165: std_logic; attribute dont_touch of WX8165: signal is true;
	signal WX8166: std_logic; attribute dont_touch of WX8166: signal is true;
	signal WX8167: std_logic; attribute dont_touch of WX8167: signal is true;
	signal WX8168: std_logic; attribute dont_touch of WX8168: signal is true;
	signal WX8169: std_logic; attribute dont_touch of WX8169: signal is true;
	signal WX8170: std_logic; attribute dont_touch of WX8170: signal is true;
	signal WX8171: std_logic; attribute dont_touch of WX8171: signal is true;
	signal WX8172: std_logic; attribute dont_touch of WX8172: signal is true;
	signal WX8173: std_logic; attribute dont_touch of WX8173: signal is true;
	signal WX8174: std_logic; attribute dont_touch of WX8174: signal is true;
	signal WX8175: std_logic; attribute dont_touch of WX8175: signal is true;
	signal WX8176: std_logic; attribute dont_touch of WX8176: signal is true;
	signal WX8177: std_logic; attribute dont_touch of WX8177: signal is true;
	signal WX8178: std_logic; attribute dont_touch of WX8178: signal is true;
	signal WX8179: std_logic; attribute dont_touch of WX8179: signal is true;
	signal WX8180: std_logic; attribute dont_touch of WX8180: signal is true;
	signal WX8181: std_logic; attribute dont_touch of WX8181: signal is true;
	signal WX8182: std_logic; attribute dont_touch of WX8182: signal is true;
	signal WX8183: std_logic; attribute dont_touch of WX8183: signal is true;
	signal WX8184: std_logic; attribute dont_touch of WX8184: signal is true;
	signal WX8185: std_logic; attribute dont_touch of WX8185: signal is true;
	signal WX8186: std_logic; attribute dont_touch of WX8186: signal is true;
	signal WX8187: std_logic; attribute dont_touch of WX8187: signal is true;
	signal WX8188: std_logic; attribute dont_touch of WX8188: signal is true;
	signal WX8189: std_logic; attribute dont_touch of WX8189: signal is true;
	signal WX8190: std_logic; attribute dont_touch of WX8190: signal is true;
	signal WX8191: std_logic; attribute dont_touch of WX8191: signal is true;
	signal WX8192: std_logic; attribute dont_touch of WX8192: signal is true;
	signal WX8193: std_logic; attribute dont_touch of WX8193: signal is true;
	signal WX8194: std_logic; attribute dont_touch of WX8194: signal is true;
	signal WX8195: std_logic; attribute dont_touch of WX8195: signal is true;
	signal WX8196: std_logic; attribute dont_touch of WX8196: signal is true;
	signal WX8197: std_logic; attribute dont_touch of WX8197: signal is true;
	signal WX8198: std_logic; attribute dont_touch of WX8198: signal is true;
	signal WX8199: std_logic; attribute dont_touch of WX8199: signal is true;
	signal WX8200: std_logic; attribute dont_touch of WX8200: signal is true;
	signal WX8201: std_logic; attribute dont_touch of WX8201: signal is true;
	signal WX8202: std_logic; attribute dont_touch of WX8202: signal is true;
	signal WX8203: std_logic; attribute dont_touch of WX8203: signal is true;
	signal WX8204: std_logic; attribute dont_touch of WX8204: signal is true;
	signal WX8205: std_logic; attribute dont_touch of WX8205: signal is true;
	signal WX8206: std_logic; attribute dont_touch of WX8206: signal is true;
	signal WX8207: std_logic; attribute dont_touch of WX8207: signal is true;
	signal WX8208: std_logic; attribute dont_touch of WX8208: signal is true;
	signal WX8209: std_logic; attribute dont_touch of WX8209: signal is true;
	signal WX8210: std_logic; attribute dont_touch of WX8210: signal is true;
	signal WX8211: std_logic; attribute dont_touch of WX8211: signal is true;
	signal WX8212: std_logic; attribute dont_touch of WX8212: signal is true;
	signal WX8213: std_logic; attribute dont_touch of WX8213: signal is true;
	signal WX8214: std_logic; attribute dont_touch of WX8214: signal is true;
	signal WX8215: std_logic; attribute dont_touch of WX8215: signal is true;
	signal WX8216: std_logic; attribute dont_touch of WX8216: signal is true;
	signal WX8217: std_logic; attribute dont_touch of WX8217: signal is true;
	signal WX8218: std_logic; attribute dont_touch of WX8218: signal is true;
	signal WX8219: std_logic; attribute dont_touch of WX8219: signal is true;
	signal WX8220: std_logic; attribute dont_touch of WX8220: signal is true;
	signal WX8221: std_logic; attribute dont_touch of WX8221: signal is true;
	signal WX8222: std_logic; attribute dont_touch of WX8222: signal is true;
	signal WX8223: std_logic; attribute dont_touch of WX8223: signal is true;
	signal WX8224: std_logic; attribute dont_touch of WX8224: signal is true;
	signal WX8225: std_logic; attribute dont_touch of WX8225: signal is true;
	signal WX8226: std_logic; attribute dont_touch of WX8226: signal is true;
	signal WX8227: std_logic; attribute dont_touch of WX8227: signal is true;
	signal WX8228: std_logic; attribute dont_touch of WX8228: signal is true;
	signal WX8229: std_logic; attribute dont_touch of WX8229: signal is true;
	signal WX8230: std_logic; attribute dont_touch of WX8230: signal is true;
	signal WX8231: std_logic; attribute dont_touch of WX8231: signal is true;
	signal WX8232: std_logic; attribute dont_touch of WX8232: signal is true;
	signal WX8233: std_logic; attribute dont_touch of WX8233: signal is true;
	signal WX8234: std_logic; attribute dont_touch of WX8234: signal is true;
	signal WX8235: std_logic; attribute dont_touch of WX8235: signal is true;
	signal WX8236: std_logic; attribute dont_touch of WX8236: signal is true;
	signal WX8237: std_logic; attribute dont_touch of WX8237: signal is true;
	signal WX8238: std_logic; attribute dont_touch of WX8238: signal is true;
	signal WX8239: std_logic; attribute dont_touch of WX8239: signal is true;
	signal WX8240: std_logic; attribute dont_touch of WX8240: signal is true;
	signal WX8241: std_logic; attribute dont_touch of WX8241: signal is true;
	signal WX8242: std_logic; attribute dont_touch of WX8242: signal is true;
	signal WX8243: std_logic; attribute dont_touch of WX8243: signal is true;
	signal WX8244: std_logic; attribute dont_touch of WX8244: signal is true;
	signal WX8245: std_logic; attribute dont_touch of WX8245: signal is true;
	signal WX8246: std_logic; attribute dont_touch of WX8246: signal is true;
	signal WX8247: std_logic; attribute dont_touch of WX8247: signal is true;
	signal WX8248: std_logic; attribute dont_touch of WX8248: signal is true;
	signal WX8249: std_logic; attribute dont_touch of WX8249: signal is true;
	signal WX8250: std_logic; attribute dont_touch of WX8250: signal is true;
	signal WX8251: std_logic; attribute dont_touch of WX8251: signal is true;
	signal WX8252: std_logic; attribute dont_touch of WX8252: signal is true;
	signal WX8253: std_logic; attribute dont_touch of WX8253: signal is true;
	signal WX8254: std_logic; attribute dont_touch of WX8254: signal is true;
	signal WX8255: std_logic; attribute dont_touch of WX8255: signal is true;
	signal WX8256: std_logic; attribute dont_touch of WX8256: signal is true;
	signal WX8257: std_logic; attribute dont_touch of WX8257: signal is true;
	signal WX8258: std_logic; attribute dont_touch of WX8258: signal is true;
	signal WX8259: std_logic; attribute dont_touch of WX8259: signal is true;
	signal WX8260: std_logic; attribute dont_touch of WX8260: signal is true;
	signal WX8261: std_logic; attribute dont_touch of WX8261: signal is true;
	signal WX8262: std_logic; attribute dont_touch of WX8262: signal is true;
	signal WX8263: std_logic; attribute dont_touch of WX8263: signal is true;
	signal WX8264: std_logic; attribute dont_touch of WX8264: signal is true;
	signal WX8265: std_logic; attribute dont_touch of WX8265: signal is true;
	signal WX8266: std_logic; attribute dont_touch of WX8266: signal is true;
	signal WX8267: std_logic; attribute dont_touch of WX8267: signal is true;
	signal WX8268: std_logic; attribute dont_touch of WX8268: signal is true;
	signal WX8269: std_logic; attribute dont_touch of WX8269: signal is true;
	signal WX8270: std_logic; attribute dont_touch of WX8270: signal is true;
	signal WX8271: std_logic; attribute dont_touch of WX8271: signal is true;
	signal WX8272: std_logic; attribute dont_touch of WX8272: signal is true;
	signal WX8273: std_logic; attribute dont_touch of WX8273: signal is true;
	signal WX8274: std_logic; attribute dont_touch of WX8274: signal is true;
	signal WX8275: std_logic; attribute dont_touch of WX8275: signal is true;
	signal WX8276: std_logic; attribute dont_touch of WX8276: signal is true;
	signal WX8277: std_logic; attribute dont_touch of WX8277: signal is true;
	signal WX8278: std_logic; attribute dont_touch of WX8278: signal is true;
	signal WX8279: std_logic; attribute dont_touch of WX8279: signal is true;
	signal WX8280: std_logic; attribute dont_touch of WX8280: signal is true;
	signal WX8281: std_logic; attribute dont_touch of WX8281: signal is true;
	signal WX8282: std_logic; attribute dont_touch of WX8282: signal is true;
	signal WX8283: std_logic; attribute dont_touch of WX8283: signal is true;
	signal WX8284: std_logic; attribute dont_touch of WX8284: signal is true;
	signal WX8285: std_logic; attribute dont_touch of WX8285: signal is true;
	signal WX8286: std_logic; attribute dont_touch of WX8286: signal is true;
	signal WX8287: std_logic; attribute dont_touch of WX8287: signal is true;
	signal WX8288: std_logic; attribute dont_touch of WX8288: signal is true;
	signal WX8289: std_logic; attribute dont_touch of WX8289: signal is true;
	signal WX8290: std_logic; attribute dont_touch of WX8290: signal is true;
	signal WX8291: std_logic; attribute dont_touch of WX8291: signal is true;
	signal WX8292: std_logic; attribute dont_touch of WX8292: signal is true;
	signal WX8293: std_logic; attribute dont_touch of WX8293: signal is true;
	signal WX8294: std_logic; attribute dont_touch of WX8294: signal is true;
	signal WX8295: std_logic; attribute dont_touch of WX8295: signal is true;
	signal WX8296: std_logic; attribute dont_touch of WX8296: signal is true;
	signal WX8297: std_logic; attribute dont_touch of WX8297: signal is true;
	signal WX8298: std_logic; attribute dont_touch of WX8298: signal is true;
	signal WX8299: std_logic; attribute dont_touch of WX8299: signal is true;
	signal WX8300: std_logic; attribute dont_touch of WX8300: signal is true;
	signal WX8301: std_logic; attribute dont_touch of WX8301: signal is true;
	signal WX8302: std_logic; attribute dont_touch of WX8302: signal is true;
	signal WX8303: std_logic; attribute dont_touch of WX8303: signal is true;
	signal WX8304: std_logic; attribute dont_touch of WX8304: signal is true;
	signal WX8305: std_logic; attribute dont_touch of WX8305: signal is true;
	signal WX8306: std_logic; attribute dont_touch of WX8306: signal is true;
	signal WX8307: std_logic; attribute dont_touch of WX8307: signal is true;
	signal WX8308: std_logic; attribute dont_touch of WX8308: signal is true;
	signal WX8309: std_logic; attribute dont_touch of WX8309: signal is true;
	signal WX8310: std_logic; attribute dont_touch of WX8310: signal is true;
	signal WX8311: std_logic; attribute dont_touch of WX8311: signal is true;
	signal WX8312: std_logic; attribute dont_touch of WX8312: signal is true;
	signal WX8313: std_logic; attribute dont_touch of WX8313: signal is true;
	signal WX8314: std_logic; attribute dont_touch of WX8314: signal is true;
	signal WX8315: std_logic; attribute dont_touch of WX8315: signal is true;
	signal WX8316: std_logic; attribute dont_touch of WX8316: signal is true;
	signal WX8317: std_logic; attribute dont_touch of WX8317: signal is true;
	signal WX8318: std_logic; attribute dont_touch of WX8318: signal is true;
	signal WX8319: std_logic; attribute dont_touch of WX8319: signal is true;
	signal WX8320: std_logic; attribute dont_touch of WX8320: signal is true;
	signal WX8321: std_logic; attribute dont_touch of WX8321: signal is true;
	signal WX8322: std_logic; attribute dont_touch of WX8322: signal is true;
	signal WX8323: std_logic; attribute dont_touch of WX8323: signal is true;
	signal WX8324: std_logic; attribute dont_touch of WX8324: signal is true;
	signal WX8325: std_logic; attribute dont_touch of WX8325: signal is true;
	signal WX8326: std_logic; attribute dont_touch of WX8326: signal is true;
	signal WX8327: std_logic; attribute dont_touch of WX8327: signal is true;
	signal WX8328: std_logic; attribute dont_touch of WX8328: signal is true;
	signal WX8329: std_logic; attribute dont_touch of WX8329: signal is true;
	signal WX8330: std_logic; attribute dont_touch of WX8330: signal is true;
	signal WX8331: std_logic; attribute dont_touch of WX8331: signal is true;
	signal WX8332: std_logic; attribute dont_touch of WX8332: signal is true;
	signal WX8333: std_logic; attribute dont_touch of WX8333: signal is true;
	signal WX8334: std_logic; attribute dont_touch of WX8334: signal is true;
	signal WX8335: std_logic; attribute dont_touch of WX8335: signal is true;
	signal WX8336: std_logic; attribute dont_touch of WX8336: signal is true;
	signal WX8337: std_logic; attribute dont_touch of WX8337: signal is true;
	signal WX8338: std_logic; attribute dont_touch of WX8338: signal is true;
	signal WX8339: std_logic; attribute dont_touch of WX8339: signal is true;
	signal WX8340: std_logic; attribute dont_touch of WX8340: signal is true;
	signal WX8341: std_logic; attribute dont_touch of WX8341: signal is true;
	signal WX8342: std_logic; attribute dont_touch of WX8342: signal is true;
	signal WX8343: std_logic; attribute dont_touch of WX8343: signal is true;
	signal WX8344: std_logic; attribute dont_touch of WX8344: signal is true;
	signal WX8345: std_logic; attribute dont_touch of WX8345: signal is true;
	signal WX8346: std_logic; attribute dont_touch of WX8346: signal is true;
	signal WX8347: std_logic; attribute dont_touch of WX8347: signal is true;
	signal WX8348: std_logic; attribute dont_touch of WX8348: signal is true;
	signal WX8349: std_logic; attribute dont_touch of WX8349: signal is true;
	signal WX8350: std_logic; attribute dont_touch of WX8350: signal is true;
	signal WX8351: std_logic; attribute dont_touch of WX8351: signal is true;
	signal WX8352: std_logic; attribute dont_touch of WX8352: signal is true;
	signal WX8353: std_logic; attribute dont_touch of WX8353: signal is true;
	signal WX8354: std_logic; attribute dont_touch of WX8354: signal is true;
	signal WX8355: std_logic; attribute dont_touch of WX8355: signal is true;
	signal WX8356: std_logic; attribute dont_touch of WX8356: signal is true;
	signal WX8357: std_logic; attribute dont_touch of WX8357: signal is true;
	signal WX8358: std_logic; attribute dont_touch of WX8358: signal is true;
	signal WX8359: std_logic; attribute dont_touch of WX8359: signal is true;
	signal WX8360: std_logic; attribute dont_touch of WX8360: signal is true;
	signal WX8361: std_logic; attribute dont_touch of WX8361: signal is true;
	signal WX8362: std_logic; attribute dont_touch of WX8362: signal is true;
	signal WX8363: std_logic; attribute dont_touch of WX8363: signal is true;
	signal WX8364: std_logic; attribute dont_touch of WX8364: signal is true;
	signal WX8365: std_logic; attribute dont_touch of WX8365: signal is true;
	signal WX8366: std_logic; attribute dont_touch of WX8366: signal is true;
	signal WX8367: std_logic; attribute dont_touch of WX8367: signal is true;
	signal WX8368: std_logic; attribute dont_touch of WX8368: signal is true;
	signal WX8369: std_logic; attribute dont_touch of WX8369: signal is true;
	signal WX8370: std_logic; attribute dont_touch of WX8370: signal is true;
	signal WX8371: std_logic; attribute dont_touch of WX8371: signal is true;
	signal WX8372: std_logic; attribute dont_touch of WX8372: signal is true;
	signal WX8373: std_logic; attribute dont_touch of WX8373: signal is true;
	signal WX8374: std_logic; attribute dont_touch of WX8374: signal is true;
	signal WX8375: std_logic; attribute dont_touch of WX8375: signal is true;
	signal WX8376: std_logic; attribute dont_touch of WX8376: signal is true;
	signal WX8377: std_logic; attribute dont_touch of WX8377: signal is true;
	signal WX8378: std_logic; attribute dont_touch of WX8378: signal is true;
	signal WX8379: std_logic; attribute dont_touch of WX8379: signal is true;
	signal WX8380: std_logic; attribute dont_touch of WX8380: signal is true;
	signal WX8381: std_logic; attribute dont_touch of WX8381: signal is true;
	signal WX8382: std_logic; attribute dont_touch of WX8382: signal is true;
	signal WX8383: std_logic; attribute dont_touch of WX8383: signal is true;
	signal WX8384: std_logic; attribute dont_touch of WX8384: signal is true;
	signal WX8385: std_logic; attribute dont_touch of WX8385: signal is true;
	signal WX8386: std_logic; attribute dont_touch of WX8386: signal is true;
	signal WX8387: std_logic; attribute dont_touch of WX8387: signal is true;
	signal WX8388: std_logic; attribute dont_touch of WX8388: signal is true;
	signal WX8389: std_logic; attribute dont_touch of WX8389: signal is true;
	signal WX8390: std_logic; attribute dont_touch of WX8390: signal is true;
	signal WX8391: std_logic; attribute dont_touch of WX8391: signal is true;
	signal WX8392: std_logic; attribute dont_touch of WX8392: signal is true;
	signal WX8393: std_logic; attribute dont_touch of WX8393: signal is true;
	signal WX8394: std_logic; attribute dont_touch of WX8394: signal is true;
	signal WX8395: std_logic; attribute dont_touch of WX8395: signal is true;
	signal WX8396: std_logic; attribute dont_touch of WX8396: signal is true;
	signal WX8397: std_logic; attribute dont_touch of WX8397: signal is true;
	signal WX8398: std_logic; attribute dont_touch of WX8398: signal is true;
	signal WX8399: std_logic; attribute dont_touch of WX8399: signal is true;
	signal WX8400: std_logic; attribute dont_touch of WX8400: signal is true;
	signal WX8401: std_logic; attribute dont_touch of WX8401: signal is true;
	signal WX8402: std_logic; attribute dont_touch of WX8402: signal is true;
	signal WX8403: std_logic; attribute dont_touch of WX8403: signal is true;
	signal WX8404: std_logic; attribute dont_touch of WX8404: signal is true;
	signal WX8405: std_logic; attribute dont_touch of WX8405: signal is true;
	signal WX8406: std_logic; attribute dont_touch of WX8406: signal is true;
	signal WX8407: std_logic; attribute dont_touch of WX8407: signal is true;
	signal WX8408: std_logic; attribute dont_touch of WX8408: signal is true;
	signal WX8409: std_logic; attribute dont_touch of WX8409: signal is true;
	signal WX8410: std_logic; attribute dont_touch of WX8410: signal is true;
	signal WX8411: std_logic; attribute dont_touch of WX8411: signal is true;
	signal WX8412: std_logic; attribute dont_touch of WX8412: signal is true;
	signal WX8413: std_logic; attribute dont_touch of WX8413: signal is true;
	signal WX8414: std_logic; attribute dont_touch of WX8414: signal is true;
	signal WX8415: std_logic; attribute dont_touch of WX8415: signal is true;
	signal WX8416: std_logic; attribute dont_touch of WX8416: signal is true;
	signal WX8417: std_logic; attribute dont_touch of WX8417: signal is true;
	signal WX8418: std_logic; attribute dont_touch of WX8418: signal is true;
	signal WX8419: std_logic; attribute dont_touch of WX8419: signal is true;
	signal WX8420: std_logic; attribute dont_touch of WX8420: signal is true;
	signal WX8421: std_logic; attribute dont_touch of WX8421: signal is true;
	signal WX8422: std_logic; attribute dont_touch of WX8422: signal is true;
	signal WX8423: std_logic; attribute dont_touch of WX8423: signal is true;
	signal WX8424: std_logic; attribute dont_touch of WX8424: signal is true;
	signal WX8425: std_logic; attribute dont_touch of WX8425: signal is true;
	signal WX8426: std_logic; attribute dont_touch of WX8426: signal is true;
	signal WX8427: std_logic; attribute dont_touch of WX8427: signal is true;
	signal WX8428: std_logic; attribute dont_touch of WX8428: signal is true;
	signal WX8429: std_logic; attribute dont_touch of WX8429: signal is true;
	signal WX8430: std_logic; attribute dont_touch of WX8430: signal is true;
	signal WX8431: std_logic; attribute dont_touch of WX8431: signal is true;
	signal WX8432: std_logic; attribute dont_touch of WX8432: signal is true;
	signal WX8433: std_logic; attribute dont_touch of WX8433: signal is true;
	signal WX8434: std_logic; attribute dont_touch of WX8434: signal is true;
	signal WX8435: std_logic; attribute dont_touch of WX8435: signal is true;
	signal WX8436: std_logic; attribute dont_touch of WX8436: signal is true;
	signal WX8437: std_logic; attribute dont_touch of WX8437: signal is true;
	signal WX8438: std_logic; attribute dont_touch of WX8438: signal is true;
	signal WX8439: std_logic; attribute dont_touch of WX8439: signal is true;
	signal WX8440: std_logic; attribute dont_touch of WX8440: signal is true;
	signal WX8441: std_logic; attribute dont_touch of WX8441: signal is true;
	signal WX8442: std_logic; attribute dont_touch of WX8442: signal is true;
	signal WX8443: std_logic; attribute dont_touch of WX8443: signal is true;
	signal WX8444: std_logic; attribute dont_touch of WX8444: signal is true;
	signal WX8445: std_logic; attribute dont_touch of WX8445: signal is true;
	signal WX8446: std_logic; attribute dont_touch of WX8446: signal is true;
	signal WX8447: std_logic; attribute dont_touch of WX8447: signal is true;
	signal WX8448: std_logic; attribute dont_touch of WX8448: signal is true;
	signal WX8449: std_logic; attribute dont_touch of WX8449: signal is true;
	signal WX8450: std_logic; attribute dont_touch of WX8450: signal is true;
	signal WX8451: std_logic; attribute dont_touch of WX8451: signal is true;
	signal WX8452: std_logic; attribute dont_touch of WX8452: signal is true;
	signal WX8453: std_logic; attribute dont_touch of WX8453: signal is true;
	signal WX8454: std_logic; attribute dont_touch of WX8454: signal is true;
	signal WX8455: std_logic; attribute dont_touch of WX8455: signal is true;
	signal WX8456: std_logic; attribute dont_touch of WX8456: signal is true;
	signal WX8457: std_logic; attribute dont_touch of WX8457: signal is true;
	signal WX8458: std_logic; attribute dont_touch of WX8458: signal is true;
	signal WX8459: std_logic; attribute dont_touch of WX8459: signal is true;
	signal WX8460: std_logic; attribute dont_touch of WX8460: signal is true;
	signal WX8461: std_logic; attribute dont_touch of WX8461: signal is true;
	signal WX8462: std_logic; attribute dont_touch of WX8462: signal is true;
	signal WX8463: std_logic; attribute dont_touch of WX8463: signal is true;
	signal WX8464: std_logic; attribute dont_touch of WX8464: signal is true;
	signal WX8465: std_logic; attribute dont_touch of WX8465: signal is true;
	signal WX8466: std_logic; attribute dont_touch of WX8466: signal is true;
	signal WX8467: std_logic; attribute dont_touch of WX8467: signal is true;
	signal WX8468: std_logic; attribute dont_touch of WX8468: signal is true;
	signal WX8469: std_logic; attribute dont_touch of WX8469: signal is true;
	signal WX8470: std_logic; attribute dont_touch of WX8470: signal is true;
	signal WX8471: std_logic; attribute dont_touch of WX8471: signal is true;
	signal WX8472: std_logic; attribute dont_touch of WX8472: signal is true;
	signal WX8473: std_logic; attribute dont_touch of WX8473: signal is true;
	signal WX8474: std_logic; attribute dont_touch of WX8474: signal is true;
	signal WX8475: std_logic; attribute dont_touch of WX8475: signal is true;
	signal WX8476: std_logic; attribute dont_touch of WX8476: signal is true;
	signal WX8477: std_logic; attribute dont_touch of WX8477: signal is true;
	signal WX8478: std_logic; attribute dont_touch of WX8478: signal is true;
	signal WX8479: std_logic; attribute dont_touch of WX8479: signal is true;
	signal WX8480: std_logic; attribute dont_touch of WX8480: signal is true;
	signal WX8481: std_logic; attribute dont_touch of WX8481: signal is true;
	signal WX8482: std_logic; attribute dont_touch of WX8482: signal is true;
	signal WX8483: std_logic; attribute dont_touch of WX8483: signal is true;
	signal WX8484: std_logic; attribute dont_touch of WX8484: signal is true;
	signal WX8485: std_logic; attribute dont_touch of WX8485: signal is true;
	signal WX8486: std_logic; attribute dont_touch of WX8486: signal is true;
	signal WX8487: std_logic; attribute dont_touch of WX8487: signal is true;
	signal WX8488: std_logic; attribute dont_touch of WX8488: signal is true;
	signal WX8489: std_logic; attribute dont_touch of WX8489: signal is true;
	signal WX8490: std_logic; attribute dont_touch of WX8490: signal is true;
	signal WX8491: std_logic; attribute dont_touch of WX8491: signal is true;
	signal WX8492: std_logic; attribute dont_touch of WX8492: signal is true;
	signal WX8493: std_logic; attribute dont_touch of WX8493: signal is true;
	signal WX8494: std_logic; attribute dont_touch of WX8494: signal is true;
	signal WX8495: std_logic; attribute dont_touch of WX8495: signal is true;
	signal WX8496: std_logic; attribute dont_touch of WX8496: signal is true;
	signal WX8497: std_logic; attribute dont_touch of WX8497: signal is true;
	signal WX8498: std_logic; attribute dont_touch of WX8498: signal is true;
	signal WX8499: std_logic; attribute dont_touch of WX8499: signal is true;
	signal WX8500: std_logic; attribute dont_touch of WX8500: signal is true;
	signal WX8501: std_logic; attribute dont_touch of WX8501: signal is true;
	signal WX8502: std_logic; attribute dont_touch of WX8502: signal is true;
	signal WX8503: std_logic; attribute dont_touch of WX8503: signal is true;
	signal WX8504: std_logic; attribute dont_touch of WX8504: signal is true;
	signal WX8505: std_logic; attribute dont_touch of WX8505: signal is true;
	signal WX8506: std_logic; attribute dont_touch of WX8506: signal is true;
	signal WX8507: std_logic; attribute dont_touch of WX8507: signal is true;
	signal WX8508: std_logic; attribute dont_touch of WX8508: signal is true;
	signal WX8509: std_logic; attribute dont_touch of WX8509: signal is true;
	signal WX8510: std_logic; attribute dont_touch of WX8510: signal is true;
	signal WX8511: std_logic; attribute dont_touch of WX8511: signal is true;
	signal WX8512: std_logic; attribute dont_touch of WX8512: signal is true;
	signal WX8513: std_logic; attribute dont_touch of WX8513: signal is true;
	signal WX8514: std_logic; attribute dont_touch of WX8514: signal is true;
	signal WX8515: std_logic; attribute dont_touch of WX8515: signal is true;
	signal WX8516: std_logic; attribute dont_touch of WX8516: signal is true;
	signal WX8517: std_logic; attribute dont_touch of WX8517: signal is true;
	signal WX8518: std_logic; attribute dont_touch of WX8518: signal is true;
	signal WX8519: std_logic; attribute dont_touch of WX8519: signal is true;
	signal WX8520: std_logic; attribute dont_touch of WX8520: signal is true;
	signal WX8521: std_logic; attribute dont_touch of WX8521: signal is true;
	signal WX8522: std_logic; attribute dont_touch of WX8522: signal is true;
	signal WX8523: std_logic; attribute dont_touch of WX8523: signal is true;
	signal WX8524: std_logic; attribute dont_touch of WX8524: signal is true;
	signal WX8525: std_logic; attribute dont_touch of WX8525: signal is true;
	signal WX8526: std_logic; attribute dont_touch of WX8526: signal is true;
	signal WX8527: std_logic; attribute dont_touch of WX8527: signal is true;
	signal WX8528: std_logic; attribute dont_touch of WX8528: signal is true;
	signal WX8529: std_logic; attribute dont_touch of WX8529: signal is true;
	signal WX8530: std_logic; attribute dont_touch of WX8530: signal is true;
	signal WX8531: std_logic; attribute dont_touch of WX8531: signal is true;
	signal WX8532: std_logic; attribute dont_touch of WX8532: signal is true;
	signal WX8533: std_logic; attribute dont_touch of WX8533: signal is true;
	signal WX8534: std_logic; attribute dont_touch of WX8534: signal is true;
	signal WX8535: std_logic; attribute dont_touch of WX8535: signal is true;
	signal WX8536: std_logic; attribute dont_touch of WX8536: signal is true;
	signal WX8537: std_logic; attribute dont_touch of WX8537: signal is true;
	signal WX8538: std_logic; attribute dont_touch of WX8538: signal is true;
	signal WX8539: std_logic; attribute dont_touch of WX8539: signal is true;
	signal WX8540: std_logic; attribute dont_touch of WX8540: signal is true;
	signal WX8541: std_logic; attribute dont_touch of WX8541: signal is true;
	signal WX8542: std_logic; attribute dont_touch of WX8542: signal is true;
	signal WX8543: std_logic; attribute dont_touch of WX8543: signal is true;
	signal WX8544: std_logic; attribute dont_touch of WX8544: signal is true;
	signal WX8545: std_logic; attribute dont_touch of WX8545: signal is true;
	signal WX8546: std_logic; attribute dont_touch of WX8546: signal is true;
	signal WX8547: std_logic; attribute dont_touch of WX8547: signal is true;
	signal WX8548: std_logic; attribute dont_touch of WX8548: signal is true;
	signal WX8549: std_logic; attribute dont_touch of WX8549: signal is true;
	signal WX8550: std_logic; attribute dont_touch of WX8550: signal is true;
	signal WX8551: std_logic; attribute dont_touch of WX8551: signal is true;
	signal WX8552: std_logic; attribute dont_touch of WX8552: signal is true;
	signal WX8553: std_logic; attribute dont_touch of WX8553: signal is true;
	signal WX8554: std_logic; attribute dont_touch of WX8554: signal is true;
	signal WX8555: std_logic; attribute dont_touch of WX8555: signal is true;
	signal WX8556: std_logic; attribute dont_touch of WX8556: signal is true;
	signal WX8557: std_logic; attribute dont_touch of WX8557: signal is true;
	signal WX8558: std_logic; attribute dont_touch of WX8558: signal is true;
	signal WX8559: std_logic; attribute dont_touch of WX8559: signal is true;
	signal WX8560: std_logic; attribute dont_touch of WX8560: signal is true;
	signal WX8561: std_logic; attribute dont_touch of WX8561: signal is true;
	signal WX8562: std_logic; attribute dont_touch of WX8562: signal is true;
	signal WX8563: std_logic; attribute dont_touch of WX8563: signal is true;
	signal WX8564: std_logic; attribute dont_touch of WX8564: signal is true;
	signal WX8565: std_logic; attribute dont_touch of WX8565: signal is true;
	signal WX8566: std_logic; attribute dont_touch of WX8566: signal is true;
	signal WX8567: std_logic; attribute dont_touch of WX8567: signal is true;
	signal WX8568: std_logic; attribute dont_touch of WX8568: signal is true;
	signal WX8569: std_logic; attribute dont_touch of WX8569: signal is true;
	signal WX8570: std_logic; attribute dont_touch of WX8570: signal is true;
	signal WX8571: std_logic; attribute dont_touch of WX8571: signal is true;
	signal WX8572: std_logic; attribute dont_touch of WX8572: signal is true;
	signal WX8573: std_logic; attribute dont_touch of WX8573: signal is true;
	signal WX8574: std_logic; attribute dont_touch of WX8574: signal is true;
	signal WX8575: std_logic; attribute dont_touch of WX8575: signal is true;
	signal WX8576: std_logic; attribute dont_touch of WX8576: signal is true;
	signal WX8577: std_logic; attribute dont_touch of WX8577: signal is true;
	signal WX8578: std_logic; attribute dont_touch of WX8578: signal is true;
	signal WX8579: std_logic; attribute dont_touch of WX8579: signal is true;
	signal WX8580: std_logic; attribute dont_touch of WX8580: signal is true;
	signal WX8581: std_logic; attribute dont_touch of WX8581: signal is true;
	signal WX8582: std_logic; attribute dont_touch of WX8582: signal is true;
	signal WX8583: std_logic; attribute dont_touch of WX8583: signal is true;
	signal WX8584: std_logic; attribute dont_touch of WX8584: signal is true;
	signal WX8585: std_logic; attribute dont_touch of WX8585: signal is true;
	signal WX8586: std_logic; attribute dont_touch of WX8586: signal is true;
	signal WX8587: std_logic; attribute dont_touch of WX8587: signal is true;
	signal WX8588: std_logic; attribute dont_touch of WX8588: signal is true;
	signal WX8589: std_logic; attribute dont_touch of WX8589: signal is true;
	signal WX8590: std_logic; attribute dont_touch of WX8590: signal is true;
	signal WX8591: std_logic; attribute dont_touch of WX8591: signal is true;
	signal WX8592: std_logic; attribute dont_touch of WX8592: signal is true;
	signal WX8593: std_logic; attribute dont_touch of WX8593: signal is true;
	signal WX8594: std_logic; attribute dont_touch of WX8594: signal is true;
	signal WX8595: std_logic; attribute dont_touch of WX8595: signal is true;
	signal WX8596: std_logic; attribute dont_touch of WX8596: signal is true;
	signal WX8597: std_logic; attribute dont_touch of WX8597: signal is true;
	signal WX8598: std_logic; attribute dont_touch of WX8598: signal is true;
	signal WX8599: std_logic; attribute dont_touch of WX8599: signal is true;
	signal WX8600: std_logic; attribute dont_touch of WX8600: signal is true;
	signal WX8601: std_logic; attribute dont_touch of WX8601: signal is true;
	signal WX8602: std_logic; attribute dont_touch of WX8602: signal is true;
	signal WX8603: std_logic; attribute dont_touch of WX8603: signal is true;
	signal WX8604: std_logic; attribute dont_touch of WX8604: signal is true;
	signal WX8605: std_logic; attribute dont_touch of WX8605: signal is true;
	signal WX8606: std_logic; attribute dont_touch of WX8606: signal is true;
	signal WX8607: std_logic; attribute dont_touch of WX8607: signal is true;
	signal WX8608: std_logic; attribute dont_touch of WX8608: signal is true;
	signal WX8609: std_logic; attribute dont_touch of WX8609: signal is true;
	signal WX8610: std_logic; attribute dont_touch of WX8610: signal is true;
	signal WX8611: std_logic; attribute dont_touch of WX8611: signal is true;
	signal WX8612: std_logic; attribute dont_touch of WX8612: signal is true;
	signal WX8613: std_logic; attribute dont_touch of WX8613: signal is true;
	signal WX8614: std_logic; attribute dont_touch of WX8614: signal is true;
	signal WX8615: std_logic; attribute dont_touch of WX8615: signal is true;
	signal WX8616: std_logic; attribute dont_touch of WX8616: signal is true;
	signal WX8617: std_logic; attribute dont_touch of WX8617: signal is true;
	signal WX8618: std_logic; attribute dont_touch of WX8618: signal is true;
	signal WX8619: std_logic; attribute dont_touch of WX8619: signal is true;
	signal WX8620: std_logic; attribute dont_touch of WX8620: signal is true;
	signal WX8621: std_logic; attribute dont_touch of WX8621: signal is true;
	signal WX8622: std_logic; attribute dont_touch of WX8622: signal is true;
	signal WX8623: std_logic; attribute dont_touch of WX8623: signal is true;
	signal WX8624: std_logic; attribute dont_touch of WX8624: signal is true;
	signal WX8625: std_logic; attribute dont_touch of WX8625: signal is true;
	signal WX8626: std_logic; attribute dont_touch of WX8626: signal is true;
	signal WX8627: std_logic; attribute dont_touch of WX8627: signal is true;
	signal WX8628: std_logic; attribute dont_touch of WX8628: signal is true;
	signal WX8629: std_logic; attribute dont_touch of WX8629: signal is true;
	signal WX8630: std_logic; attribute dont_touch of WX8630: signal is true;
	signal WX8631: std_logic; attribute dont_touch of WX8631: signal is true;
	signal WX8632: std_logic; attribute dont_touch of WX8632: signal is true;
	signal WX8633: std_logic; attribute dont_touch of WX8633: signal is true;
	signal WX8634: std_logic; attribute dont_touch of WX8634: signal is true;
	signal WX8635: std_logic; attribute dont_touch of WX8635: signal is true;
	signal WX8636: std_logic; attribute dont_touch of WX8636: signal is true;
	signal WX8637: std_logic; attribute dont_touch of WX8637: signal is true;
	signal WX8638: std_logic; attribute dont_touch of WX8638: signal is true;
	signal WX8639: std_logic; attribute dont_touch of WX8639: signal is true;
	signal WX8640: std_logic; attribute dont_touch of WX8640: signal is true;
	signal WX8641: std_logic; attribute dont_touch of WX8641: signal is true;
	signal WX8642: std_logic; attribute dont_touch of WX8642: signal is true;
	signal WX8643: std_logic; attribute dont_touch of WX8643: signal is true;
	signal WX8644: std_logic; attribute dont_touch of WX8644: signal is true;
	signal WX8645: std_logic; attribute dont_touch of WX8645: signal is true;
	signal WX8646: std_logic; attribute dont_touch of WX8646: signal is true;
	signal WX8647: std_logic; attribute dont_touch of WX8647: signal is true;
	signal WX8648: std_logic; attribute dont_touch of WX8648: signal is true;
	signal WX8649: std_logic; attribute dont_touch of WX8649: signal is true;
	signal WX8650: std_logic; attribute dont_touch of WX8650: signal is true;
	signal WX8651: std_logic; attribute dont_touch of WX8651: signal is true;
	signal WX8652: std_logic; attribute dont_touch of WX8652: signal is true;
	signal WX8653: std_logic; attribute dont_touch of WX8653: signal is true;
	signal WX8654: std_logic; attribute dont_touch of WX8654: signal is true;
	signal WX8655: std_logic; attribute dont_touch of WX8655: signal is true;
	signal WX8656: std_logic; attribute dont_touch of WX8656: signal is true;
	signal WX8657: std_logic; attribute dont_touch of WX8657: signal is true;
	signal WX8658: std_logic; attribute dont_touch of WX8658: signal is true;
	signal WX8659: std_logic; attribute dont_touch of WX8659: signal is true;
	signal WX8660: std_logic; attribute dont_touch of WX8660: signal is true;
	signal WX8661: std_logic; attribute dont_touch of WX8661: signal is true;
	signal WX8662: std_logic; attribute dont_touch of WX8662: signal is true;
	signal WX8663: std_logic; attribute dont_touch of WX8663: signal is true;
	signal WX8664: std_logic; attribute dont_touch of WX8664: signal is true;
	signal WX8665: std_logic; attribute dont_touch of WX8665: signal is true;
	signal WX8666: std_logic; attribute dont_touch of WX8666: signal is true;
	signal WX8667: std_logic; attribute dont_touch of WX8667: signal is true;
	signal WX8668: std_logic; attribute dont_touch of WX8668: signal is true;
	signal WX8669: std_logic; attribute dont_touch of WX8669: signal is true;
	signal WX8670: std_logic; attribute dont_touch of WX8670: signal is true;
	signal WX8671: std_logic; attribute dont_touch of WX8671: signal is true;
	signal WX8672: std_logic; attribute dont_touch of WX8672: signal is true;
	signal WX8673: std_logic; attribute dont_touch of WX8673: signal is true;
	signal WX8674: std_logic; attribute dont_touch of WX8674: signal is true;
	signal WX8675: std_logic; attribute dont_touch of WX8675: signal is true;
	signal WX8676: std_logic; attribute dont_touch of WX8676: signal is true;
	signal WX8677: std_logic; attribute dont_touch of WX8677: signal is true;
	signal WX8678: std_logic; attribute dont_touch of WX8678: signal is true;
	signal WX8679: std_logic; attribute dont_touch of WX8679: signal is true;
	signal WX8680: std_logic; attribute dont_touch of WX8680: signal is true;
	signal WX8681: std_logic; attribute dont_touch of WX8681: signal is true;
	signal WX8682: std_logic; attribute dont_touch of WX8682: signal is true;
	signal WX8683: std_logic; attribute dont_touch of WX8683: signal is true;
	signal WX8684: std_logic; attribute dont_touch of WX8684: signal is true;
	signal WX8685: std_logic; attribute dont_touch of WX8685: signal is true;
	signal WX8686: std_logic; attribute dont_touch of WX8686: signal is true;
	signal WX8687: std_logic; attribute dont_touch of WX8687: signal is true;
	signal WX8688: std_logic; attribute dont_touch of WX8688: signal is true;
	signal WX8689: std_logic; attribute dont_touch of WX8689: signal is true;
	signal WX8690: std_logic; attribute dont_touch of WX8690: signal is true;
	signal WX8691: std_logic; attribute dont_touch of WX8691: signal is true;
	signal WX8692: std_logic; attribute dont_touch of WX8692: signal is true;
	signal WX8693: std_logic; attribute dont_touch of WX8693: signal is true;
	signal WX8694: std_logic; attribute dont_touch of WX8694: signal is true;
	signal WX8695: std_logic; attribute dont_touch of WX8695: signal is true;
	signal WX8696: std_logic; attribute dont_touch of WX8696: signal is true;
	signal WX8697: std_logic; attribute dont_touch of WX8697: signal is true;
	signal WX8698: std_logic; attribute dont_touch of WX8698: signal is true;
	signal WX8699: std_logic; attribute dont_touch of WX8699: signal is true;
	signal WX8700: std_logic; attribute dont_touch of WX8700: signal is true;
	signal WX8701: std_logic; attribute dont_touch of WX8701: signal is true;
	signal WX8702: std_logic; attribute dont_touch of WX8702: signal is true;
	signal WX8703: std_logic; attribute dont_touch of WX8703: signal is true;
	signal WX8704: std_logic; attribute dont_touch of WX8704: signal is true;
	signal WX8705: std_logic; attribute dont_touch of WX8705: signal is true;
	signal WX8706: std_logic; attribute dont_touch of WX8706: signal is true;
	signal WX8707: std_logic; attribute dont_touch of WX8707: signal is true;
	signal WX8708: std_logic; attribute dont_touch of WX8708: signal is true;
	signal WX8709: std_logic; attribute dont_touch of WX8709: signal is true;
	signal WX8710: std_logic; attribute dont_touch of WX8710: signal is true;
	signal WX8711: std_logic; attribute dont_touch of WX8711: signal is true;
	signal WX8712: std_logic; attribute dont_touch of WX8712: signal is true;
	signal WX8713: std_logic; attribute dont_touch of WX8713: signal is true;
	signal WX8714: std_logic; attribute dont_touch of WX8714: signal is true;
	signal WX8715: std_logic; attribute dont_touch of WX8715: signal is true;
	signal WX8716: std_logic; attribute dont_touch of WX8716: signal is true;
	signal WX8717: std_logic; attribute dont_touch of WX8717: signal is true;
	signal WX8718: std_logic; attribute dont_touch of WX8718: signal is true;
	signal WX8719: std_logic; attribute dont_touch of WX8719: signal is true;
	signal WX8720: std_logic; attribute dont_touch of WX8720: signal is true;
	signal WX8721: std_logic; attribute dont_touch of WX8721: signal is true;
	signal WX8722: std_logic; attribute dont_touch of WX8722: signal is true;
	signal WX8723: std_logic; attribute dont_touch of WX8723: signal is true;
	signal WX8724: std_logic; attribute dont_touch of WX8724: signal is true;
	signal WX8725: std_logic; attribute dont_touch of WX8725: signal is true;
	signal WX8726: std_logic; attribute dont_touch of WX8726: signal is true;
	signal WX8727: std_logic; attribute dont_touch of WX8727: signal is true;
	signal WX8728: std_logic; attribute dont_touch of WX8728: signal is true;
	signal WX8729: std_logic; attribute dont_touch of WX8729: signal is true;
	signal WX8730: std_logic; attribute dont_touch of WX8730: signal is true;
	signal WX8731: std_logic; attribute dont_touch of WX8731: signal is true;
	signal WX8732: std_logic; attribute dont_touch of WX8732: signal is true;
	signal WX8733: std_logic; attribute dont_touch of WX8733: signal is true;
	signal WX8734: std_logic; attribute dont_touch of WX8734: signal is true;
	signal WX8735: std_logic; attribute dont_touch of WX8735: signal is true;
	signal WX8736: std_logic; attribute dont_touch of WX8736: signal is true;
	signal WX8737: std_logic; attribute dont_touch of WX8737: signal is true;
	signal WX8738: std_logic; attribute dont_touch of WX8738: signal is true;
	signal WX8739: std_logic; attribute dont_touch of WX8739: signal is true;
	signal WX8740: std_logic; attribute dont_touch of WX8740: signal is true;
	signal WX8741: std_logic; attribute dont_touch of WX8741: signal is true;
	signal WX8742: std_logic; attribute dont_touch of WX8742: signal is true;
	signal WX8743: std_logic; attribute dont_touch of WX8743: signal is true;
	signal WX8744: std_logic; attribute dont_touch of WX8744: signal is true;
	signal WX8745: std_logic; attribute dont_touch of WX8745: signal is true;
	signal WX8746: std_logic; attribute dont_touch of WX8746: signal is true;
	signal WX8747: std_logic; attribute dont_touch of WX8747: signal is true;
	signal WX8748: std_logic; attribute dont_touch of WX8748: signal is true;
	signal WX8749: std_logic; attribute dont_touch of WX8749: signal is true;
	signal WX8750: std_logic; attribute dont_touch of WX8750: signal is true;
	signal WX8751: std_logic; attribute dont_touch of WX8751: signal is true;
	signal WX8752: std_logic; attribute dont_touch of WX8752: signal is true;
	signal WX8753: std_logic; attribute dont_touch of WX8753: signal is true;
	signal WX8754: std_logic; attribute dont_touch of WX8754: signal is true;
	signal WX8755: std_logic; attribute dont_touch of WX8755: signal is true;
	signal WX8756: std_logic; attribute dont_touch of WX8756: signal is true;
	signal WX8757: std_logic; attribute dont_touch of WX8757: signal is true;
	signal WX8758: std_logic; attribute dont_touch of WX8758: signal is true;
	signal WX8759: std_logic; attribute dont_touch of WX8759: signal is true;
	signal WX8760: std_logic; attribute dont_touch of WX8760: signal is true;
	signal WX8761: std_logic; attribute dont_touch of WX8761: signal is true;
	signal WX8762: std_logic; attribute dont_touch of WX8762: signal is true;
	signal WX8763: std_logic; attribute dont_touch of WX8763: signal is true;
	signal WX8764: std_logic; attribute dont_touch of WX8764: signal is true;
	signal WX8765: std_logic; attribute dont_touch of WX8765: signal is true;
	signal WX8766: std_logic; attribute dont_touch of WX8766: signal is true;
	signal WX8767: std_logic; attribute dont_touch of WX8767: signal is true;
	signal WX8768: std_logic; attribute dont_touch of WX8768: signal is true;
	signal WX8769: std_logic; attribute dont_touch of WX8769: signal is true;
	signal WX8770: std_logic; attribute dont_touch of WX8770: signal is true;
	signal WX8771: std_logic; attribute dont_touch of WX8771: signal is true;
	signal WX8772: std_logic; attribute dont_touch of WX8772: signal is true;
	signal WX8773: std_logic; attribute dont_touch of WX8773: signal is true;
	signal WX8774: std_logic; attribute dont_touch of WX8774: signal is true;
	signal WX8775: std_logic; attribute dont_touch of WX8775: signal is true;
	signal WX8776: std_logic; attribute dont_touch of WX8776: signal is true;
	signal WX8777: std_logic; attribute dont_touch of WX8777: signal is true;
	signal WX8778: std_logic; attribute dont_touch of WX8778: signal is true;
	signal WX8779: std_logic; attribute dont_touch of WX8779: signal is true;
	signal WX8780: std_logic; attribute dont_touch of WX8780: signal is true;
	signal WX8781: std_logic; attribute dont_touch of WX8781: signal is true;
	signal WX8782: std_logic; attribute dont_touch of WX8782: signal is true;
	signal WX8783: std_logic; attribute dont_touch of WX8783: signal is true;
	signal WX8784: std_logic; attribute dont_touch of WX8784: signal is true;
	signal WX8785: std_logic; attribute dont_touch of WX8785: signal is true;
	signal WX8786: std_logic; attribute dont_touch of WX8786: signal is true;
	signal WX8787: std_logic; attribute dont_touch of WX8787: signal is true;
	signal WX8788: std_logic; attribute dont_touch of WX8788: signal is true;
	signal WX8789: std_logic; attribute dont_touch of WX8789: signal is true;
	signal WX8790: std_logic; attribute dont_touch of WX8790: signal is true;
	signal WX8791: std_logic; attribute dont_touch of WX8791: signal is true;
	signal WX8792: std_logic; attribute dont_touch of WX8792: signal is true;
	signal WX8793: std_logic; attribute dont_touch of WX8793: signal is true;
	signal WX8794: std_logic; attribute dont_touch of WX8794: signal is true;
	signal WX8795: std_logic; attribute dont_touch of WX8795: signal is true;
	signal WX8796: std_logic; attribute dont_touch of WX8796: signal is true;
	signal WX8797: std_logic; attribute dont_touch of WX8797: signal is true;
	signal WX8798: std_logic; attribute dont_touch of WX8798: signal is true;
	signal WX8799: std_logic; attribute dont_touch of WX8799: signal is true;
	signal WX8800: std_logic; attribute dont_touch of WX8800: signal is true;
	signal WX8801: std_logic; attribute dont_touch of WX8801: signal is true;
	signal WX8802: std_logic; attribute dont_touch of WX8802: signal is true;
	signal WX8803: std_logic; attribute dont_touch of WX8803: signal is true;
	signal WX8804: std_logic; attribute dont_touch of WX8804: signal is true;
	signal WX8805: std_logic; attribute dont_touch of WX8805: signal is true;
	signal WX8806: std_logic; attribute dont_touch of WX8806: signal is true;
	signal WX8807: std_logic; attribute dont_touch of WX8807: signal is true;
	signal WX8808: std_logic; attribute dont_touch of WX8808: signal is true;
	signal WX8809: std_logic; attribute dont_touch of WX8809: signal is true;
	signal WX8810: std_logic; attribute dont_touch of WX8810: signal is true;
	signal WX8811: std_logic; attribute dont_touch of WX8811: signal is true;
	signal WX8812: std_logic; attribute dont_touch of WX8812: signal is true;
	signal WX8813: std_logic; attribute dont_touch of WX8813: signal is true;
	signal WX8814: std_logic; attribute dont_touch of WX8814: signal is true;
	signal WX8815: std_logic; attribute dont_touch of WX8815: signal is true;
	signal WX8816: std_logic; attribute dont_touch of WX8816: signal is true;
	signal WX8817: std_logic; attribute dont_touch of WX8817: signal is true;
	signal WX8818: std_logic; attribute dont_touch of WX8818: signal is true;
	signal WX8819: std_logic; attribute dont_touch of WX8819: signal is true;
	signal WX8820: std_logic; attribute dont_touch of WX8820: signal is true;
	signal WX8821: std_logic; attribute dont_touch of WX8821: signal is true;
	signal WX8822: std_logic; attribute dont_touch of WX8822: signal is true;
	signal WX8823: std_logic; attribute dont_touch of WX8823: signal is true;
	signal WX8824: std_logic; attribute dont_touch of WX8824: signal is true;
	signal WX8825: std_logic; attribute dont_touch of WX8825: signal is true;
	signal WX8826: std_logic; attribute dont_touch of WX8826: signal is true;
	signal WX8827: std_logic; attribute dont_touch of WX8827: signal is true;
	signal WX8828: std_logic; attribute dont_touch of WX8828: signal is true;
	signal WX8829: std_logic; attribute dont_touch of WX8829: signal is true;
	signal WX8830: std_logic; attribute dont_touch of WX8830: signal is true;
	signal WX8831: std_logic; attribute dont_touch of WX8831: signal is true;
	signal WX8832: std_logic; attribute dont_touch of WX8832: signal is true;
	signal WX8833: std_logic; attribute dont_touch of WX8833: signal is true;
	signal WX8834: std_logic; attribute dont_touch of WX8834: signal is true;
	signal WX8835: std_logic; attribute dont_touch of WX8835: signal is true;
	signal WX8836: std_logic; attribute dont_touch of WX8836: signal is true;
	signal WX8837: std_logic; attribute dont_touch of WX8837: signal is true;
	signal WX8838: std_logic; attribute dont_touch of WX8838: signal is true;
	signal WX8839: std_logic; attribute dont_touch of WX8839: signal is true;
	signal WX8840: std_logic; attribute dont_touch of WX8840: signal is true;
	signal WX8841: std_logic; attribute dont_touch of WX8841: signal is true;
	signal WX8842: std_logic; attribute dont_touch of WX8842: signal is true;
	signal WX8843: std_logic; attribute dont_touch of WX8843: signal is true;
	signal WX8844: std_logic; attribute dont_touch of WX8844: signal is true;
	signal WX8845: std_logic; attribute dont_touch of WX8845: signal is true;
	signal WX8846: std_logic; attribute dont_touch of WX8846: signal is true;
	signal WX8847: std_logic; attribute dont_touch of WX8847: signal is true;
	signal WX8848: std_logic; attribute dont_touch of WX8848: signal is true;
	signal WX8849: std_logic; attribute dont_touch of WX8849: signal is true;
	signal WX8850: std_logic; attribute dont_touch of WX8850: signal is true;
	signal WX8851: std_logic; attribute dont_touch of WX8851: signal is true;
	signal WX8852: std_logic; attribute dont_touch of WX8852: signal is true;
	signal WX8853: std_logic; attribute dont_touch of WX8853: signal is true;
	signal WX8854: std_logic; attribute dont_touch of WX8854: signal is true;
	signal WX8855: std_logic; attribute dont_touch of WX8855: signal is true;
	signal WX8856: std_logic; attribute dont_touch of WX8856: signal is true;
	signal WX8857: std_logic; attribute dont_touch of WX8857: signal is true;
	signal WX8858: std_logic; attribute dont_touch of WX8858: signal is true;
	signal WX8859: std_logic; attribute dont_touch of WX8859: signal is true;
	signal WX8860: std_logic; attribute dont_touch of WX8860: signal is true;
	signal WX8861: std_logic; attribute dont_touch of WX8861: signal is true;
	signal WX8862: std_logic; attribute dont_touch of WX8862: signal is true;
	signal WX8863: std_logic; attribute dont_touch of WX8863: signal is true;
	signal WX8864: std_logic; attribute dont_touch of WX8864: signal is true;
	signal WX8865: std_logic; attribute dont_touch of WX8865: signal is true;
	signal WX8866: std_logic; attribute dont_touch of WX8866: signal is true;
	signal WX8867: std_logic; attribute dont_touch of WX8867: signal is true;
	signal WX8868: std_logic; attribute dont_touch of WX8868: signal is true;
	signal WX8869: std_logic; attribute dont_touch of WX8869: signal is true;
	signal WX8870: std_logic; attribute dont_touch of WX8870: signal is true;
	signal WX8871: std_logic; attribute dont_touch of WX8871: signal is true;
	signal WX8872: std_logic; attribute dont_touch of WX8872: signal is true;
	signal WX8873: std_logic; attribute dont_touch of WX8873: signal is true;
	signal WX8874: std_logic; attribute dont_touch of WX8874: signal is true;
	signal WX8875: std_logic; attribute dont_touch of WX8875: signal is true;
	signal WX8876: std_logic; attribute dont_touch of WX8876: signal is true;
	signal WX8877: std_logic; attribute dont_touch of WX8877: signal is true;
	signal WX8878: std_logic; attribute dont_touch of WX8878: signal is true;
	signal WX8879: std_logic; attribute dont_touch of WX8879: signal is true;
	signal WX8880: std_logic; attribute dont_touch of WX8880: signal is true;
	signal WX8881: std_logic; attribute dont_touch of WX8881: signal is true;
	signal WX8882: std_logic; attribute dont_touch of WX8882: signal is true;
	signal WX8883: std_logic; attribute dont_touch of WX8883: signal is true;
	signal WX8884: std_logic; attribute dont_touch of WX8884: signal is true;
	signal WX8885: std_logic; attribute dont_touch of WX8885: signal is true;
	signal WX8886: std_logic; attribute dont_touch of WX8886: signal is true;
	signal WX8887: std_logic; attribute dont_touch of WX8887: signal is true;
	signal WX8888: std_logic; attribute dont_touch of WX8888: signal is true;
	signal WX8889: std_logic; attribute dont_touch of WX8889: signal is true;
	signal WX8890: std_logic; attribute dont_touch of WX8890: signal is true;
	signal WX8891: std_logic; attribute dont_touch of WX8891: signal is true;
	signal WX8892: std_logic; attribute dont_touch of WX8892: signal is true;
	signal WX8893: std_logic; attribute dont_touch of WX8893: signal is true;
	signal WX8894: std_logic; attribute dont_touch of WX8894: signal is true;
	signal WX8895: std_logic; attribute dont_touch of WX8895: signal is true;
	signal WX8896: std_logic; attribute dont_touch of WX8896: signal is true;
	signal WX8897: std_logic; attribute dont_touch of WX8897: signal is true;
	signal WX8898: std_logic; attribute dont_touch of WX8898: signal is true;
	signal WX8899: std_logic; attribute dont_touch of WX8899: signal is true;
	signal WX8900: std_logic; attribute dont_touch of WX8900: signal is true;
	signal WX8901: std_logic; attribute dont_touch of WX8901: signal is true;
	signal WX8902: std_logic; attribute dont_touch of WX8902: signal is true;
	signal WX8903: std_logic; attribute dont_touch of WX8903: signal is true;
	signal WX8904: std_logic; attribute dont_touch of WX8904: signal is true;
	signal WX8905: std_logic; attribute dont_touch of WX8905: signal is true;
	signal WX8906: std_logic; attribute dont_touch of WX8906: signal is true;
	signal WX8907: std_logic; attribute dont_touch of WX8907: signal is true;
	signal WX8908: std_logic; attribute dont_touch of WX8908: signal is true;
	signal WX8909: std_logic; attribute dont_touch of WX8909: signal is true;
	signal WX8910: std_logic; attribute dont_touch of WX8910: signal is true;
	signal WX8911: std_logic; attribute dont_touch of WX8911: signal is true;
	signal WX8912: std_logic; attribute dont_touch of WX8912: signal is true;
	signal WX8913: std_logic; attribute dont_touch of WX8913: signal is true;
	signal WX8914: std_logic; attribute dont_touch of WX8914: signal is true;
	signal WX8915: std_logic; attribute dont_touch of WX8915: signal is true;
	signal WX8916: std_logic; attribute dont_touch of WX8916: signal is true;
	signal WX8917: std_logic; attribute dont_touch of WX8917: signal is true;
	signal WX8918: std_logic; attribute dont_touch of WX8918: signal is true;
	signal WX8919: std_logic; attribute dont_touch of WX8919: signal is true;
	signal WX8920: std_logic; attribute dont_touch of WX8920: signal is true;
	signal WX8921: std_logic; attribute dont_touch of WX8921: signal is true;
	signal WX8922: std_logic; attribute dont_touch of WX8922: signal is true;
	signal WX8923: std_logic; attribute dont_touch of WX8923: signal is true;
	signal WX8924: std_logic; attribute dont_touch of WX8924: signal is true;
	signal WX8925: std_logic; attribute dont_touch of WX8925: signal is true;
	signal WX8926: std_logic; attribute dont_touch of WX8926: signal is true;
	signal WX8927: std_logic; attribute dont_touch of WX8927: signal is true;
	signal WX8928: std_logic; attribute dont_touch of WX8928: signal is true;
	signal WX8929: std_logic; attribute dont_touch of WX8929: signal is true;
	signal WX8930: std_logic; attribute dont_touch of WX8930: signal is true;
	signal WX8931: std_logic; attribute dont_touch of WX8931: signal is true;
	signal WX8932: std_logic; attribute dont_touch of WX8932: signal is true;
	signal WX8933: std_logic; attribute dont_touch of WX8933: signal is true;
	signal WX8934: std_logic; attribute dont_touch of WX8934: signal is true;
	signal WX8935: std_logic; attribute dont_touch of WX8935: signal is true;
	signal WX8936: std_logic; attribute dont_touch of WX8936: signal is true;
	signal WX8937: std_logic; attribute dont_touch of WX8937: signal is true;
	signal WX8938: std_logic; attribute dont_touch of WX8938: signal is true;
	signal WX8939: std_logic; attribute dont_touch of WX8939: signal is true;
	signal WX8940: std_logic; attribute dont_touch of WX8940: signal is true;
	signal WX8941: std_logic; attribute dont_touch of WX8941: signal is true;
	signal WX8942: std_logic; attribute dont_touch of WX8942: signal is true;
	signal WX8943: std_logic; attribute dont_touch of WX8943: signal is true;
	signal WX8944: std_logic; attribute dont_touch of WX8944: signal is true;
	signal WX8945: std_logic; attribute dont_touch of WX8945: signal is true;
	signal WX8946: std_logic; attribute dont_touch of WX8946: signal is true;
	signal WX8947: std_logic; attribute dont_touch of WX8947: signal is true;
	signal WX8948: std_logic; attribute dont_touch of WX8948: signal is true;
	signal WX8949: std_logic; attribute dont_touch of WX8949: signal is true;
	signal WX8950: std_logic; attribute dont_touch of WX8950: signal is true;
	signal WX8951: std_logic; attribute dont_touch of WX8951: signal is true;
	signal WX8952: std_logic; attribute dont_touch of WX8952: signal is true;
	signal WX8953: std_logic; attribute dont_touch of WX8953: signal is true;
	signal WX8954: std_logic; attribute dont_touch of WX8954: signal is true;
	signal WX8955: std_logic; attribute dont_touch of WX8955: signal is true;
	signal WX8956: std_logic; attribute dont_touch of WX8956: signal is true;
	signal WX8957: std_logic; attribute dont_touch of WX8957: signal is true;
	signal WX8958: std_logic; attribute dont_touch of WX8958: signal is true;
	signal WX8959: std_logic; attribute dont_touch of WX8959: signal is true;
	signal WX8960: std_logic; attribute dont_touch of WX8960: signal is true;
	signal WX8961: std_logic; attribute dont_touch of WX8961: signal is true;
	signal WX8962: std_logic; attribute dont_touch of WX8962: signal is true;
	signal WX8963: std_logic; attribute dont_touch of WX8963: signal is true;
	signal WX8964: std_logic; attribute dont_touch of WX8964: signal is true;
	signal WX8965: std_logic; attribute dont_touch of WX8965: signal is true;
	signal WX8966: std_logic; attribute dont_touch of WX8966: signal is true;
	signal WX8967: std_logic; attribute dont_touch of WX8967: signal is true;
	signal WX8968: std_logic; attribute dont_touch of WX8968: signal is true;
	signal WX8969: std_logic; attribute dont_touch of WX8969: signal is true;
	signal WX8970: std_logic; attribute dont_touch of WX8970: signal is true;
	signal WX8971: std_logic; attribute dont_touch of WX8971: signal is true;
	signal WX8972: std_logic; attribute dont_touch of WX8972: signal is true;
	signal WX8973: std_logic; attribute dont_touch of WX8973: signal is true;
	signal WX8974: std_logic; attribute dont_touch of WX8974: signal is true;
	signal WX8975: std_logic; attribute dont_touch of WX8975: signal is true;
	signal WX8976: std_logic; attribute dont_touch of WX8976: signal is true;
	signal WX8977: std_logic; attribute dont_touch of WX8977: signal is true;
	signal WX8978: std_logic; attribute dont_touch of WX8978: signal is true;
	signal WX8979: std_logic; attribute dont_touch of WX8979: signal is true;
	signal WX8980: std_logic; attribute dont_touch of WX8980: signal is true;
	signal WX8981: std_logic; attribute dont_touch of WX8981: signal is true;
	signal WX8982: std_logic; attribute dont_touch of WX8982: signal is true;
	signal WX8983: std_logic; attribute dont_touch of WX8983: signal is true;
	signal WX8984: std_logic; attribute dont_touch of WX8984: signal is true;
	signal WX8985: std_logic; attribute dont_touch of WX8985: signal is true;
	signal WX8986: std_logic; attribute dont_touch of WX8986: signal is true;
	signal WX8987: std_logic; attribute dont_touch of WX8987: signal is true;
	signal WX8988: std_logic; attribute dont_touch of WX8988: signal is true;
	signal WX8989: std_logic; attribute dont_touch of WX8989: signal is true;
	signal WX8990: std_logic; attribute dont_touch of WX8990: signal is true;
	signal WX8991: std_logic; attribute dont_touch of WX8991: signal is true;
	signal WX8992: std_logic; attribute dont_touch of WX8992: signal is true;
	signal WX8993: std_logic; attribute dont_touch of WX8993: signal is true;
	signal WX8994: std_logic; attribute dont_touch of WX8994: signal is true;
	signal WX8995: std_logic; attribute dont_touch of WX8995: signal is true;
	signal WX8996: std_logic; attribute dont_touch of WX8996: signal is true;
	signal WX8997: std_logic; attribute dont_touch of WX8997: signal is true;
	signal WX8998: std_logic; attribute dont_touch of WX8998: signal is true;
	signal WX8999: std_logic; attribute dont_touch of WX8999: signal is true;
	signal WX9000: std_logic; attribute dont_touch of WX9000: signal is true;
	signal WX9001: std_logic; attribute dont_touch of WX9001: signal is true;
	signal WX9002: std_logic; attribute dont_touch of WX9002: signal is true;
	signal WX9003: std_logic; attribute dont_touch of WX9003: signal is true;
	signal WX9004: std_logic; attribute dont_touch of WX9004: signal is true;
	signal WX9005: std_logic; attribute dont_touch of WX9005: signal is true;
	signal WX9006: std_logic; attribute dont_touch of WX9006: signal is true;
	signal WX9007: std_logic; attribute dont_touch of WX9007: signal is true;
	signal WX9008: std_logic; attribute dont_touch of WX9008: signal is true;
	signal WX9009: std_logic; attribute dont_touch of WX9009: signal is true;
	signal WX9010: std_logic; attribute dont_touch of WX9010: signal is true;
	signal WX9011: std_logic; attribute dont_touch of WX9011: signal is true;
	signal WX9012: std_logic; attribute dont_touch of WX9012: signal is true;
	signal WX9013: std_logic; attribute dont_touch of WX9013: signal is true;
	signal WX9014: std_logic; attribute dont_touch of WX9014: signal is true;
	signal WX9015: std_logic; attribute dont_touch of WX9015: signal is true;
	signal WX9016: std_logic; attribute dont_touch of WX9016: signal is true;
	signal WX9017: std_logic; attribute dont_touch of WX9017: signal is true;
	signal WX9018: std_logic; attribute dont_touch of WX9018: signal is true;
	signal WX9019: std_logic; attribute dont_touch of WX9019: signal is true;
	signal WX9020: std_logic; attribute dont_touch of WX9020: signal is true;
	signal WX9021: std_logic; attribute dont_touch of WX9021: signal is true;
	signal WX9022: std_logic; attribute dont_touch of WX9022: signal is true;
	signal WX9024: std_logic; attribute dont_touch of WX9024: signal is true;
	signal WX9026: std_logic; attribute dont_touch of WX9026: signal is true;
	signal WX9028: std_logic; attribute dont_touch of WX9028: signal is true;
	signal WX9030: std_logic; attribute dont_touch of WX9030: signal is true;
	signal WX9032: std_logic; attribute dont_touch of WX9032: signal is true;
	signal WX9034: std_logic; attribute dont_touch of WX9034: signal is true;
	signal WX9036: std_logic; attribute dont_touch of WX9036: signal is true;
	signal WX9038: std_logic; attribute dont_touch of WX9038: signal is true;
	signal WX9040: std_logic; attribute dont_touch of WX9040: signal is true;
	signal WX9042: std_logic; attribute dont_touch of WX9042: signal is true;
	signal WX9044: std_logic; attribute dont_touch of WX9044: signal is true;
	signal WX9046: std_logic; attribute dont_touch of WX9046: signal is true;
	signal WX9048: std_logic; attribute dont_touch of WX9048: signal is true;
	signal WX9050: std_logic; attribute dont_touch of WX9050: signal is true;
	signal WX9052: std_logic; attribute dont_touch of WX9052: signal is true;
	signal WX9054: std_logic; attribute dont_touch of WX9054: signal is true;
	signal WX9056: std_logic; attribute dont_touch of WX9056: signal is true;
	signal WX9058: std_logic; attribute dont_touch of WX9058: signal is true;
	signal WX9060: std_logic; attribute dont_touch of WX9060: signal is true;
	signal WX9062: std_logic; attribute dont_touch of WX9062: signal is true;
	signal WX9064: std_logic; attribute dont_touch of WX9064: signal is true;
	signal WX9066: std_logic; attribute dont_touch of WX9066: signal is true;
	signal WX9068: std_logic; attribute dont_touch of WX9068: signal is true;
	signal WX9070: std_logic; attribute dont_touch of WX9070: signal is true;
	signal WX9072: std_logic; attribute dont_touch of WX9072: signal is true;
	signal WX9074: std_logic; attribute dont_touch of WX9074: signal is true;
	signal WX9076: std_logic; attribute dont_touch of WX9076: signal is true;
	signal WX9078: std_logic; attribute dont_touch of WX9078: signal is true;
	signal WX9080: std_logic; attribute dont_touch of WX9080: signal is true;
	signal WX9082: std_logic; attribute dont_touch of WX9082: signal is true;
	signal WX9084: std_logic; attribute dont_touch of WX9084: signal is true;
	signal WX9086: std_logic; attribute dont_touch of WX9086: signal is true;
	signal WX9087: std_logic; attribute dont_touch of WX9087: signal is true;
	signal WX9088: std_logic; attribute dont_touch of WX9088: signal is true;
	signal WX9089: std_logic; attribute dont_touch of WX9089: signal is true;
	signal WX9090: std_logic; attribute dont_touch of WX9090: signal is true;
	signal WX9091: std_logic; attribute dont_touch of WX9091: signal is true;
	signal WX9092: std_logic; attribute dont_touch of WX9092: signal is true;
	signal WX9093: std_logic; attribute dont_touch of WX9093: signal is true;
	signal WX9094: std_logic; attribute dont_touch of WX9094: signal is true;
	signal WX9095: std_logic; attribute dont_touch of WX9095: signal is true;
	signal WX9096: std_logic; attribute dont_touch of WX9096: signal is true;
	signal WX9097: std_logic; attribute dont_touch of WX9097: signal is true;
	signal WX9098: std_logic; attribute dont_touch of WX9098: signal is true;
	signal WX9099: std_logic; attribute dont_touch of WX9099: signal is true;
	signal WX9100: std_logic; attribute dont_touch of WX9100: signal is true;
	signal WX9101: std_logic; attribute dont_touch of WX9101: signal is true;
	signal WX9102: std_logic; attribute dont_touch of WX9102: signal is true;
	signal WX9103: std_logic; attribute dont_touch of WX9103: signal is true;
	signal WX9104: std_logic; attribute dont_touch of WX9104: signal is true;
	signal WX9105: std_logic; attribute dont_touch of WX9105: signal is true;
	signal WX9106: std_logic; attribute dont_touch of WX9106: signal is true;
	signal WX9107: std_logic; attribute dont_touch of WX9107: signal is true;
	signal WX9108: std_logic; attribute dont_touch of WX9108: signal is true;
	signal WX9109: std_logic; attribute dont_touch of WX9109: signal is true;
	signal WX9110: std_logic; attribute dont_touch of WX9110: signal is true;
	signal WX9111: std_logic; attribute dont_touch of WX9111: signal is true;
	signal WX9112: std_logic; attribute dont_touch of WX9112: signal is true;
	signal WX9113: std_logic; attribute dont_touch of WX9113: signal is true;
	signal WX9114: std_logic; attribute dont_touch of WX9114: signal is true;
	signal WX9115: std_logic; attribute dont_touch of WX9115: signal is true;
	signal WX9116: std_logic; attribute dont_touch of WX9116: signal is true;
	signal WX9117: std_logic; attribute dont_touch of WX9117: signal is true;
	signal WX9118: std_logic; attribute dont_touch of WX9118: signal is true;
	signal WX9119: std_logic; attribute dont_touch of WX9119: signal is true;
	signal WX9120: std_logic; attribute dont_touch of WX9120: signal is true;
	signal WX9121: std_logic; attribute dont_touch of WX9121: signal is true;
	signal WX9122: std_logic; attribute dont_touch of WX9122: signal is true;
	signal WX9123: std_logic; attribute dont_touch of WX9123: signal is true;
	signal WX9124: std_logic; attribute dont_touch of WX9124: signal is true;
	signal WX9125: std_logic; attribute dont_touch of WX9125: signal is true;
	signal WX9126: std_logic; attribute dont_touch of WX9126: signal is true;
	signal WX9127: std_logic; attribute dont_touch of WX9127: signal is true;
	signal WX9128: std_logic; attribute dont_touch of WX9128: signal is true;
	signal WX9129: std_logic; attribute dont_touch of WX9129: signal is true;
	signal WX9130: std_logic; attribute dont_touch of WX9130: signal is true;
	signal WX9131: std_logic; attribute dont_touch of WX9131: signal is true;
	signal WX9132: std_logic; attribute dont_touch of WX9132: signal is true;
	signal WX9133: std_logic; attribute dont_touch of WX9133: signal is true;
	signal WX9134: std_logic; attribute dont_touch of WX9134: signal is true;
	signal WX9135: std_logic; attribute dont_touch of WX9135: signal is true;
	signal WX9136: std_logic; attribute dont_touch of WX9136: signal is true;
	signal WX9137: std_logic; attribute dont_touch of WX9137: signal is true;
	signal WX9138: std_logic; attribute dont_touch of WX9138: signal is true;
	signal WX9139: std_logic; attribute dont_touch of WX9139: signal is true;
	signal WX9140: std_logic; attribute dont_touch of WX9140: signal is true;
	signal WX9141: std_logic; attribute dont_touch of WX9141: signal is true;
	signal WX9142: std_logic; attribute dont_touch of WX9142: signal is true;
	signal WX9143: std_logic; attribute dont_touch of WX9143: signal is true;
	signal WX9144: std_logic; attribute dont_touch of WX9144: signal is true;
	signal WX9145: std_logic; attribute dont_touch of WX9145: signal is true;
	signal WX9146: std_logic; attribute dont_touch of WX9146: signal is true;
	signal WX9147: std_logic; attribute dont_touch of WX9147: signal is true;
	signal WX9148: std_logic; attribute dont_touch of WX9148: signal is true;
	signal WX9149: std_logic; attribute dont_touch of WX9149: signal is true;
	signal WX9150: std_logic; attribute dont_touch of WX9150: signal is true;
	signal WX9151: std_logic; attribute dont_touch of WX9151: signal is true;
	signal WX9152: std_logic; attribute dont_touch of WX9152: signal is true;
	signal WX9153: std_logic; attribute dont_touch of WX9153: signal is true;
	signal WX9154: std_logic; attribute dont_touch of WX9154: signal is true;
	signal WX9155: std_logic; attribute dont_touch of WX9155: signal is true;
	signal WX9156: std_logic; attribute dont_touch of WX9156: signal is true;
	signal WX9157: std_logic; attribute dont_touch of WX9157: signal is true;
	signal WX9158: std_logic; attribute dont_touch of WX9158: signal is true;
	signal WX9159: std_logic; attribute dont_touch of WX9159: signal is true;
	signal WX9160: std_logic; attribute dont_touch of WX9160: signal is true;
	signal WX9161: std_logic; attribute dont_touch of WX9161: signal is true;
	signal WX9162: std_logic; attribute dont_touch of WX9162: signal is true;
	signal WX9163: std_logic; attribute dont_touch of WX9163: signal is true;
	signal WX9164: std_logic; attribute dont_touch of WX9164: signal is true;
	signal WX9165: std_logic; attribute dont_touch of WX9165: signal is true;
	signal WX9166: std_logic; attribute dont_touch of WX9166: signal is true;
	signal WX9167: std_logic; attribute dont_touch of WX9167: signal is true;
	signal WX9168: std_logic; attribute dont_touch of WX9168: signal is true;
	signal WX9169: std_logic; attribute dont_touch of WX9169: signal is true;
	signal WX9170: std_logic; attribute dont_touch of WX9170: signal is true;
	signal WX9171: std_logic; attribute dont_touch of WX9171: signal is true;
	signal WX9172: std_logic; attribute dont_touch of WX9172: signal is true;
	signal WX9173: std_logic; attribute dont_touch of WX9173: signal is true;
	signal WX9174: std_logic; attribute dont_touch of WX9174: signal is true;
	signal WX9175: std_logic; attribute dont_touch of WX9175: signal is true;
	signal WX9176: std_logic; attribute dont_touch of WX9176: signal is true;
	signal WX9177: std_logic; attribute dont_touch of WX9177: signal is true;
	signal WX9178: std_logic; attribute dont_touch of WX9178: signal is true;
	signal WX9179: std_logic; attribute dont_touch of WX9179: signal is true;
	signal WX9180: std_logic; attribute dont_touch of WX9180: signal is true;
	signal WX9181: std_logic; attribute dont_touch of WX9181: signal is true;
	signal WX9182: std_logic; attribute dont_touch of WX9182: signal is true;
	signal WX9183: std_logic; attribute dont_touch of WX9183: signal is true;
	signal WX9184: std_logic; attribute dont_touch of WX9184: signal is true;
	signal WX9185: std_logic; attribute dont_touch of WX9185: signal is true;
	signal WX9186: std_logic; attribute dont_touch of WX9186: signal is true;
	signal WX9187: std_logic; attribute dont_touch of WX9187: signal is true;
	signal WX9188: std_logic; attribute dont_touch of WX9188: signal is true;
	signal WX9189: std_logic; attribute dont_touch of WX9189: signal is true;
	signal WX9190: std_logic; attribute dont_touch of WX9190: signal is true;
	signal WX9191: std_logic; attribute dont_touch of WX9191: signal is true;
	signal WX9192: std_logic; attribute dont_touch of WX9192: signal is true;
	signal WX9193: std_logic; attribute dont_touch of WX9193: signal is true;
	signal WX9194: std_logic; attribute dont_touch of WX9194: signal is true;
	signal WX9195: std_logic; attribute dont_touch of WX9195: signal is true;
	signal WX9196: std_logic; attribute dont_touch of WX9196: signal is true;
	signal WX9197: std_logic; attribute dont_touch of WX9197: signal is true;
	signal WX9198: std_logic; attribute dont_touch of WX9198: signal is true;
	signal WX9199: std_logic; attribute dont_touch of WX9199: signal is true;
	signal WX9200: std_logic; attribute dont_touch of WX9200: signal is true;
	signal WX9201: std_logic; attribute dont_touch of WX9201: signal is true;
	signal WX9202: std_logic; attribute dont_touch of WX9202: signal is true;
	signal WX9203: std_logic; attribute dont_touch of WX9203: signal is true;
	signal WX9204: std_logic; attribute dont_touch of WX9204: signal is true;
	signal WX9205: std_logic; attribute dont_touch of WX9205: signal is true;
	signal WX9206: std_logic; attribute dont_touch of WX9206: signal is true;
	signal WX9207: std_logic; attribute dont_touch of WX9207: signal is true;
	signal WX9208: std_logic; attribute dont_touch of WX9208: signal is true;
	signal WX9209: std_logic; attribute dont_touch of WX9209: signal is true;
	signal WX9210: std_logic; attribute dont_touch of WX9210: signal is true;
	signal WX9211: std_logic; attribute dont_touch of WX9211: signal is true;
	signal WX9212: std_logic; attribute dont_touch of WX9212: signal is true;
	signal WX9213: std_logic; attribute dont_touch of WX9213: signal is true;
	signal WX9214: std_logic; attribute dont_touch of WX9214: signal is true;
	signal WX9215: std_logic; attribute dont_touch of WX9215: signal is true;
	signal WX9216: std_logic; attribute dont_touch of WX9216: signal is true;
	signal WX9217: std_logic; attribute dont_touch of WX9217: signal is true;
	signal WX9218: std_logic; attribute dont_touch of WX9218: signal is true;
	signal WX9219: std_logic; attribute dont_touch of WX9219: signal is true;
	signal WX9220: std_logic; attribute dont_touch of WX9220: signal is true;
	signal WX9221: std_logic; attribute dont_touch of WX9221: signal is true;
	signal WX9222: std_logic; attribute dont_touch of WX9222: signal is true;
	signal WX9223: std_logic; attribute dont_touch of WX9223: signal is true;
	signal WX9224: std_logic; attribute dont_touch of WX9224: signal is true;
	signal WX9225: std_logic; attribute dont_touch of WX9225: signal is true;
	signal WX9226: std_logic; attribute dont_touch of WX9226: signal is true;
	signal WX9227: std_logic; attribute dont_touch of WX9227: signal is true;
	signal WX9228: std_logic; attribute dont_touch of WX9228: signal is true;
	signal WX9229: std_logic; attribute dont_touch of WX9229: signal is true;
	signal WX9230: std_logic; attribute dont_touch of WX9230: signal is true;
	signal WX9231: std_logic; attribute dont_touch of WX9231: signal is true;
	signal WX9232: std_logic; attribute dont_touch of WX9232: signal is true;
	signal WX9233: std_logic; attribute dont_touch of WX9233: signal is true;
	signal WX9234: std_logic; attribute dont_touch of WX9234: signal is true;
	signal WX9235: std_logic; attribute dont_touch of WX9235: signal is true;
	signal WX9236: std_logic; attribute dont_touch of WX9236: signal is true;
	signal WX9237: std_logic; attribute dont_touch of WX9237: signal is true;
	signal WX9238: std_logic; attribute dont_touch of WX9238: signal is true;
	signal WX9239: std_logic; attribute dont_touch of WX9239: signal is true;
	signal WX9240: std_logic; attribute dont_touch of WX9240: signal is true;
	signal WX9241: std_logic; attribute dont_touch of WX9241: signal is true;
	signal WX9242: std_logic; attribute dont_touch of WX9242: signal is true;
	signal WX9243: std_logic; attribute dont_touch of WX9243: signal is true;
	signal WX9244: std_logic; attribute dont_touch of WX9244: signal is true;
	signal WX9245: std_logic; attribute dont_touch of WX9245: signal is true;
	signal WX9246: std_logic; attribute dont_touch of WX9246: signal is true;
	signal WX9247: std_logic; attribute dont_touch of WX9247: signal is true;
	signal WX9248: std_logic; attribute dont_touch of WX9248: signal is true;
	signal WX9249: std_logic; attribute dont_touch of WX9249: signal is true;
	signal WX9250: std_logic; attribute dont_touch of WX9250: signal is true;
	signal WX9251: std_logic; attribute dont_touch of WX9251: signal is true;
	signal WX9252: std_logic; attribute dont_touch of WX9252: signal is true;
	signal WX9253: std_logic; attribute dont_touch of WX9253: signal is true;
	signal WX9254: std_logic; attribute dont_touch of WX9254: signal is true;
	signal WX9255: std_logic; attribute dont_touch of WX9255: signal is true;
	signal WX9256: std_logic; attribute dont_touch of WX9256: signal is true;
	signal WX9257: std_logic; attribute dont_touch of WX9257: signal is true;
	signal WX9258: std_logic; attribute dont_touch of WX9258: signal is true;
	signal WX9259: std_logic; attribute dont_touch of WX9259: signal is true;
	signal WX9260: std_logic; attribute dont_touch of WX9260: signal is true;
	signal WX9261: std_logic; attribute dont_touch of WX9261: signal is true;
	signal WX9262: std_logic; attribute dont_touch of WX9262: signal is true;
	signal WX9263: std_logic; attribute dont_touch of WX9263: signal is true;
	signal WX9264: std_logic; attribute dont_touch of WX9264: signal is true;
	signal WX9265: std_logic; attribute dont_touch of WX9265: signal is true;
	signal WX9266: std_logic; attribute dont_touch of WX9266: signal is true;
	signal WX9267: std_logic; attribute dont_touch of WX9267: signal is true;
	signal WX9268: std_logic; attribute dont_touch of WX9268: signal is true;
	signal WX9269: std_logic; attribute dont_touch of WX9269: signal is true;
	signal WX9270: std_logic; attribute dont_touch of WX9270: signal is true;
	signal WX9271: std_logic; attribute dont_touch of WX9271: signal is true;
	signal WX9272: std_logic; attribute dont_touch of WX9272: signal is true;
	signal WX9273: std_logic; attribute dont_touch of WX9273: signal is true;
	signal WX9274: std_logic; attribute dont_touch of WX9274: signal is true;
	signal WX9275: std_logic; attribute dont_touch of WX9275: signal is true;
	signal WX9276: std_logic; attribute dont_touch of WX9276: signal is true;
	signal WX9277: std_logic; attribute dont_touch of WX9277: signal is true;
	signal WX9278: std_logic; attribute dont_touch of WX9278: signal is true;
	signal WX9279: std_logic; attribute dont_touch of WX9279: signal is true;
	signal WX9280: std_logic; attribute dont_touch of WX9280: signal is true;
	signal WX9281: std_logic; attribute dont_touch of WX9281: signal is true;
	signal WX9282: std_logic; attribute dont_touch of WX9282: signal is true;
	signal WX9283: std_logic; attribute dont_touch of WX9283: signal is true;
	signal WX9284: std_logic; attribute dont_touch of WX9284: signal is true;
	signal WX9285: std_logic; attribute dont_touch of WX9285: signal is true;
	signal WX9286: std_logic; attribute dont_touch of WX9286: signal is true;
	signal WX9287: std_logic; attribute dont_touch of WX9287: signal is true;
	signal WX9288: std_logic; attribute dont_touch of WX9288: signal is true;
	signal WX9289: std_logic; attribute dont_touch of WX9289: signal is true;
	signal WX9290: std_logic; attribute dont_touch of WX9290: signal is true;
	signal WX9291: std_logic; attribute dont_touch of WX9291: signal is true;
	signal WX9292: std_logic; attribute dont_touch of WX9292: signal is true;
	signal WX9293: std_logic; attribute dont_touch of WX9293: signal is true;
	signal WX9294: std_logic; attribute dont_touch of WX9294: signal is true;
	signal WX9295: std_logic; attribute dont_touch of WX9295: signal is true;
	signal WX9296: std_logic; attribute dont_touch of WX9296: signal is true;
	signal WX9297: std_logic; attribute dont_touch of WX9297: signal is true;
	signal WX9298: std_logic; attribute dont_touch of WX9298: signal is true;
	signal WX9299: std_logic; attribute dont_touch of WX9299: signal is true;
	signal WX9300: std_logic; attribute dont_touch of WX9300: signal is true;
	signal WX9301: std_logic; attribute dont_touch of WX9301: signal is true;
	signal WX9302: std_logic; attribute dont_touch of WX9302: signal is true;
	signal WX9303: std_logic; attribute dont_touch of WX9303: signal is true;
	signal WX9304: std_logic; attribute dont_touch of WX9304: signal is true;
	signal WX9305: std_logic; attribute dont_touch of WX9305: signal is true;
	signal WX9306: std_logic; attribute dont_touch of WX9306: signal is true;
	signal WX9307: std_logic; attribute dont_touch of WX9307: signal is true;
	signal WX9308: std_logic; attribute dont_touch of WX9308: signal is true;
	signal WX9309: std_logic; attribute dont_touch of WX9309: signal is true;
	signal WX9310: std_logic; attribute dont_touch of WX9310: signal is true;
	signal WX9311: std_logic; attribute dont_touch of WX9311: signal is true;
	signal WX9312: std_logic; attribute dont_touch of WX9312: signal is true;
	signal WX9313: std_logic; attribute dont_touch of WX9313: signal is true;
	signal WX9314: std_logic; attribute dont_touch of WX9314: signal is true;
	signal WX9315: std_logic; attribute dont_touch of WX9315: signal is true;
	signal WX9316: std_logic; attribute dont_touch of WX9316: signal is true;
	signal WX9317: std_logic; attribute dont_touch of WX9317: signal is true;
	signal WX9318: std_logic; attribute dont_touch of WX9318: signal is true;
	signal WX9319: std_logic; attribute dont_touch of WX9319: signal is true;
	signal WX9320: std_logic; attribute dont_touch of WX9320: signal is true;
	signal WX9321: std_logic; attribute dont_touch of WX9321: signal is true;
	signal WX9322: std_logic; attribute dont_touch of WX9322: signal is true;
	signal WX9323: std_logic; attribute dont_touch of WX9323: signal is true;
	signal WX9324: std_logic; attribute dont_touch of WX9324: signal is true;
	signal WX9325: std_logic; attribute dont_touch of WX9325: signal is true;
	signal WX9326: std_logic; attribute dont_touch of WX9326: signal is true;
	signal WX9327: std_logic; attribute dont_touch of WX9327: signal is true;
	signal WX9328: std_logic; attribute dont_touch of WX9328: signal is true;
	signal WX9329: std_logic; attribute dont_touch of WX9329: signal is true;
	signal WX9330: std_logic; attribute dont_touch of WX9330: signal is true;
	signal WX9331: std_logic; attribute dont_touch of WX9331: signal is true;
	signal WX9332: std_logic; attribute dont_touch of WX9332: signal is true;
	signal WX9333: std_logic; attribute dont_touch of WX9333: signal is true;
	signal WX9334: std_logic; attribute dont_touch of WX9334: signal is true;
	signal WX9335: std_logic; attribute dont_touch of WX9335: signal is true;
	signal WX9336: std_logic; attribute dont_touch of WX9336: signal is true;
	signal WX9337: std_logic; attribute dont_touch of WX9337: signal is true;
	signal WX9338: std_logic; attribute dont_touch of WX9338: signal is true;
	signal WX9339: std_logic; attribute dont_touch of WX9339: signal is true;
	signal WX9340: std_logic; attribute dont_touch of WX9340: signal is true;
	signal WX9341: std_logic; attribute dont_touch of WX9341: signal is true;
	signal WX9342: std_logic; attribute dont_touch of WX9342: signal is true;
	signal WX9343: std_logic; attribute dont_touch of WX9343: signal is true;
	signal WX9344: std_logic; attribute dont_touch of WX9344: signal is true;
	signal WX9345: std_logic; attribute dont_touch of WX9345: signal is true;
	signal WX9346: std_logic; attribute dont_touch of WX9346: signal is true;
	signal WX9347: std_logic; attribute dont_touch of WX9347: signal is true;
	signal WX9348: std_logic; attribute dont_touch of WX9348: signal is true;
	signal WX9349: std_logic; attribute dont_touch of WX9349: signal is true;
	signal WX9350: std_logic; attribute dont_touch of WX9350: signal is true;
	signal WX9351: std_logic; attribute dont_touch of WX9351: signal is true;
	signal WX9352: std_logic; attribute dont_touch of WX9352: signal is true;
	signal WX9353: std_logic; attribute dont_touch of WX9353: signal is true;
	signal WX9354: std_logic; attribute dont_touch of WX9354: signal is true;
	signal WX9355: std_logic; attribute dont_touch of WX9355: signal is true;
	signal WX9356: std_logic; attribute dont_touch of WX9356: signal is true;
	signal WX9357: std_logic; attribute dont_touch of WX9357: signal is true;
	signal WX9358: std_logic; attribute dont_touch of WX9358: signal is true;
	signal WX9359: std_logic; attribute dont_touch of WX9359: signal is true;
	signal WX9360: std_logic; attribute dont_touch of WX9360: signal is true;
	signal WX9361: std_logic; attribute dont_touch of WX9361: signal is true;
	signal WX9362: std_logic; attribute dont_touch of WX9362: signal is true;
	signal WX9363: std_logic; attribute dont_touch of WX9363: signal is true;
	signal WX9364: std_logic; attribute dont_touch of WX9364: signal is true;
	signal WX9365: std_logic; attribute dont_touch of WX9365: signal is true;
	signal WX9366: std_logic; attribute dont_touch of WX9366: signal is true;
	signal WX9367: std_logic; attribute dont_touch of WX9367: signal is true;
	signal WX9368: std_logic; attribute dont_touch of WX9368: signal is true;
	signal WX9369: std_logic; attribute dont_touch of WX9369: signal is true;
	signal WX9370: std_logic; attribute dont_touch of WX9370: signal is true;
	signal WX9371: std_logic; attribute dont_touch of WX9371: signal is true;
	signal WX9372: std_logic; attribute dont_touch of WX9372: signal is true;
	signal WX9373: std_logic; attribute dont_touch of WX9373: signal is true;
	signal WX9374: std_logic; attribute dont_touch of WX9374: signal is true;
	signal WX9375: std_logic; attribute dont_touch of WX9375: signal is true;
	signal WX9376: std_logic; attribute dont_touch of WX9376: signal is true;
	signal WX9377: std_logic; attribute dont_touch of WX9377: signal is true;
	signal WX9378: std_logic; attribute dont_touch of WX9378: signal is true;
	signal WX9379: std_logic; attribute dont_touch of WX9379: signal is true;
	signal WX9380: std_logic; attribute dont_touch of WX9380: signal is true;
	signal WX9381: std_logic; attribute dont_touch of WX9381: signal is true;
	signal WX9382: std_logic; attribute dont_touch of WX9382: signal is true;
	signal WX9383: std_logic; attribute dont_touch of WX9383: signal is true;
	signal WX9384: std_logic; attribute dont_touch of WX9384: signal is true;
	signal WX9385: std_logic; attribute dont_touch of WX9385: signal is true;
	signal WX9386: std_logic; attribute dont_touch of WX9386: signal is true;
	signal WX9387: std_logic; attribute dont_touch of WX9387: signal is true;
	signal WX9388: std_logic; attribute dont_touch of WX9388: signal is true;
	signal WX9389: std_logic; attribute dont_touch of WX9389: signal is true;
	signal WX9390: std_logic; attribute dont_touch of WX9390: signal is true;
	signal WX9391: std_logic; attribute dont_touch of WX9391: signal is true;
	signal WX9392: std_logic; attribute dont_touch of WX9392: signal is true;
	signal WX9393: std_logic; attribute dont_touch of WX9393: signal is true;
	signal WX9394: std_logic; attribute dont_touch of WX9394: signal is true;
	signal WX9395: std_logic; attribute dont_touch of WX9395: signal is true;
	signal WX9396: std_logic; attribute dont_touch of WX9396: signal is true;
	signal WX9397: std_logic; attribute dont_touch of WX9397: signal is true;
	signal WX9398: std_logic; attribute dont_touch of WX9398: signal is true;
	signal WX9399: std_logic; attribute dont_touch of WX9399: signal is true;
	signal WX9400: std_logic; attribute dont_touch of WX9400: signal is true;
	signal WX9401: std_logic; attribute dont_touch of WX9401: signal is true;
	signal WX9402: std_logic; attribute dont_touch of WX9402: signal is true;
	signal WX9403: std_logic; attribute dont_touch of WX9403: signal is true;
	signal WX9404: std_logic; attribute dont_touch of WX9404: signal is true;
	signal WX9405: std_logic; attribute dont_touch of WX9405: signal is true;
	signal WX9406: std_logic; attribute dont_touch of WX9406: signal is true;
	signal WX9407: std_logic; attribute dont_touch of WX9407: signal is true;
	signal WX9408: std_logic; attribute dont_touch of WX9408: signal is true;
	signal WX9409: std_logic; attribute dont_touch of WX9409: signal is true;
	signal WX9410: std_logic; attribute dont_touch of WX9410: signal is true;
	signal WX9411: std_logic; attribute dont_touch of WX9411: signal is true;
	signal WX9412: std_logic; attribute dont_touch of WX9412: signal is true;
	signal WX9413: std_logic; attribute dont_touch of WX9413: signal is true;
	signal WX9414: std_logic; attribute dont_touch of WX9414: signal is true;
	signal WX9415: std_logic; attribute dont_touch of WX9415: signal is true;
	signal WX9416: std_logic; attribute dont_touch of WX9416: signal is true;
	signal WX9417: std_logic; attribute dont_touch of WX9417: signal is true;
	signal WX9418: std_logic; attribute dont_touch of WX9418: signal is true;
	signal WX9419: std_logic; attribute dont_touch of WX9419: signal is true;
	signal WX9420: std_logic; attribute dont_touch of WX9420: signal is true;
	signal WX9421: std_logic; attribute dont_touch of WX9421: signal is true;
	signal WX9422: std_logic; attribute dont_touch of WX9422: signal is true;
	signal WX9423: std_logic; attribute dont_touch of WX9423: signal is true;
	signal WX9424: std_logic; attribute dont_touch of WX9424: signal is true;
	signal WX9425: std_logic; attribute dont_touch of WX9425: signal is true;
	signal WX9426: std_logic; attribute dont_touch of WX9426: signal is true;
	signal WX9427: std_logic; attribute dont_touch of WX9427: signal is true;
	signal WX9428: std_logic; attribute dont_touch of WX9428: signal is true;
	signal WX9429: std_logic; attribute dont_touch of WX9429: signal is true;
	signal WX9430: std_logic; attribute dont_touch of WX9430: signal is true;
	signal WX9431: std_logic; attribute dont_touch of WX9431: signal is true;
	signal WX9432: std_logic; attribute dont_touch of WX9432: signal is true;
	signal WX9433: std_logic; attribute dont_touch of WX9433: signal is true;
	signal WX9434: std_logic; attribute dont_touch of WX9434: signal is true;
	signal WX9435: std_logic; attribute dont_touch of WX9435: signal is true;
	signal WX9436: std_logic; attribute dont_touch of WX9436: signal is true;
	signal WX9437: std_logic; attribute dont_touch of WX9437: signal is true;
	signal WX9438: std_logic; attribute dont_touch of WX9438: signal is true;
	signal WX9439: std_logic; attribute dont_touch of WX9439: signal is true;
	signal WX9440: std_logic; attribute dont_touch of WX9440: signal is true;
	signal WX9441: std_logic; attribute dont_touch of WX9441: signal is true;
	signal WX9442: std_logic; attribute dont_touch of WX9442: signal is true;
	signal WX9443: std_logic; attribute dont_touch of WX9443: signal is true;
	signal WX9444: std_logic; attribute dont_touch of WX9444: signal is true;
	signal WX9445: std_logic; attribute dont_touch of WX9445: signal is true;
	signal WX9446: std_logic; attribute dont_touch of WX9446: signal is true;
	signal WX9447: std_logic; attribute dont_touch of WX9447: signal is true;
	signal WX9448: std_logic; attribute dont_touch of WX9448: signal is true;
	signal WX9449: std_logic; attribute dont_touch of WX9449: signal is true;
	signal WX9450: std_logic; attribute dont_touch of WX9450: signal is true;
	signal WX9451: std_logic; attribute dont_touch of WX9451: signal is true;
	signal WX9452: std_logic; attribute dont_touch of WX9452: signal is true;
	signal WX9453: std_logic; attribute dont_touch of WX9453: signal is true;
	signal WX9454: std_logic; attribute dont_touch of WX9454: signal is true;
	signal WX9455: std_logic; attribute dont_touch of WX9455: signal is true;
	signal WX9456: std_logic; attribute dont_touch of WX9456: signal is true;
	signal WX9457: std_logic; attribute dont_touch of WX9457: signal is true;
	signal WX9458: std_logic; attribute dont_touch of WX9458: signal is true;
	signal WX9459: std_logic; attribute dont_touch of WX9459: signal is true;
	signal WX9460: std_logic; attribute dont_touch of WX9460: signal is true;
	signal WX9461: std_logic; attribute dont_touch of WX9461: signal is true;
	signal WX9462: std_logic; attribute dont_touch of WX9462: signal is true;
	signal WX9463: std_logic; attribute dont_touch of WX9463: signal is true;
	signal WX9464: std_logic; attribute dont_touch of WX9464: signal is true;
	signal WX9465: std_logic; attribute dont_touch of WX9465: signal is true;
	signal WX9466: std_logic; attribute dont_touch of WX9466: signal is true;
	signal WX9467: std_logic; attribute dont_touch of WX9467: signal is true;
	signal WX9468: std_logic; attribute dont_touch of WX9468: signal is true;
	signal WX9469: std_logic; attribute dont_touch of WX9469: signal is true;
	signal WX9470: std_logic; attribute dont_touch of WX9470: signal is true;
	signal WX9471: std_logic; attribute dont_touch of WX9471: signal is true;
	signal WX9472: std_logic; attribute dont_touch of WX9472: signal is true;
	signal WX9473: std_logic; attribute dont_touch of WX9473: signal is true;
	signal WX9474: std_logic; attribute dont_touch of WX9474: signal is true;
	signal WX9475: std_logic; attribute dont_touch of WX9475: signal is true;
	signal WX9476: std_logic; attribute dont_touch of WX9476: signal is true;
	signal WX9477: std_logic; attribute dont_touch of WX9477: signal is true;
	signal WX9478: std_logic; attribute dont_touch of WX9478: signal is true;
	signal WX9479: std_logic; attribute dont_touch of WX9479: signal is true;
	signal WX9480: std_logic; attribute dont_touch of WX9480: signal is true;
	signal WX9481: std_logic; attribute dont_touch of WX9481: signal is true;
	signal WX9482: std_logic; attribute dont_touch of WX9482: signal is true;
	signal WX9483: std_logic; attribute dont_touch of WX9483: signal is true;
	signal WX9484: std_logic; attribute dont_touch of WX9484: signal is true;
	signal WX9485: std_logic; attribute dont_touch of WX9485: signal is true;
	signal WX9486: std_logic; attribute dont_touch of WX9486: signal is true;
	signal WX9487: std_logic; attribute dont_touch of WX9487: signal is true;
	signal WX9488: std_logic; attribute dont_touch of WX9488: signal is true;
	signal WX9489: std_logic; attribute dont_touch of WX9489: signal is true;
	signal WX9490: std_logic; attribute dont_touch of WX9490: signal is true;
	signal WX9491: std_logic; attribute dont_touch of WX9491: signal is true;
	signal WX9492: std_logic; attribute dont_touch of WX9492: signal is true;
	signal WX9493: std_logic; attribute dont_touch of WX9493: signal is true;
	signal WX9494: std_logic; attribute dont_touch of WX9494: signal is true;
	signal WX9495: std_logic; attribute dont_touch of WX9495: signal is true;
	signal WX9496: std_logic; attribute dont_touch of WX9496: signal is true;
	signal WX9497: std_logic; attribute dont_touch of WX9497: signal is true;
	signal WX9498: std_logic; attribute dont_touch of WX9498: signal is true;
	signal WX9499: std_logic; attribute dont_touch of WX9499: signal is true;
	signal WX9500: std_logic; attribute dont_touch of WX9500: signal is true;
	signal WX9501: std_logic; attribute dont_touch of WX9501: signal is true;
	signal WX9502: std_logic; attribute dont_touch of WX9502: signal is true;
	signal WX9503: std_logic; attribute dont_touch of WX9503: signal is true;
	signal WX9504: std_logic; attribute dont_touch of WX9504: signal is true;
	signal WX9505: std_logic; attribute dont_touch of WX9505: signal is true;
	signal WX9506: std_logic; attribute dont_touch of WX9506: signal is true;
	signal WX9507: std_logic; attribute dont_touch of WX9507: signal is true;
	signal WX9508: std_logic; attribute dont_touch of WX9508: signal is true;
	signal WX9509: std_logic; attribute dont_touch of WX9509: signal is true;
	signal WX9510: std_logic; attribute dont_touch of WX9510: signal is true;
	signal WX9511: std_logic; attribute dont_touch of WX9511: signal is true;
	signal WX9512: std_logic; attribute dont_touch of WX9512: signal is true;
	signal WX9513: std_logic; attribute dont_touch of WX9513: signal is true;
	signal WX9514: std_logic; attribute dont_touch of WX9514: signal is true;
	signal WX9515: std_logic; attribute dont_touch of WX9515: signal is true;
	signal WX9516: std_logic; attribute dont_touch of WX9516: signal is true;
	signal WX9517: std_logic; attribute dont_touch of WX9517: signal is true;
	signal WX9518: std_logic; attribute dont_touch of WX9518: signal is true;
	signal WX9519: std_logic; attribute dont_touch of WX9519: signal is true;
	signal WX9520: std_logic; attribute dont_touch of WX9520: signal is true;
	signal WX9521: std_logic; attribute dont_touch of WX9521: signal is true;
	signal WX9522: std_logic; attribute dont_touch of WX9522: signal is true;
	signal WX9523: std_logic; attribute dont_touch of WX9523: signal is true;
	signal WX9524: std_logic; attribute dont_touch of WX9524: signal is true;
	signal WX9525: std_logic; attribute dont_touch of WX9525: signal is true;
	signal WX9526: std_logic; attribute dont_touch of WX9526: signal is true;
	signal WX9527: std_logic; attribute dont_touch of WX9527: signal is true;
	signal WX9528: std_logic; attribute dont_touch of WX9528: signal is true;
	signal WX9529: std_logic; attribute dont_touch of WX9529: signal is true;
	signal WX9530: std_logic; attribute dont_touch of WX9530: signal is true;
	signal WX9531: std_logic; attribute dont_touch of WX9531: signal is true;
	signal WX9532: std_logic; attribute dont_touch of WX9532: signal is true;
	signal WX9533: std_logic; attribute dont_touch of WX9533: signal is true;
	signal WX9534: std_logic; attribute dont_touch of WX9534: signal is true;
	signal WX9535: std_logic; attribute dont_touch of WX9535: signal is true;
	signal WX9536: std_logic; attribute dont_touch of WX9536: signal is true;
	signal WX9537: std_logic; attribute dont_touch of WX9537: signal is true;
	signal WX9538: std_logic; attribute dont_touch of WX9538: signal is true;
	signal WX9539: std_logic; attribute dont_touch of WX9539: signal is true;
	signal WX9540: std_logic; attribute dont_touch of WX9540: signal is true;
	signal WX9541: std_logic; attribute dont_touch of WX9541: signal is true;
	signal WX9542: std_logic; attribute dont_touch of WX9542: signal is true;
	signal WX9543: std_logic; attribute dont_touch of WX9543: signal is true;
	signal WX9544: std_logic; attribute dont_touch of WX9544: signal is true;
	signal WX9545: std_logic; attribute dont_touch of WX9545: signal is true;
	signal WX9546: std_logic; attribute dont_touch of WX9546: signal is true;
	signal WX9547: std_logic; attribute dont_touch of WX9547: signal is true;
	signal WX9548: std_logic; attribute dont_touch of WX9548: signal is true;
	signal WX9549: std_logic; attribute dont_touch of WX9549: signal is true;
	signal WX9550: std_logic; attribute dont_touch of WX9550: signal is true;
	signal WX9551: std_logic; attribute dont_touch of WX9551: signal is true;
	signal WX9552: std_logic; attribute dont_touch of WX9552: signal is true;
	signal WX9553: std_logic; attribute dont_touch of WX9553: signal is true;
	signal WX9554: std_logic; attribute dont_touch of WX9554: signal is true;
	signal WX9555: std_logic; attribute dont_touch of WX9555: signal is true;
	signal WX9556: std_logic; attribute dont_touch of WX9556: signal is true;
	signal WX9557: std_logic; attribute dont_touch of WX9557: signal is true;
	signal WX9558: std_logic; attribute dont_touch of WX9558: signal is true;
	signal WX9559: std_logic; attribute dont_touch of WX9559: signal is true;
	signal WX9560: std_logic; attribute dont_touch of WX9560: signal is true;
	signal WX9561: std_logic; attribute dont_touch of WX9561: signal is true;
	signal WX9562: std_logic; attribute dont_touch of WX9562: signal is true;
	signal WX9563: std_logic; attribute dont_touch of WX9563: signal is true;
	signal WX9564: std_logic; attribute dont_touch of WX9564: signal is true;
	signal WX9565: std_logic; attribute dont_touch of WX9565: signal is true;
	signal WX9566: std_logic; attribute dont_touch of WX9566: signal is true;
	signal WX9567: std_logic; attribute dont_touch of WX9567: signal is true;
	signal WX9568: std_logic; attribute dont_touch of WX9568: signal is true;
	signal WX9569: std_logic; attribute dont_touch of WX9569: signal is true;
	signal WX9570: std_logic; attribute dont_touch of WX9570: signal is true;
	signal WX9571: std_logic; attribute dont_touch of WX9571: signal is true;
	signal WX9572: std_logic; attribute dont_touch of WX9572: signal is true;
	signal WX9573: std_logic; attribute dont_touch of WX9573: signal is true;
	signal WX9574: std_logic; attribute dont_touch of WX9574: signal is true;
	signal WX9575: std_logic; attribute dont_touch of WX9575: signal is true;
	signal WX9576: std_logic; attribute dont_touch of WX9576: signal is true;
	signal WX9577: std_logic; attribute dont_touch of WX9577: signal is true;
	signal WX9578: std_logic; attribute dont_touch of WX9578: signal is true;
	signal WX9579: std_logic; attribute dont_touch of WX9579: signal is true;
	signal WX9580: std_logic; attribute dont_touch of WX9580: signal is true;
	signal WX9581: std_logic; attribute dont_touch of WX9581: signal is true;
	signal WX9582: std_logic; attribute dont_touch of WX9582: signal is true;
	signal WX9583: std_logic; attribute dont_touch of WX9583: signal is true;
	signal WX9584: std_logic; attribute dont_touch of WX9584: signal is true;
	signal WX9585: std_logic; attribute dont_touch of WX9585: signal is true;
	signal WX9586: std_logic; attribute dont_touch of WX9586: signal is true;
	signal WX9587: std_logic; attribute dont_touch of WX9587: signal is true;
	signal WX9588: std_logic; attribute dont_touch of WX9588: signal is true;
	signal WX9589: std_logic; attribute dont_touch of WX9589: signal is true;
	signal WX9590: std_logic; attribute dont_touch of WX9590: signal is true;
	signal WX9591: std_logic; attribute dont_touch of WX9591: signal is true;
	signal WX9592: std_logic; attribute dont_touch of WX9592: signal is true;
	signal WX9593: std_logic; attribute dont_touch of WX9593: signal is true;
	signal WX9594: std_logic; attribute dont_touch of WX9594: signal is true;
	signal WX9595: std_logic; attribute dont_touch of WX9595: signal is true;
	signal WX9596: std_logic; attribute dont_touch of WX9596: signal is true;
	signal WX9597: std_logic; attribute dont_touch of WX9597: signal is true;
	signal WX9598: std_logic; attribute dont_touch of WX9598: signal is true;
	signal WX9599: std_logic; attribute dont_touch of WX9599: signal is true;
	signal WX9600: std_logic; attribute dont_touch of WX9600: signal is true;
	signal WX9601: std_logic; attribute dont_touch of WX9601: signal is true;
	signal WX9602: std_logic; attribute dont_touch of WX9602: signal is true;
	signal WX9603: std_logic; attribute dont_touch of WX9603: signal is true;
	signal WX9604: std_logic; attribute dont_touch of WX9604: signal is true;
	signal WX9605: std_logic; attribute dont_touch of WX9605: signal is true;
	signal WX9606: std_logic; attribute dont_touch of WX9606: signal is true;
	signal WX9607: std_logic; attribute dont_touch of WX9607: signal is true;
	signal WX9608: std_logic; attribute dont_touch of WX9608: signal is true;
	signal WX9609: std_logic; attribute dont_touch of WX9609: signal is true;
	signal WX9610: std_logic; attribute dont_touch of WX9610: signal is true;
	signal WX9611: std_logic; attribute dont_touch of WX9611: signal is true;
	signal WX9612: std_logic; attribute dont_touch of WX9612: signal is true;
	signal WX9613: std_logic; attribute dont_touch of WX9613: signal is true;
	signal WX9614: std_logic; attribute dont_touch of WX9614: signal is true;
	signal WX9615: std_logic; attribute dont_touch of WX9615: signal is true;
	signal WX9616: std_logic; attribute dont_touch of WX9616: signal is true;
	signal WX9617: std_logic; attribute dont_touch of WX9617: signal is true;
	signal WX9618: std_logic; attribute dont_touch of WX9618: signal is true;
	signal WX9619: std_logic; attribute dont_touch of WX9619: signal is true;
	signal WX9620: std_logic; attribute dont_touch of WX9620: signal is true;
	signal WX9621: std_logic; attribute dont_touch of WX9621: signal is true;
	signal WX9622: std_logic; attribute dont_touch of WX9622: signal is true;
	signal WX9623: std_logic; attribute dont_touch of WX9623: signal is true;
	signal WX9624: std_logic; attribute dont_touch of WX9624: signal is true;
	signal WX9625: std_logic; attribute dont_touch of WX9625: signal is true;
	signal WX9626: std_logic; attribute dont_touch of WX9626: signal is true;
	signal WX9627: std_logic; attribute dont_touch of WX9627: signal is true;
	signal WX9628: std_logic; attribute dont_touch of WX9628: signal is true;
	signal WX9629: std_logic; attribute dont_touch of WX9629: signal is true;
	signal WX9630: std_logic; attribute dont_touch of WX9630: signal is true;
	signal WX9631: std_logic; attribute dont_touch of WX9631: signal is true;
	signal WX9632: std_logic; attribute dont_touch of WX9632: signal is true;
	signal WX9633: std_logic; attribute dont_touch of WX9633: signal is true;
	signal WX9634: std_logic; attribute dont_touch of WX9634: signal is true;
	signal WX9635: std_logic; attribute dont_touch of WX9635: signal is true;
	signal WX9636: std_logic; attribute dont_touch of WX9636: signal is true;
	signal WX9637: std_logic; attribute dont_touch of WX9637: signal is true;
	signal WX9638: std_logic; attribute dont_touch of WX9638: signal is true;
	signal WX9639: std_logic; attribute dont_touch of WX9639: signal is true;
	signal WX9640: std_logic; attribute dont_touch of WX9640: signal is true;
	signal WX9641: std_logic; attribute dont_touch of WX9641: signal is true;
	signal WX9642: std_logic; attribute dont_touch of WX9642: signal is true;
	signal WX9643: std_logic; attribute dont_touch of WX9643: signal is true;
	signal WX9644: std_logic; attribute dont_touch of WX9644: signal is true;
	signal WX9645: std_logic; attribute dont_touch of WX9645: signal is true;
	signal WX9646: std_logic; attribute dont_touch of WX9646: signal is true;
	signal WX9647: std_logic; attribute dont_touch of WX9647: signal is true;
	signal WX9648: std_logic; attribute dont_touch of WX9648: signal is true;
	signal WX9649: std_logic; attribute dont_touch of WX9649: signal is true;
	signal WX9650: std_logic; attribute dont_touch of WX9650: signal is true;
	signal WX9651: std_logic; attribute dont_touch of WX9651: signal is true;
	signal WX9652: std_logic; attribute dont_touch of WX9652: signal is true;
	signal WX9653: std_logic; attribute dont_touch of WX9653: signal is true;
	signal WX9654: std_logic; attribute dont_touch of WX9654: signal is true;
	signal WX9655: std_logic; attribute dont_touch of WX9655: signal is true;
	signal WX9656: std_logic; attribute dont_touch of WX9656: signal is true;
	signal WX9657: std_logic; attribute dont_touch of WX9657: signal is true;
	signal WX9658: std_logic; attribute dont_touch of WX9658: signal is true;
	signal WX9659: std_logic; attribute dont_touch of WX9659: signal is true;
	signal WX9660: std_logic; attribute dont_touch of WX9660: signal is true;
	signal WX9661: std_logic; attribute dont_touch of WX9661: signal is true;
	signal WX9662: std_logic; attribute dont_touch of WX9662: signal is true;
	signal WX9663: std_logic; attribute dont_touch of WX9663: signal is true;
	signal WX9664: std_logic; attribute dont_touch of WX9664: signal is true;
	signal WX9665: std_logic; attribute dont_touch of WX9665: signal is true;
	signal WX9666: std_logic; attribute dont_touch of WX9666: signal is true;
	signal WX9667: std_logic; attribute dont_touch of WX9667: signal is true;
	signal WX9668: std_logic; attribute dont_touch of WX9668: signal is true;
	signal WX9669: std_logic; attribute dont_touch of WX9669: signal is true;
	signal WX9670: std_logic; attribute dont_touch of WX9670: signal is true;
	signal WX9671: std_logic; attribute dont_touch of WX9671: signal is true;
	signal WX9672: std_logic; attribute dont_touch of WX9672: signal is true;
	signal WX9673: std_logic; attribute dont_touch of WX9673: signal is true;
	signal WX9674: std_logic; attribute dont_touch of WX9674: signal is true;
	signal WX9675: std_logic; attribute dont_touch of WX9675: signal is true;
	signal WX9676: std_logic; attribute dont_touch of WX9676: signal is true;
	signal WX9677: std_logic; attribute dont_touch of WX9677: signal is true;
	signal WX9678: std_logic; attribute dont_touch of WX9678: signal is true;
	signal WX9679: std_logic; attribute dont_touch of WX9679: signal is true;
	signal WX9680: std_logic; attribute dont_touch of WX9680: signal is true;
	signal WX9681: std_logic; attribute dont_touch of WX9681: signal is true;
	signal WX9682: std_logic; attribute dont_touch of WX9682: signal is true;
	signal WX9683: std_logic; attribute dont_touch of WX9683: signal is true;
	signal WX9684: std_logic; attribute dont_touch of WX9684: signal is true;
	signal WX9685: std_logic; attribute dont_touch of WX9685: signal is true;
	signal WX9686: std_logic; attribute dont_touch of WX9686: signal is true;
	signal WX9687: std_logic; attribute dont_touch of WX9687: signal is true;
	signal WX9688: std_logic; attribute dont_touch of WX9688: signal is true;
	signal WX9689: std_logic; attribute dont_touch of WX9689: signal is true;
	signal WX9690: std_logic; attribute dont_touch of WX9690: signal is true;
	signal WX9691: std_logic; attribute dont_touch of WX9691: signal is true;
	signal WX9692: std_logic; attribute dont_touch of WX9692: signal is true;
	signal WX9693: std_logic; attribute dont_touch of WX9693: signal is true;
	signal WX9694: std_logic; attribute dont_touch of WX9694: signal is true;
	signal WX9695: std_logic; attribute dont_touch of WX9695: signal is true;
	signal WX9696: std_logic; attribute dont_touch of WX9696: signal is true;
	signal WX9697: std_logic; attribute dont_touch of WX9697: signal is true;
	signal WX9698: std_logic; attribute dont_touch of WX9698: signal is true;
	signal WX9699: std_logic; attribute dont_touch of WX9699: signal is true;
	signal WX9700: std_logic; attribute dont_touch of WX9700: signal is true;
	signal WX9701: std_logic; attribute dont_touch of WX9701: signal is true;
	signal WX9702: std_logic; attribute dont_touch of WX9702: signal is true;
	signal WX9703: std_logic; attribute dont_touch of WX9703: signal is true;
	signal WX9704: std_logic; attribute dont_touch of WX9704: signal is true;
	signal WX9705: std_logic; attribute dont_touch of WX9705: signal is true;
	signal WX9706: std_logic; attribute dont_touch of WX9706: signal is true;
	signal WX9707: std_logic; attribute dont_touch of WX9707: signal is true;
	signal WX9708: std_logic; attribute dont_touch of WX9708: signal is true;
	signal WX9709: std_logic; attribute dont_touch of WX9709: signal is true;
	signal WX9710: std_logic; attribute dont_touch of WX9710: signal is true;
	signal WX9711: std_logic; attribute dont_touch of WX9711: signal is true;
	signal WX9712: std_logic; attribute dont_touch of WX9712: signal is true;
	signal WX9713: std_logic; attribute dont_touch of WX9713: signal is true;
	signal WX9714: std_logic; attribute dont_touch of WX9714: signal is true;
	signal WX9715: std_logic; attribute dont_touch of WX9715: signal is true;
	signal WX9716: std_logic; attribute dont_touch of WX9716: signal is true;
	signal WX9717: std_logic; attribute dont_touch of WX9717: signal is true;
	signal WX9718: std_logic; attribute dont_touch of WX9718: signal is true;
	signal WX9719: std_logic; attribute dont_touch of WX9719: signal is true;
	signal WX9720: std_logic; attribute dont_touch of WX9720: signal is true;
	signal WX9721: std_logic; attribute dont_touch of WX9721: signal is true;
	signal WX9722: std_logic; attribute dont_touch of WX9722: signal is true;
	signal WX9723: std_logic; attribute dont_touch of WX9723: signal is true;
	signal WX9724: std_logic; attribute dont_touch of WX9724: signal is true;
	signal WX9725: std_logic; attribute dont_touch of WX9725: signal is true;
	signal WX9726: std_logic; attribute dont_touch of WX9726: signal is true;
	signal WX9727: std_logic; attribute dont_touch of WX9727: signal is true;
	signal WX9728: std_logic; attribute dont_touch of WX9728: signal is true;
	signal WX9729: std_logic; attribute dont_touch of WX9729: signal is true;
	signal WX9730: std_logic; attribute dont_touch of WX9730: signal is true;
	signal WX9731: std_logic; attribute dont_touch of WX9731: signal is true;
	signal WX9732: std_logic; attribute dont_touch of WX9732: signal is true;
	signal WX9733: std_logic; attribute dont_touch of WX9733: signal is true;
	signal WX9734: std_logic; attribute dont_touch of WX9734: signal is true;
	signal WX9735: std_logic; attribute dont_touch of WX9735: signal is true;
	signal WX9736: std_logic; attribute dont_touch of WX9736: signal is true;
	signal WX9737: std_logic; attribute dont_touch of WX9737: signal is true;
	signal WX9738: std_logic; attribute dont_touch of WX9738: signal is true;
	signal WX9739: std_logic; attribute dont_touch of WX9739: signal is true;
	signal WX9740: std_logic; attribute dont_touch of WX9740: signal is true;
	signal WX9741: std_logic; attribute dont_touch of WX9741: signal is true;
	signal WX9742: std_logic; attribute dont_touch of WX9742: signal is true;
	signal WX9743: std_logic; attribute dont_touch of WX9743: signal is true;
	signal WX9744: std_logic; attribute dont_touch of WX9744: signal is true;
	signal WX9745: std_logic; attribute dont_touch of WX9745: signal is true;
	signal WX9746: std_logic; attribute dont_touch of WX9746: signal is true;
	signal WX9747: std_logic; attribute dont_touch of WX9747: signal is true;
	signal WX9748: std_logic; attribute dont_touch of WX9748: signal is true;
	signal WX9749: std_logic; attribute dont_touch of WX9749: signal is true;
	signal WX9750: std_logic; attribute dont_touch of WX9750: signal is true;
	signal WX9751: std_logic; attribute dont_touch of WX9751: signal is true;
	signal WX9752: std_logic; attribute dont_touch of WX9752: signal is true;
	signal WX9753: std_logic; attribute dont_touch of WX9753: signal is true;
	signal WX9754: std_logic; attribute dont_touch of WX9754: signal is true;
	signal WX9755: std_logic; attribute dont_touch of WX9755: signal is true;
	signal WX9756: std_logic; attribute dont_touch of WX9756: signal is true;
	signal WX9757: std_logic; attribute dont_touch of WX9757: signal is true;
	signal WX9758: std_logic; attribute dont_touch of WX9758: signal is true;
	signal WX9759: std_logic; attribute dont_touch of WX9759: signal is true;
	signal WX9760: std_logic; attribute dont_touch of WX9760: signal is true;
	signal WX9761: std_logic; attribute dont_touch of WX9761: signal is true;
	signal WX9762: std_logic; attribute dont_touch of WX9762: signal is true;
	signal WX9763: std_logic; attribute dont_touch of WX9763: signal is true;
	signal WX9764: std_logic; attribute dont_touch of WX9764: signal is true;
	signal WX9765: std_logic; attribute dont_touch of WX9765: signal is true;
	signal WX9766: std_logic; attribute dont_touch of WX9766: signal is true;
	signal WX9767: std_logic; attribute dont_touch of WX9767: signal is true;
	signal WX9768: std_logic; attribute dont_touch of WX9768: signal is true;
	signal WX9769: std_logic; attribute dont_touch of WX9769: signal is true;
	signal WX9770: std_logic; attribute dont_touch of WX9770: signal is true;
	signal WX9771: std_logic; attribute dont_touch of WX9771: signal is true;
	signal WX9772: std_logic; attribute dont_touch of WX9772: signal is true;
	signal WX9773: std_logic; attribute dont_touch of WX9773: signal is true;
	signal WX9774: std_logic; attribute dont_touch of WX9774: signal is true;
	signal WX9775: std_logic; attribute dont_touch of WX9775: signal is true;
	signal WX9776: std_logic; attribute dont_touch of WX9776: signal is true;
	signal WX9777: std_logic; attribute dont_touch of WX9777: signal is true;
	signal WX9778: std_logic; attribute dont_touch of WX9778: signal is true;
	signal WX9779: std_logic; attribute dont_touch of WX9779: signal is true;
	signal WX9780: std_logic; attribute dont_touch of WX9780: signal is true;
	signal WX9781: std_logic; attribute dont_touch of WX9781: signal is true;
	signal WX9782: std_logic; attribute dont_touch of WX9782: signal is true;
	signal WX9783: std_logic; attribute dont_touch of WX9783: signal is true;
	signal WX9784: std_logic; attribute dont_touch of WX9784: signal is true;
	signal WX9785: std_logic; attribute dont_touch of WX9785: signal is true;
	signal WX9786: std_logic; attribute dont_touch of WX9786: signal is true;
	signal WX9787: std_logic; attribute dont_touch of WX9787: signal is true;
	signal WX9788: std_logic; attribute dont_touch of WX9788: signal is true;
	signal WX9789: std_logic; attribute dont_touch of WX9789: signal is true;
	signal WX9790: std_logic; attribute dont_touch of WX9790: signal is true;
	signal WX9791: std_logic; attribute dont_touch of WX9791: signal is true;
	signal WX9792: std_logic; attribute dont_touch of WX9792: signal is true;
	signal WX9793: std_logic; attribute dont_touch of WX9793: signal is true;
	signal WX9794: std_logic; attribute dont_touch of WX9794: signal is true;
	signal WX9795: std_logic; attribute dont_touch of WX9795: signal is true;
	signal WX9796: std_logic; attribute dont_touch of WX9796: signal is true;
	signal WX9797: std_logic; attribute dont_touch of WX9797: signal is true;
	signal WX9798: std_logic; attribute dont_touch of WX9798: signal is true;
	signal WX9799: std_logic; attribute dont_touch of WX9799: signal is true;
	signal WX9800: std_logic; attribute dont_touch of WX9800: signal is true;
	signal WX9801: std_logic; attribute dont_touch of WX9801: signal is true;
	signal WX9802: std_logic; attribute dont_touch of WX9802: signal is true;
	signal WX9803: std_logic; attribute dont_touch of WX9803: signal is true;
	signal WX9804: std_logic; attribute dont_touch of WX9804: signal is true;
	signal WX9805: std_logic; attribute dont_touch of WX9805: signal is true;
	signal WX9806: std_logic; attribute dont_touch of WX9806: signal is true;
	signal WX9807: std_logic; attribute dont_touch of WX9807: signal is true;
	signal WX9808: std_logic; attribute dont_touch of WX9808: signal is true;
	signal WX9809: std_logic; attribute dont_touch of WX9809: signal is true;
	signal WX9810: std_logic; attribute dont_touch of WX9810: signal is true;
	signal WX9811: std_logic; attribute dont_touch of WX9811: signal is true;
	signal WX9812: std_logic; attribute dont_touch of WX9812: signal is true;
	signal WX9813: std_logic; attribute dont_touch of WX9813: signal is true;
	signal WX9814: std_logic; attribute dont_touch of WX9814: signal is true;
	signal WX9815: std_logic; attribute dont_touch of WX9815: signal is true;
	signal WX9816: std_logic; attribute dont_touch of WX9816: signal is true;
	signal WX9817: std_logic; attribute dont_touch of WX9817: signal is true;
	signal WX9818: std_logic; attribute dont_touch of WX9818: signal is true;
	signal WX9819: std_logic; attribute dont_touch of WX9819: signal is true;
	signal WX9820: std_logic; attribute dont_touch of WX9820: signal is true;
	signal WX9821: std_logic; attribute dont_touch of WX9821: signal is true;
	signal WX9822: std_logic; attribute dont_touch of WX9822: signal is true;
	signal WX9823: std_logic; attribute dont_touch of WX9823: signal is true;
	signal WX9824: std_logic; attribute dont_touch of WX9824: signal is true;
	signal WX9825: std_logic; attribute dont_touch of WX9825: signal is true;
	signal WX9826: std_logic; attribute dont_touch of WX9826: signal is true;
	signal WX9827: std_logic; attribute dont_touch of WX9827: signal is true;
	signal WX9828: std_logic; attribute dont_touch of WX9828: signal is true;
	signal WX9829: std_logic; attribute dont_touch of WX9829: signal is true;
	signal WX9830: std_logic; attribute dont_touch of WX9830: signal is true;
	signal WX9831: std_logic; attribute dont_touch of WX9831: signal is true;
	signal WX9832: std_logic; attribute dont_touch of WX9832: signal is true;
	signal WX9833: std_logic; attribute dont_touch of WX9833: signal is true;
	signal WX9834: std_logic; attribute dont_touch of WX9834: signal is true;
	signal WX9835: std_logic; attribute dont_touch of WX9835: signal is true;
	signal WX9836: std_logic; attribute dont_touch of WX9836: signal is true;
	signal WX9837: std_logic; attribute dont_touch of WX9837: signal is true;
	signal WX9838: std_logic; attribute dont_touch of WX9838: signal is true;
	signal WX9839: std_logic; attribute dont_touch of WX9839: signal is true;
	signal WX9840: std_logic; attribute dont_touch of WX9840: signal is true;
	signal WX9841: std_logic; attribute dont_touch of WX9841: signal is true;
	signal WX9842: std_logic; attribute dont_touch of WX9842: signal is true;
	signal WX9843: std_logic; attribute dont_touch of WX9843: signal is true;
	signal WX9844: std_logic; attribute dont_touch of WX9844: signal is true;
	signal WX9845: std_logic; attribute dont_touch of WX9845: signal is true;
	signal WX9846: std_logic; attribute dont_touch of WX9846: signal is true;
	signal WX9847: std_logic; attribute dont_touch of WX9847: signal is true;
	signal WX9848: std_logic; attribute dont_touch of WX9848: signal is true;
	signal WX9849: std_logic; attribute dont_touch of WX9849: signal is true;
	signal WX9850: std_logic; attribute dont_touch of WX9850: signal is true;
	signal WX9851: std_logic; attribute dont_touch of WX9851: signal is true;
	signal WX9852: std_logic; attribute dont_touch of WX9852: signal is true;
	signal WX9853: std_logic; attribute dont_touch of WX9853: signal is true;
	signal WX9854: std_logic; attribute dont_touch of WX9854: signal is true;
	signal WX9855: std_logic; attribute dont_touch of WX9855: signal is true;
	signal WX9856: std_logic; attribute dont_touch of WX9856: signal is true;
	signal WX9857: std_logic; attribute dont_touch of WX9857: signal is true;
	signal WX9858: std_logic; attribute dont_touch of WX9858: signal is true;
	signal WX9859: std_logic; attribute dont_touch of WX9859: signal is true;
	signal WX9860: std_logic; attribute dont_touch of WX9860: signal is true;
	signal WX9861: std_logic; attribute dont_touch of WX9861: signal is true;
	signal WX9862: std_logic; attribute dont_touch of WX9862: signal is true;
	signal WX9863: std_logic; attribute dont_touch of WX9863: signal is true;
	signal WX9864: std_logic; attribute dont_touch of WX9864: signal is true;
	signal WX9865: std_logic; attribute dont_touch of WX9865: signal is true;
	signal WX9866: std_logic; attribute dont_touch of WX9866: signal is true;
	signal WX9867: std_logic; attribute dont_touch of WX9867: signal is true;
	signal WX9868: std_logic; attribute dont_touch of WX9868: signal is true;
	signal WX9869: std_logic; attribute dont_touch of WX9869: signal is true;
	signal WX9870: std_logic; attribute dont_touch of WX9870: signal is true;
	signal WX9871: std_logic; attribute dont_touch of WX9871: signal is true;
	signal WX9872: std_logic; attribute dont_touch of WX9872: signal is true;
	signal WX9873: std_logic; attribute dont_touch of WX9873: signal is true;
	signal WX9874: std_logic; attribute dont_touch of WX9874: signal is true;
	signal WX9875: std_logic; attribute dont_touch of WX9875: signal is true;
	signal WX9876: std_logic; attribute dont_touch of WX9876: signal is true;
	signal WX9877: std_logic; attribute dont_touch of WX9877: signal is true;
	signal WX9878: std_logic; attribute dont_touch of WX9878: signal is true;
	signal WX9879: std_logic; attribute dont_touch of WX9879: signal is true;
	signal WX9880: std_logic; attribute dont_touch of WX9880: signal is true;
	signal WX9881: std_logic; attribute dont_touch of WX9881: signal is true;
	signal WX9882: std_logic; attribute dont_touch of WX9882: signal is true;
	signal WX9883: std_logic; attribute dont_touch of WX9883: signal is true;
	signal WX9884: std_logic; attribute dont_touch of WX9884: signal is true;
	signal WX9885: std_logic; attribute dont_touch of WX9885: signal is true;
	signal WX9886: std_logic; attribute dont_touch of WX9886: signal is true;
	signal WX9887: std_logic; attribute dont_touch of WX9887: signal is true;
	signal WX9888: std_logic; attribute dont_touch of WX9888: signal is true;
	signal WX9889: std_logic; attribute dont_touch of WX9889: signal is true;
	signal WX9890: std_logic; attribute dont_touch of WX9890: signal is true;
	signal WX9891: std_logic; attribute dont_touch of WX9891: signal is true;
	signal WX9892: std_logic; attribute dont_touch of WX9892: signal is true;
	signal WX9893: std_logic; attribute dont_touch of WX9893: signal is true;
	signal WX9894: std_logic; attribute dont_touch of WX9894: signal is true;
	signal WX9895: std_logic; attribute dont_touch of WX9895: signal is true;
	signal WX9896: std_logic; attribute dont_touch of WX9896: signal is true;
	signal WX9897: std_logic; attribute dont_touch of WX9897: signal is true;
	signal WX9898: std_logic; attribute dont_touch of WX9898: signal is true;
	signal WX9899: std_logic; attribute dont_touch of WX9899: signal is true;
	signal WX9900: std_logic; attribute dont_touch of WX9900: signal is true;
	signal WX9901: std_logic; attribute dont_touch of WX9901: signal is true;
	signal WX9902: std_logic; attribute dont_touch of WX9902: signal is true;
	signal WX9903: std_logic; attribute dont_touch of WX9903: signal is true;
	signal WX9904: std_logic; attribute dont_touch of WX9904: signal is true;
	signal WX9905: std_logic; attribute dont_touch of WX9905: signal is true;
	signal WX9906: std_logic; attribute dont_touch of WX9906: signal is true;
	signal WX9907: std_logic; attribute dont_touch of WX9907: signal is true;
	signal WX9908: std_logic; attribute dont_touch of WX9908: signal is true;
	signal WX9909: std_logic; attribute dont_touch of WX9909: signal is true;
	signal WX9910: std_logic; attribute dont_touch of WX9910: signal is true;
	signal WX9911: std_logic; attribute dont_touch of WX9911: signal is true;
	signal WX9912: std_logic; attribute dont_touch of WX9912: signal is true;
	signal WX9913: std_logic; attribute dont_touch of WX9913: signal is true;
	signal WX9914: std_logic; attribute dont_touch of WX9914: signal is true;
	signal WX9915: std_logic; attribute dont_touch of WX9915: signal is true;
	signal WX9916: std_logic; attribute dont_touch of WX9916: signal is true;
	signal WX9917: std_logic; attribute dont_touch of WX9917: signal is true;
	signal WX9918: std_logic; attribute dont_touch of WX9918: signal is true;
	signal WX9919: std_logic; attribute dont_touch of WX9919: signal is true;
	signal WX9920: std_logic; attribute dont_touch of WX9920: signal is true;
	signal WX9921: std_logic; attribute dont_touch of WX9921: signal is true;
	signal WX9922: std_logic; attribute dont_touch of WX9922: signal is true;
	signal WX9923: std_logic; attribute dont_touch of WX9923: signal is true;
	signal WX9924: std_logic; attribute dont_touch of WX9924: signal is true;
	signal WX9925: std_logic; attribute dont_touch of WX9925: signal is true;
	signal WX9926: std_logic; attribute dont_touch of WX9926: signal is true;
	signal WX9927: std_logic; attribute dont_touch of WX9927: signal is true;
	signal WX9928: std_logic; attribute dont_touch of WX9928: signal is true;
	signal WX9929: std_logic; attribute dont_touch of WX9929: signal is true;
	signal WX9930: std_logic; attribute dont_touch of WX9930: signal is true;
	signal WX9931: std_logic; attribute dont_touch of WX9931: signal is true;
	signal WX9932: std_logic; attribute dont_touch of WX9932: signal is true;
	signal WX9933: std_logic; attribute dont_touch of WX9933: signal is true;
	signal WX9934: std_logic; attribute dont_touch of WX9934: signal is true;
	signal WX9935: std_logic; attribute dont_touch of WX9935: signal is true;
	signal WX9936: std_logic; attribute dont_touch of WX9936: signal is true;
	signal WX9937: std_logic; attribute dont_touch of WX9937: signal is true;
	signal WX9938: std_logic; attribute dont_touch of WX9938: signal is true;
	signal WX9939: std_logic; attribute dont_touch of WX9939: signal is true;
	signal WX9940: std_logic; attribute dont_touch of WX9940: signal is true;
	signal WX9941: std_logic; attribute dont_touch of WX9941: signal is true;
	signal WX9942: std_logic; attribute dont_touch of WX9942: signal is true;
	signal WX9943: std_logic; attribute dont_touch of WX9943: signal is true;
	signal WX9944: std_logic; attribute dont_touch of WX9944: signal is true;
	signal WX9945: std_logic; attribute dont_touch of WX9945: signal is true;
	signal WX9946: std_logic; attribute dont_touch of WX9946: signal is true;
	signal WX9947: std_logic; attribute dont_touch of WX9947: signal is true;
	signal WX9948: std_logic; attribute dont_touch of WX9948: signal is true;
	signal WX9949: std_logic; attribute dont_touch of WX9949: signal is true;
	signal WX9950: std_logic; attribute dont_touch of WX9950: signal is true;
	signal WX9951: std_logic; attribute dont_touch of WX9951: signal is true;
	signal WX9952: std_logic; attribute dont_touch of WX9952: signal is true;
	signal WX9953: std_logic; attribute dont_touch of WX9953: signal is true;
	signal WX9954: std_logic; attribute dont_touch of WX9954: signal is true;
	signal WX9955: std_logic; attribute dont_touch of WX9955: signal is true;
	signal WX9956: std_logic; attribute dont_touch of WX9956: signal is true;
	signal WX9957: std_logic; attribute dont_touch of WX9957: signal is true;
	signal WX9958: std_logic; attribute dont_touch of WX9958: signal is true;
	signal WX9959: std_logic; attribute dont_touch of WX9959: signal is true;
	signal WX9960: std_logic; attribute dont_touch of WX9960: signal is true;
	signal WX9961: std_logic; attribute dont_touch of WX9961: signal is true;
	signal WX9962: std_logic; attribute dont_touch of WX9962: signal is true;
	signal WX9963: std_logic; attribute dont_touch of WX9963: signal is true;
	signal WX9964: std_logic; attribute dont_touch of WX9964: signal is true;
	signal WX9965: std_logic; attribute dont_touch of WX9965: signal is true;
	signal WX9966: std_logic; attribute dont_touch of WX9966: signal is true;
	signal WX9967: std_logic; attribute dont_touch of WX9967: signal is true;
	signal WX9968: std_logic; attribute dont_touch of WX9968: signal is true;
	signal WX9969: std_logic; attribute dont_touch of WX9969: signal is true;
	signal WX9970: std_logic; attribute dont_touch of WX9970: signal is true;
	signal WX9971: std_logic; attribute dont_touch of WX9971: signal is true;
	signal WX9972: std_logic; attribute dont_touch of WX9972: signal is true;
	signal WX9973: std_logic; attribute dont_touch of WX9973: signal is true;
	signal WX9974: std_logic; attribute dont_touch of WX9974: signal is true;
	signal WX9975: std_logic; attribute dont_touch of WX9975: signal is true;
	signal WX9976: std_logic; attribute dont_touch of WX9976: signal is true;
	signal WX9977: std_logic; attribute dont_touch of WX9977: signal is true;
	signal WX9978: std_logic; attribute dont_touch of WX9978: signal is true;
	signal WX9979: std_logic; attribute dont_touch of WX9979: signal is true;
	signal WX9980: std_logic; attribute dont_touch of WX9980: signal is true;
	signal WX9981: std_logic; attribute dont_touch of WX9981: signal is true;
	signal WX9982: std_logic; attribute dont_touch of WX9982: signal is true;
	signal WX9983: std_logic; attribute dont_touch of WX9983: signal is true;
	signal WX9984: std_logic; attribute dont_touch of WX9984: signal is true;
	signal WX9985: std_logic; attribute dont_touch of WX9985: signal is true;
	signal WX9986: std_logic; attribute dont_touch of WX9986: signal is true;
	signal WX9987: std_logic; attribute dont_touch of WX9987: signal is true;
	signal WX9988: std_logic; attribute dont_touch of WX9988: signal is true;
	signal WX9989: std_logic; attribute dont_touch of WX9989: signal is true;
	signal WX9990: std_logic; attribute dont_touch of WX9990: signal is true;
	signal WX9991: std_logic; attribute dont_touch of WX9991: signal is true;
	signal WX9992: std_logic; attribute dont_touch of WX9992: signal is true;
	signal WX9993: std_logic; attribute dont_touch of WX9993: signal is true;
	signal WX9994: std_logic; attribute dont_touch of WX9994: signal is true;
	signal WX9995: std_logic; attribute dont_touch of WX9995: signal is true;
	signal WX9996: std_logic; attribute dont_touch of WX9996: signal is true;
	signal WX9997: std_logic; attribute dont_touch of WX9997: signal is true;
	signal WX9998: std_logic; attribute dont_touch of WX9998: signal is true;
	signal WX9999: std_logic; attribute dont_touch of WX9999: signal is true;
	signal WX10000: std_logic; attribute dont_touch of WX10000: signal is true;
	signal WX10001: std_logic; attribute dont_touch of WX10001: signal is true;
	signal WX10002: std_logic; attribute dont_touch of WX10002: signal is true;
	signal WX10003: std_logic; attribute dont_touch of WX10003: signal is true;
	signal WX10004: std_logic; attribute dont_touch of WX10004: signal is true;
	signal WX10005: std_logic; attribute dont_touch of WX10005: signal is true;
	signal WX10006: std_logic; attribute dont_touch of WX10006: signal is true;
	signal WX10007: std_logic; attribute dont_touch of WX10007: signal is true;
	signal WX10008: std_logic; attribute dont_touch of WX10008: signal is true;
	signal WX10009: std_logic; attribute dont_touch of WX10009: signal is true;
	signal WX10010: std_logic; attribute dont_touch of WX10010: signal is true;
	signal WX10011: std_logic; attribute dont_touch of WX10011: signal is true;
	signal WX10012: std_logic; attribute dont_touch of WX10012: signal is true;
	signal WX10013: std_logic; attribute dont_touch of WX10013: signal is true;
	signal WX10014: std_logic; attribute dont_touch of WX10014: signal is true;
	signal WX10015: std_logic; attribute dont_touch of WX10015: signal is true;
	signal WX10016: std_logic; attribute dont_touch of WX10016: signal is true;
	signal WX10017: std_logic; attribute dont_touch of WX10017: signal is true;
	signal WX10018: std_logic; attribute dont_touch of WX10018: signal is true;
	signal WX10019: std_logic; attribute dont_touch of WX10019: signal is true;
	signal WX10020: std_logic; attribute dont_touch of WX10020: signal is true;
	signal WX10021: std_logic; attribute dont_touch of WX10021: signal is true;
	signal WX10022: std_logic; attribute dont_touch of WX10022: signal is true;
	signal WX10023: std_logic; attribute dont_touch of WX10023: signal is true;
	signal WX10024: std_logic; attribute dont_touch of WX10024: signal is true;
	signal WX10025: std_logic; attribute dont_touch of WX10025: signal is true;
	signal WX10026: std_logic; attribute dont_touch of WX10026: signal is true;
	signal WX10027: std_logic; attribute dont_touch of WX10027: signal is true;
	signal WX10028: std_logic; attribute dont_touch of WX10028: signal is true;
	signal WX10029: std_logic; attribute dont_touch of WX10029: signal is true;
	signal WX10030: std_logic; attribute dont_touch of WX10030: signal is true;
	signal WX10031: std_logic; attribute dont_touch of WX10031: signal is true;
	signal WX10032: std_logic; attribute dont_touch of WX10032: signal is true;
	signal WX10033: std_logic; attribute dont_touch of WX10033: signal is true;
	signal WX10034: std_logic; attribute dont_touch of WX10034: signal is true;
	signal WX10035: std_logic; attribute dont_touch of WX10035: signal is true;
	signal WX10036: std_logic; attribute dont_touch of WX10036: signal is true;
	signal WX10037: std_logic; attribute dont_touch of WX10037: signal is true;
	signal WX10038: std_logic; attribute dont_touch of WX10038: signal is true;
	signal WX10039: std_logic; attribute dont_touch of WX10039: signal is true;
	signal WX10040: std_logic; attribute dont_touch of WX10040: signal is true;
	signal WX10041: std_logic; attribute dont_touch of WX10041: signal is true;
	signal WX10042: std_logic; attribute dont_touch of WX10042: signal is true;
	signal WX10043: std_logic; attribute dont_touch of WX10043: signal is true;
	signal WX10044: std_logic; attribute dont_touch of WX10044: signal is true;
	signal WX10045: std_logic; attribute dont_touch of WX10045: signal is true;
	signal WX10046: std_logic; attribute dont_touch of WX10046: signal is true;
	signal WX10047: std_logic; attribute dont_touch of WX10047: signal is true;
	signal WX10048: std_logic; attribute dont_touch of WX10048: signal is true;
	signal WX10049: std_logic; attribute dont_touch of WX10049: signal is true;
	signal WX10050: std_logic; attribute dont_touch of WX10050: signal is true;
	signal WX10051: std_logic; attribute dont_touch of WX10051: signal is true;
	signal WX10052: std_logic; attribute dont_touch of WX10052: signal is true;
	signal WX10053: std_logic; attribute dont_touch of WX10053: signal is true;
	signal WX10054: std_logic; attribute dont_touch of WX10054: signal is true;
	signal WX10055: std_logic; attribute dont_touch of WX10055: signal is true;
	signal WX10056: std_logic; attribute dont_touch of WX10056: signal is true;
	signal WX10057: std_logic; attribute dont_touch of WX10057: signal is true;
	signal WX10058: std_logic; attribute dont_touch of WX10058: signal is true;
	signal WX10059: std_logic; attribute dont_touch of WX10059: signal is true;
	signal WX10060: std_logic; attribute dont_touch of WX10060: signal is true;
	signal WX10061: std_logic; attribute dont_touch of WX10061: signal is true;
	signal WX10062: std_logic; attribute dont_touch of WX10062: signal is true;
	signal WX10063: std_logic; attribute dont_touch of WX10063: signal is true;
	signal WX10064: std_logic; attribute dont_touch of WX10064: signal is true;
	signal WX10065: std_logic; attribute dont_touch of WX10065: signal is true;
	signal WX10066: std_logic; attribute dont_touch of WX10066: signal is true;
	signal WX10067: std_logic; attribute dont_touch of WX10067: signal is true;
	signal WX10068: std_logic; attribute dont_touch of WX10068: signal is true;
	signal WX10069: std_logic; attribute dont_touch of WX10069: signal is true;
	signal WX10070: std_logic; attribute dont_touch of WX10070: signal is true;
	signal WX10071: std_logic; attribute dont_touch of WX10071: signal is true;
	signal WX10072: std_logic; attribute dont_touch of WX10072: signal is true;
	signal WX10073: std_logic; attribute dont_touch of WX10073: signal is true;
	signal WX10074: std_logic; attribute dont_touch of WX10074: signal is true;
	signal WX10075: std_logic; attribute dont_touch of WX10075: signal is true;
	signal WX10076: std_logic; attribute dont_touch of WX10076: signal is true;
	signal WX10077: std_logic; attribute dont_touch of WX10077: signal is true;
	signal WX10078: std_logic; attribute dont_touch of WX10078: signal is true;
	signal WX10079: std_logic; attribute dont_touch of WX10079: signal is true;
	signal WX10080: std_logic; attribute dont_touch of WX10080: signal is true;
	signal WX10081: std_logic; attribute dont_touch of WX10081: signal is true;
	signal WX10082: std_logic; attribute dont_touch of WX10082: signal is true;
	signal WX10083: std_logic; attribute dont_touch of WX10083: signal is true;
	signal WX10084: std_logic; attribute dont_touch of WX10084: signal is true;
	signal WX10085: std_logic; attribute dont_touch of WX10085: signal is true;
	signal WX10086: std_logic; attribute dont_touch of WX10086: signal is true;
	signal WX10087: std_logic; attribute dont_touch of WX10087: signal is true;
	signal WX10088: std_logic; attribute dont_touch of WX10088: signal is true;
	signal WX10089: std_logic; attribute dont_touch of WX10089: signal is true;
	signal WX10090: std_logic; attribute dont_touch of WX10090: signal is true;
	signal WX10091: std_logic; attribute dont_touch of WX10091: signal is true;
	signal WX10092: std_logic; attribute dont_touch of WX10092: signal is true;
	signal WX10093: std_logic; attribute dont_touch of WX10093: signal is true;
	signal WX10094: std_logic; attribute dont_touch of WX10094: signal is true;
	signal WX10095: std_logic; attribute dont_touch of WX10095: signal is true;
	signal WX10096: std_logic; attribute dont_touch of WX10096: signal is true;
	signal WX10097: std_logic; attribute dont_touch of WX10097: signal is true;
	signal WX10098: std_logic; attribute dont_touch of WX10098: signal is true;
	signal WX10099: std_logic; attribute dont_touch of WX10099: signal is true;
	signal WX10100: std_logic; attribute dont_touch of WX10100: signal is true;
	signal WX10101: std_logic; attribute dont_touch of WX10101: signal is true;
	signal WX10102: std_logic; attribute dont_touch of WX10102: signal is true;
	signal WX10103: std_logic; attribute dont_touch of WX10103: signal is true;
	signal WX10104: std_logic; attribute dont_touch of WX10104: signal is true;
	signal WX10105: std_logic; attribute dont_touch of WX10105: signal is true;
	signal WX10106: std_logic; attribute dont_touch of WX10106: signal is true;
	signal WX10107: std_logic; attribute dont_touch of WX10107: signal is true;
	signal WX10108: std_logic; attribute dont_touch of WX10108: signal is true;
	signal WX10109: std_logic; attribute dont_touch of WX10109: signal is true;
	signal WX10110: std_logic; attribute dont_touch of WX10110: signal is true;
	signal WX10111: std_logic; attribute dont_touch of WX10111: signal is true;
	signal WX10112: std_logic; attribute dont_touch of WX10112: signal is true;
	signal WX10113: std_logic; attribute dont_touch of WX10113: signal is true;
	signal WX10114: std_logic; attribute dont_touch of WX10114: signal is true;
	signal WX10115: std_logic; attribute dont_touch of WX10115: signal is true;
	signal WX10116: std_logic; attribute dont_touch of WX10116: signal is true;
	signal WX10117: std_logic; attribute dont_touch of WX10117: signal is true;
	signal WX10118: std_logic; attribute dont_touch of WX10118: signal is true;
	signal WX10119: std_logic; attribute dont_touch of WX10119: signal is true;
	signal WX10120: std_logic; attribute dont_touch of WX10120: signal is true;
	signal WX10121: std_logic; attribute dont_touch of WX10121: signal is true;
	signal WX10122: std_logic; attribute dont_touch of WX10122: signal is true;
	signal WX10123: std_logic; attribute dont_touch of WX10123: signal is true;
	signal WX10124: std_logic; attribute dont_touch of WX10124: signal is true;
	signal WX10125: std_logic; attribute dont_touch of WX10125: signal is true;
	signal WX10126: std_logic; attribute dont_touch of WX10126: signal is true;
	signal WX10127: std_logic; attribute dont_touch of WX10127: signal is true;
	signal WX10128: std_logic; attribute dont_touch of WX10128: signal is true;
	signal WX10129: std_logic; attribute dont_touch of WX10129: signal is true;
	signal WX10130: std_logic; attribute dont_touch of WX10130: signal is true;
	signal WX10131: std_logic; attribute dont_touch of WX10131: signal is true;
	signal WX10132: std_logic; attribute dont_touch of WX10132: signal is true;
	signal WX10133: std_logic; attribute dont_touch of WX10133: signal is true;
	signal WX10134: std_logic; attribute dont_touch of WX10134: signal is true;
	signal WX10135: std_logic; attribute dont_touch of WX10135: signal is true;
	signal WX10136: std_logic; attribute dont_touch of WX10136: signal is true;
	signal WX10137: std_logic; attribute dont_touch of WX10137: signal is true;
	signal WX10138: std_logic; attribute dont_touch of WX10138: signal is true;
	signal WX10139: std_logic; attribute dont_touch of WX10139: signal is true;
	signal WX10140: std_logic; attribute dont_touch of WX10140: signal is true;
	signal WX10141: std_logic; attribute dont_touch of WX10141: signal is true;
	signal WX10142: std_logic; attribute dont_touch of WX10142: signal is true;
	signal WX10143: std_logic; attribute dont_touch of WX10143: signal is true;
	signal WX10144: std_logic; attribute dont_touch of WX10144: signal is true;
	signal WX10145: std_logic; attribute dont_touch of WX10145: signal is true;
	signal WX10146: std_logic; attribute dont_touch of WX10146: signal is true;
	signal WX10147: std_logic; attribute dont_touch of WX10147: signal is true;
	signal WX10148: std_logic; attribute dont_touch of WX10148: signal is true;
	signal WX10149: std_logic; attribute dont_touch of WX10149: signal is true;
	signal WX10150: std_logic; attribute dont_touch of WX10150: signal is true;
	signal WX10151: std_logic; attribute dont_touch of WX10151: signal is true;
	signal WX10152: std_logic; attribute dont_touch of WX10152: signal is true;
	signal WX10153: std_logic; attribute dont_touch of WX10153: signal is true;
	signal WX10154: std_logic; attribute dont_touch of WX10154: signal is true;
	signal WX10155: std_logic; attribute dont_touch of WX10155: signal is true;
	signal WX10156: std_logic; attribute dont_touch of WX10156: signal is true;
	signal WX10157: std_logic; attribute dont_touch of WX10157: signal is true;
	signal WX10158: std_logic; attribute dont_touch of WX10158: signal is true;
	signal WX10159: std_logic; attribute dont_touch of WX10159: signal is true;
	signal WX10160: std_logic; attribute dont_touch of WX10160: signal is true;
	signal WX10161: std_logic; attribute dont_touch of WX10161: signal is true;
	signal WX10162: std_logic; attribute dont_touch of WX10162: signal is true;
	signal WX10163: std_logic; attribute dont_touch of WX10163: signal is true;
	signal WX10164: std_logic; attribute dont_touch of WX10164: signal is true;
	signal WX10165: std_logic; attribute dont_touch of WX10165: signal is true;
	signal WX10166: std_logic; attribute dont_touch of WX10166: signal is true;
	signal WX10167: std_logic; attribute dont_touch of WX10167: signal is true;
	signal WX10168: std_logic; attribute dont_touch of WX10168: signal is true;
	signal WX10169: std_logic; attribute dont_touch of WX10169: signal is true;
	signal WX10170: std_logic; attribute dont_touch of WX10170: signal is true;
	signal WX10171: std_logic; attribute dont_touch of WX10171: signal is true;
	signal WX10172: std_logic; attribute dont_touch of WX10172: signal is true;
	signal WX10173: std_logic; attribute dont_touch of WX10173: signal is true;
	signal WX10174: std_logic; attribute dont_touch of WX10174: signal is true;
	signal WX10175: std_logic; attribute dont_touch of WX10175: signal is true;
	signal WX10176: std_logic; attribute dont_touch of WX10176: signal is true;
	signal WX10177: std_logic; attribute dont_touch of WX10177: signal is true;
	signal WX10178: std_logic; attribute dont_touch of WX10178: signal is true;
	signal WX10179: std_logic; attribute dont_touch of WX10179: signal is true;
	signal WX10180: std_logic; attribute dont_touch of WX10180: signal is true;
	signal WX10181: std_logic; attribute dont_touch of WX10181: signal is true;
	signal WX10182: std_logic; attribute dont_touch of WX10182: signal is true;
	signal WX10183: std_logic; attribute dont_touch of WX10183: signal is true;
	signal WX10184: std_logic; attribute dont_touch of WX10184: signal is true;
	signal WX10185: std_logic; attribute dont_touch of WX10185: signal is true;
	signal WX10186: std_logic; attribute dont_touch of WX10186: signal is true;
	signal WX10187: std_logic; attribute dont_touch of WX10187: signal is true;
	signal WX10188: std_logic; attribute dont_touch of WX10188: signal is true;
	signal WX10189: std_logic; attribute dont_touch of WX10189: signal is true;
	signal WX10190: std_logic; attribute dont_touch of WX10190: signal is true;
	signal WX10191: std_logic; attribute dont_touch of WX10191: signal is true;
	signal WX10192: std_logic; attribute dont_touch of WX10192: signal is true;
	signal WX10193: std_logic; attribute dont_touch of WX10193: signal is true;
	signal WX10194: std_logic; attribute dont_touch of WX10194: signal is true;
	signal WX10195: std_logic; attribute dont_touch of WX10195: signal is true;
	signal WX10196: std_logic; attribute dont_touch of WX10196: signal is true;
	signal WX10197: std_logic; attribute dont_touch of WX10197: signal is true;
	signal WX10198: std_logic; attribute dont_touch of WX10198: signal is true;
	signal WX10199: std_logic; attribute dont_touch of WX10199: signal is true;
	signal WX10200: std_logic; attribute dont_touch of WX10200: signal is true;
	signal WX10201: std_logic; attribute dont_touch of WX10201: signal is true;
	signal WX10202: std_logic; attribute dont_touch of WX10202: signal is true;
	signal WX10203: std_logic; attribute dont_touch of WX10203: signal is true;
	signal WX10204: std_logic; attribute dont_touch of WX10204: signal is true;
	signal WX10205: std_logic; attribute dont_touch of WX10205: signal is true;
	signal WX10206: std_logic; attribute dont_touch of WX10206: signal is true;
	signal WX10207: std_logic; attribute dont_touch of WX10207: signal is true;
	signal WX10208: std_logic; attribute dont_touch of WX10208: signal is true;
	signal WX10209: std_logic; attribute dont_touch of WX10209: signal is true;
	signal WX10210: std_logic; attribute dont_touch of WX10210: signal is true;
	signal WX10211: std_logic; attribute dont_touch of WX10211: signal is true;
	signal WX10212: std_logic; attribute dont_touch of WX10212: signal is true;
	signal WX10213: std_logic; attribute dont_touch of WX10213: signal is true;
	signal WX10214: std_logic; attribute dont_touch of WX10214: signal is true;
	signal WX10215: std_logic; attribute dont_touch of WX10215: signal is true;
	signal WX10216: std_logic; attribute dont_touch of WX10216: signal is true;
	signal WX10217: std_logic; attribute dont_touch of WX10217: signal is true;
	signal WX10218: std_logic; attribute dont_touch of WX10218: signal is true;
	signal WX10219: std_logic; attribute dont_touch of WX10219: signal is true;
	signal WX10220: std_logic; attribute dont_touch of WX10220: signal is true;
	signal WX10221: std_logic; attribute dont_touch of WX10221: signal is true;
	signal WX10222: std_logic; attribute dont_touch of WX10222: signal is true;
	signal WX10223: std_logic; attribute dont_touch of WX10223: signal is true;
	signal WX10224: std_logic; attribute dont_touch of WX10224: signal is true;
	signal WX10225: std_logic; attribute dont_touch of WX10225: signal is true;
	signal WX10226: std_logic; attribute dont_touch of WX10226: signal is true;
	signal WX10227: std_logic; attribute dont_touch of WX10227: signal is true;
	signal WX10228: std_logic; attribute dont_touch of WX10228: signal is true;
	signal WX10229: std_logic; attribute dont_touch of WX10229: signal is true;
	signal WX10230: std_logic; attribute dont_touch of WX10230: signal is true;
	signal WX10231: std_logic; attribute dont_touch of WX10231: signal is true;
	signal WX10232: std_logic; attribute dont_touch of WX10232: signal is true;
	signal WX10233: std_logic; attribute dont_touch of WX10233: signal is true;
	signal WX10234: std_logic; attribute dont_touch of WX10234: signal is true;
	signal WX10235: std_logic; attribute dont_touch of WX10235: signal is true;
	signal WX10236: std_logic; attribute dont_touch of WX10236: signal is true;
	signal WX10237: std_logic; attribute dont_touch of WX10237: signal is true;
	signal WX10238: std_logic; attribute dont_touch of WX10238: signal is true;
	signal WX10239: std_logic; attribute dont_touch of WX10239: signal is true;
	signal WX10240: std_logic; attribute dont_touch of WX10240: signal is true;
	signal WX10241: std_logic; attribute dont_touch of WX10241: signal is true;
	signal WX10242: std_logic; attribute dont_touch of WX10242: signal is true;
	signal WX10243: std_logic; attribute dont_touch of WX10243: signal is true;
	signal WX10244: std_logic; attribute dont_touch of WX10244: signal is true;
	signal WX10245: std_logic; attribute dont_touch of WX10245: signal is true;
	signal WX10246: std_logic; attribute dont_touch of WX10246: signal is true;
	signal WX10247: std_logic; attribute dont_touch of WX10247: signal is true;
	signal WX10248: std_logic; attribute dont_touch of WX10248: signal is true;
	signal WX10249: std_logic; attribute dont_touch of WX10249: signal is true;
	signal WX10250: std_logic; attribute dont_touch of WX10250: signal is true;
	signal WX10251: std_logic; attribute dont_touch of WX10251: signal is true;
	signal WX10252: std_logic; attribute dont_touch of WX10252: signal is true;
	signal WX10253: std_logic; attribute dont_touch of WX10253: signal is true;
	signal WX10254: std_logic; attribute dont_touch of WX10254: signal is true;
	signal WX10255: std_logic; attribute dont_touch of WX10255: signal is true;
	signal WX10256: std_logic; attribute dont_touch of WX10256: signal is true;
	signal WX10257: std_logic; attribute dont_touch of WX10257: signal is true;
	signal WX10258: std_logic; attribute dont_touch of WX10258: signal is true;
	signal WX10259: std_logic; attribute dont_touch of WX10259: signal is true;
	signal WX10260: std_logic; attribute dont_touch of WX10260: signal is true;
	signal WX10261: std_logic; attribute dont_touch of WX10261: signal is true;
	signal WX10262: std_logic; attribute dont_touch of WX10262: signal is true;
	signal WX10263: std_logic; attribute dont_touch of WX10263: signal is true;
	signal WX10264: std_logic; attribute dont_touch of WX10264: signal is true;
	signal WX10265: std_logic; attribute dont_touch of WX10265: signal is true;
	signal WX10266: std_logic; attribute dont_touch of WX10266: signal is true;
	signal WX10267: std_logic; attribute dont_touch of WX10267: signal is true;
	signal WX10268: std_logic; attribute dont_touch of WX10268: signal is true;
	signal WX10269: std_logic; attribute dont_touch of WX10269: signal is true;
	signal WX10270: std_logic; attribute dont_touch of WX10270: signal is true;
	signal WX10271: std_logic; attribute dont_touch of WX10271: signal is true;
	signal WX10272: std_logic; attribute dont_touch of WX10272: signal is true;
	signal WX10273: std_logic; attribute dont_touch of WX10273: signal is true;
	signal WX10274: std_logic; attribute dont_touch of WX10274: signal is true;
	signal WX10275: std_logic; attribute dont_touch of WX10275: signal is true;
	signal WX10276: std_logic; attribute dont_touch of WX10276: signal is true;
	signal WX10277: std_logic; attribute dont_touch of WX10277: signal is true;
	signal WX10278: std_logic; attribute dont_touch of WX10278: signal is true;
	signal WX10279: std_logic; attribute dont_touch of WX10279: signal is true;
	signal WX10280: std_logic; attribute dont_touch of WX10280: signal is true;
	signal WX10281: std_logic; attribute dont_touch of WX10281: signal is true;
	signal WX10282: std_logic; attribute dont_touch of WX10282: signal is true;
	signal WX10283: std_logic; attribute dont_touch of WX10283: signal is true;
	signal WX10284: std_logic; attribute dont_touch of WX10284: signal is true;
	signal WX10285: std_logic; attribute dont_touch of WX10285: signal is true;
	signal WX10286: std_logic; attribute dont_touch of WX10286: signal is true;
	signal WX10287: std_logic; attribute dont_touch of WX10287: signal is true;
	signal WX10288: std_logic; attribute dont_touch of WX10288: signal is true;
	signal WX10289: std_logic; attribute dont_touch of WX10289: signal is true;
	signal WX10290: std_logic; attribute dont_touch of WX10290: signal is true;
	signal WX10291: std_logic; attribute dont_touch of WX10291: signal is true;
	signal WX10292: std_logic; attribute dont_touch of WX10292: signal is true;
	signal WX10293: std_logic; attribute dont_touch of WX10293: signal is true;
	signal WX10294: std_logic; attribute dont_touch of WX10294: signal is true;
	signal WX10295: std_logic; attribute dont_touch of WX10295: signal is true;
	signal WX10296: std_logic; attribute dont_touch of WX10296: signal is true;
	signal WX10297: std_logic; attribute dont_touch of WX10297: signal is true;
	signal WX10298: std_logic; attribute dont_touch of WX10298: signal is true;
	signal WX10299: std_logic; attribute dont_touch of WX10299: signal is true;
	signal WX10300: std_logic; attribute dont_touch of WX10300: signal is true;
	signal WX10301: std_logic; attribute dont_touch of WX10301: signal is true;
	signal WX10302: std_logic; attribute dont_touch of WX10302: signal is true;
	signal WX10303: std_logic; attribute dont_touch of WX10303: signal is true;
	signal WX10304: std_logic; attribute dont_touch of WX10304: signal is true;
	signal WX10305: std_logic; attribute dont_touch of WX10305: signal is true;
	signal WX10306: std_logic; attribute dont_touch of WX10306: signal is true;
	signal WX10307: std_logic; attribute dont_touch of WX10307: signal is true;
	signal WX10308: std_logic; attribute dont_touch of WX10308: signal is true;
	signal WX10309: std_logic; attribute dont_touch of WX10309: signal is true;
	signal WX10310: std_logic; attribute dont_touch of WX10310: signal is true;
	signal WX10311: std_logic; attribute dont_touch of WX10311: signal is true;
	signal WX10312: std_logic; attribute dont_touch of WX10312: signal is true;
	signal WX10313: std_logic; attribute dont_touch of WX10313: signal is true;
	signal WX10314: std_logic; attribute dont_touch of WX10314: signal is true;
	signal WX10315: std_logic; attribute dont_touch of WX10315: signal is true;
	signal WX10317: std_logic; attribute dont_touch of WX10317: signal is true;
	signal WX10319: std_logic; attribute dont_touch of WX10319: signal is true;
	signal WX10321: std_logic; attribute dont_touch of WX10321: signal is true;
	signal WX10323: std_logic; attribute dont_touch of WX10323: signal is true;
	signal WX10325: std_logic; attribute dont_touch of WX10325: signal is true;
	signal WX10327: std_logic; attribute dont_touch of WX10327: signal is true;
	signal WX10329: std_logic; attribute dont_touch of WX10329: signal is true;
	signal WX10331: std_logic; attribute dont_touch of WX10331: signal is true;
	signal WX10333: std_logic; attribute dont_touch of WX10333: signal is true;
	signal WX10335: std_logic; attribute dont_touch of WX10335: signal is true;
	signal WX10337: std_logic; attribute dont_touch of WX10337: signal is true;
	signal WX10339: std_logic; attribute dont_touch of WX10339: signal is true;
	signal WX10341: std_logic; attribute dont_touch of WX10341: signal is true;
	signal WX10343: std_logic; attribute dont_touch of WX10343: signal is true;
	signal WX10345: std_logic; attribute dont_touch of WX10345: signal is true;
	signal WX10347: std_logic; attribute dont_touch of WX10347: signal is true;
	signal WX10349: std_logic; attribute dont_touch of WX10349: signal is true;
	signal WX10351: std_logic; attribute dont_touch of WX10351: signal is true;
	signal WX10353: std_logic; attribute dont_touch of WX10353: signal is true;
	signal WX10355: std_logic; attribute dont_touch of WX10355: signal is true;
	signal WX10357: std_logic; attribute dont_touch of WX10357: signal is true;
	signal WX10359: std_logic; attribute dont_touch of WX10359: signal is true;
	signal WX10361: std_logic; attribute dont_touch of WX10361: signal is true;
	signal WX10363: std_logic; attribute dont_touch of WX10363: signal is true;
	signal WX10365: std_logic; attribute dont_touch of WX10365: signal is true;
	signal WX10367: std_logic; attribute dont_touch of WX10367: signal is true;
	signal WX10369: std_logic; attribute dont_touch of WX10369: signal is true;
	signal WX10371: std_logic; attribute dont_touch of WX10371: signal is true;
	signal WX10373: std_logic; attribute dont_touch of WX10373: signal is true;
	signal WX10375: std_logic; attribute dont_touch of WX10375: signal is true;
	signal WX10377: std_logic; attribute dont_touch of WX10377: signal is true;
	signal WX10379: std_logic; attribute dont_touch of WX10379: signal is true;
	signal WX10380: std_logic; attribute dont_touch of WX10380: signal is true;
	signal WX10381: std_logic; attribute dont_touch of WX10381: signal is true;
	signal WX10382: std_logic; attribute dont_touch of WX10382: signal is true;
	signal WX10383: std_logic; attribute dont_touch of WX10383: signal is true;
	signal WX10384: std_logic; attribute dont_touch of WX10384: signal is true;
	signal WX10385: std_logic; attribute dont_touch of WX10385: signal is true;
	signal WX10386: std_logic; attribute dont_touch of WX10386: signal is true;
	signal WX10387: std_logic; attribute dont_touch of WX10387: signal is true;
	signal WX10388: std_logic; attribute dont_touch of WX10388: signal is true;
	signal WX10389: std_logic; attribute dont_touch of WX10389: signal is true;
	signal WX10390: std_logic; attribute dont_touch of WX10390: signal is true;
	signal WX10391: std_logic; attribute dont_touch of WX10391: signal is true;
	signal WX10392: std_logic; attribute dont_touch of WX10392: signal is true;
	signal WX10393: std_logic; attribute dont_touch of WX10393: signal is true;
	signal WX10394: std_logic; attribute dont_touch of WX10394: signal is true;
	signal WX10395: std_logic; attribute dont_touch of WX10395: signal is true;
	signal WX10396: std_logic; attribute dont_touch of WX10396: signal is true;
	signal WX10397: std_logic; attribute dont_touch of WX10397: signal is true;
	signal WX10398: std_logic; attribute dont_touch of WX10398: signal is true;
	signal WX10399: std_logic; attribute dont_touch of WX10399: signal is true;
	signal WX10400: std_logic; attribute dont_touch of WX10400: signal is true;
	signal WX10401: std_logic; attribute dont_touch of WX10401: signal is true;
	signal WX10402: std_logic; attribute dont_touch of WX10402: signal is true;
	signal WX10403: std_logic; attribute dont_touch of WX10403: signal is true;
	signal WX10404: std_logic; attribute dont_touch of WX10404: signal is true;
	signal WX10405: std_logic; attribute dont_touch of WX10405: signal is true;
	signal WX10406: std_logic; attribute dont_touch of WX10406: signal is true;
	signal WX10407: std_logic; attribute dont_touch of WX10407: signal is true;
	signal WX10408: std_logic; attribute dont_touch of WX10408: signal is true;
	signal WX10409: std_logic; attribute dont_touch of WX10409: signal is true;
	signal WX10410: std_logic; attribute dont_touch of WX10410: signal is true;
	signal WX10411: std_logic; attribute dont_touch of WX10411: signal is true;
	signal WX10412: std_logic; attribute dont_touch of WX10412: signal is true;
	signal WX10413: std_logic; attribute dont_touch of WX10413: signal is true;
	signal WX10414: std_logic; attribute dont_touch of WX10414: signal is true;
	signal WX10415: std_logic; attribute dont_touch of WX10415: signal is true;
	signal WX10416: std_logic; attribute dont_touch of WX10416: signal is true;
	signal WX10417: std_logic; attribute dont_touch of WX10417: signal is true;
	signal WX10418: std_logic; attribute dont_touch of WX10418: signal is true;
	signal WX10419: std_logic; attribute dont_touch of WX10419: signal is true;
	signal WX10420: std_logic; attribute dont_touch of WX10420: signal is true;
	signal WX10421: std_logic; attribute dont_touch of WX10421: signal is true;
	signal WX10422: std_logic; attribute dont_touch of WX10422: signal is true;
	signal WX10423: std_logic; attribute dont_touch of WX10423: signal is true;
	signal WX10424: std_logic; attribute dont_touch of WX10424: signal is true;
	signal WX10425: std_logic; attribute dont_touch of WX10425: signal is true;
	signal WX10426: std_logic; attribute dont_touch of WX10426: signal is true;
	signal WX10427: std_logic; attribute dont_touch of WX10427: signal is true;
	signal WX10428: std_logic; attribute dont_touch of WX10428: signal is true;
	signal WX10429: std_logic; attribute dont_touch of WX10429: signal is true;
	signal WX10430: std_logic; attribute dont_touch of WX10430: signal is true;
	signal WX10431: std_logic; attribute dont_touch of WX10431: signal is true;
	signal WX10432: std_logic; attribute dont_touch of WX10432: signal is true;
	signal WX10433: std_logic; attribute dont_touch of WX10433: signal is true;
	signal WX10434: std_logic; attribute dont_touch of WX10434: signal is true;
	signal WX10435: std_logic; attribute dont_touch of WX10435: signal is true;
	signal WX10436: std_logic; attribute dont_touch of WX10436: signal is true;
	signal WX10437: std_logic; attribute dont_touch of WX10437: signal is true;
	signal WX10438: std_logic; attribute dont_touch of WX10438: signal is true;
	signal WX10439: std_logic; attribute dont_touch of WX10439: signal is true;
	signal WX10440: std_logic; attribute dont_touch of WX10440: signal is true;
	signal WX10441: std_logic; attribute dont_touch of WX10441: signal is true;
	signal WX10442: std_logic; attribute dont_touch of WX10442: signal is true;
	signal WX10443: std_logic; attribute dont_touch of WX10443: signal is true;
	signal WX10444: std_logic; attribute dont_touch of WX10444: signal is true;
	signal WX10445: std_logic; attribute dont_touch of WX10445: signal is true;
	signal WX10446: std_logic; attribute dont_touch of WX10446: signal is true;
	signal WX10447: std_logic; attribute dont_touch of WX10447: signal is true;
	signal WX10448: std_logic; attribute dont_touch of WX10448: signal is true;
	signal WX10449: std_logic; attribute dont_touch of WX10449: signal is true;
	signal WX10450: std_logic; attribute dont_touch of WX10450: signal is true;
	signal WX10451: std_logic; attribute dont_touch of WX10451: signal is true;
	signal WX10452: std_logic; attribute dont_touch of WX10452: signal is true;
	signal WX10453: std_logic; attribute dont_touch of WX10453: signal is true;
	signal WX10454: std_logic; attribute dont_touch of WX10454: signal is true;
	signal WX10455: std_logic; attribute dont_touch of WX10455: signal is true;
	signal WX10456: std_logic; attribute dont_touch of WX10456: signal is true;
	signal WX10457: std_logic; attribute dont_touch of WX10457: signal is true;
	signal WX10458: std_logic; attribute dont_touch of WX10458: signal is true;
	signal WX10459: std_logic; attribute dont_touch of WX10459: signal is true;
	signal WX10460: std_logic; attribute dont_touch of WX10460: signal is true;
	signal WX10461: std_logic; attribute dont_touch of WX10461: signal is true;
	signal WX10462: std_logic; attribute dont_touch of WX10462: signal is true;
	signal WX10463: std_logic; attribute dont_touch of WX10463: signal is true;
	signal WX10464: std_logic; attribute dont_touch of WX10464: signal is true;
	signal WX10465: std_logic; attribute dont_touch of WX10465: signal is true;
	signal WX10466: std_logic; attribute dont_touch of WX10466: signal is true;
	signal WX10467: std_logic; attribute dont_touch of WX10467: signal is true;
	signal WX10468: std_logic; attribute dont_touch of WX10468: signal is true;
	signal WX10469: std_logic; attribute dont_touch of WX10469: signal is true;
	signal WX10470: std_logic; attribute dont_touch of WX10470: signal is true;
	signal WX10471: std_logic; attribute dont_touch of WX10471: signal is true;
	signal WX10472: std_logic; attribute dont_touch of WX10472: signal is true;
	signal WX10473: std_logic; attribute dont_touch of WX10473: signal is true;
	signal WX10474: std_logic; attribute dont_touch of WX10474: signal is true;
	signal WX10475: std_logic; attribute dont_touch of WX10475: signal is true;
	signal WX10476: std_logic; attribute dont_touch of WX10476: signal is true;
	signal WX10477: std_logic; attribute dont_touch of WX10477: signal is true;
	signal WX10478: std_logic; attribute dont_touch of WX10478: signal is true;
	signal WX10479: std_logic; attribute dont_touch of WX10479: signal is true;
	signal WX10480: std_logic; attribute dont_touch of WX10480: signal is true;
	signal WX10481: std_logic; attribute dont_touch of WX10481: signal is true;
	signal WX10482: std_logic; attribute dont_touch of WX10482: signal is true;
	signal WX10483: std_logic; attribute dont_touch of WX10483: signal is true;
	signal WX10484: std_logic; attribute dont_touch of WX10484: signal is true;
	signal WX10485: std_logic; attribute dont_touch of WX10485: signal is true;
	signal WX10486: std_logic; attribute dont_touch of WX10486: signal is true;
	signal WX10487: std_logic; attribute dont_touch of WX10487: signal is true;
	signal WX10488: std_logic; attribute dont_touch of WX10488: signal is true;
	signal WX10489: std_logic; attribute dont_touch of WX10489: signal is true;
	signal WX10490: std_logic; attribute dont_touch of WX10490: signal is true;
	signal WX10491: std_logic; attribute dont_touch of WX10491: signal is true;
	signal WX10492: std_logic; attribute dont_touch of WX10492: signal is true;
	signal WX10493: std_logic; attribute dont_touch of WX10493: signal is true;
	signal WX10494: std_logic; attribute dont_touch of WX10494: signal is true;
	signal WX10495: std_logic; attribute dont_touch of WX10495: signal is true;
	signal WX10496: std_logic; attribute dont_touch of WX10496: signal is true;
	signal WX10497: std_logic; attribute dont_touch of WX10497: signal is true;
	signal WX10498: std_logic; attribute dont_touch of WX10498: signal is true;
	signal WX10499: std_logic; attribute dont_touch of WX10499: signal is true;
	signal WX10500: std_logic; attribute dont_touch of WX10500: signal is true;
	signal WX10501: std_logic; attribute dont_touch of WX10501: signal is true;
	signal WX10502: std_logic; attribute dont_touch of WX10502: signal is true;
	signal WX10503: std_logic; attribute dont_touch of WX10503: signal is true;
	signal WX10504: std_logic; attribute dont_touch of WX10504: signal is true;
	signal WX10505: std_logic; attribute dont_touch of WX10505: signal is true;
	signal WX10506: std_logic; attribute dont_touch of WX10506: signal is true;
	signal WX10507: std_logic; attribute dont_touch of WX10507: signal is true;
	signal WX10508: std_logic; attribute dont_touch of WX10508: signal is true;
	signal WX10509: std_logic; attribute dont_touch of WX10509: signal is true;
	signal WX10510: std_logic; attribute dont_touch of WX10510: signal is true;
	signal WX10511: std_logic; attribute dont_touch of WX10511: signal is true;
	signal WX10512: std_logic; attribute dont_touch of WX10512: signal is true;
	signal WX10513: std_logic; attribute dont_touch of WX10513: signal is true;
	signal WX10514: std_logic; attribute dont_touch of WX10514: signal is true;
	signal WX10515: std_logic; attribute dont_touch of WX10515: signal is true;
	signal WX10516: std_logic; attribute dont_touch of WX10516: signal is true;
	signal WX10517: std_logic; attribute dont_touch of WX10517: signal is true;
	signal WX10518: std_logic; attribute dont_touch of WX10518: signal is true;
	signal WX10519: std_logic; attribute dont_touch of WX10519: signal is true;
	signal WX10520: std_logic; attribute dont_touch of WX10520: signal is true;
	signal WX10521: std_logic; attribute dont_touch of WX10521: signal is true;
	signal WX10522: std_logic; attribute dont_touch of WX10522: signal is true;
	signal WX10523: std_logic; attribute dont_touch of WX10523: signal is true;
	signal WX10524: std_logic; attribute dont_touch of WX10524: signal is true;
	signal WX10525: std_logic; attribute dont_touch of WX10525: signal is true;
	signal WX10526: std_logic; attribute dont_touch of WX10526: signal is true;
	signal WX10527: std_logic; attribute dont_touch of WX10527: signal is true;
	signal WX10528: std_logic; attribute dont_touch of WX10528: signal is true;
	signal WX10529: std_logic; attribute dont_touch of WX10529: signal is true;
	signal WX10530: std_logic; attribute dont_touch of WX10530: signal is true;
	signal WX10531: std_logic; attribute dont_touch of WX10531: signal is true;
	signal WX10532: std_logic; attribute dont_touch of WX10532: signal is true;
	signal WX10533: std_logic; attribute dont_touch of WX10533: signal is true;
	signal WX10534: std_logic; attribute dont_touch of WX10534: signal is true;
	signal WX10535: std_logic; attribute dont_touch of WX10535: signal is true;
	signal WX10536: std_logic; attribute dont_touch of WX10536: signal is true;
	signal WX10537: std_logic; attribute dont_touch of WX10537: signal is true;
	signal WX10538: std_logic; attribute dont_touch of WX10538: signal is true;
	signal WX10539: std_logic; attribute dont_touch of WX10539: signal is true;
	signal WX10540: std_logic; attribute dont_touch of WX10540: signal is true;
	signal WX10541: std_logic; attribute dont_touch of WX10541: signal is true;
	signal WX10542: std_logic; attribute dont_touch of WX10542: signal is true;
	signal WX10543: std_logic; attribute dont_touch of WX10543: signal is true;
	signal WX10544: std_logic; attribute dont_touch of WX10544: signal is true;
	signal WX10545: std_logic; attribute dont_touch of WX10545: signal is true;
	signal WX10546: std_logic; attribute dont_touch of WX10546: signal is true;
	signal WX10547: std_logic; attribute dont_touch of WX10547: signal is true;
	signal WX10548: std_logic; attribute dont_touch of WX10548: signal is true;
	signal WX10549: std_logic; attribute dont_touch of WX10549: signal is true;
	signal WX10550: std_logic; attribute dont_touch of WX10550: signal is true;
	signal WX10551: std_logic; attribute dont_touch of WX10551: signal is true;
	signal WX10552: std_logic; attribute dont_touch of WX10552: signal is true;
	signal WX10553: std_logic; attribute dont_touch of WX10553: signal is true;
	signal WX10554: std_logic; attribute dont_touch of WX10554: signal is true;
	signal WX10555: std_logic; attribute dont_touch of WX10555: signal is true;
	signal WX10556: std_logic; attribute dont_touch of WX10556: signal is true;
	signal WX10557: std_logic; attribute dont_touch of WX10557: signal is true;
	signal WX10558: std_logic; attribute dont_touch of WX10558: signal is true;
	signal WX10559: std_logic; attribute dont_touch of WX10559: signal is true;
	signal WX10560: std_logic; attribute dont_touch of WX10560: signal is true;
	signal WX10561: std_logic; attribute dont_touch of WX10561: signal is true;
	signal WX10562: std_logic; attribute dont_touch of WX10562: signal is true;
	signal WX10563: std_logic; attribute dont_touch of WX10563: signal is true;
	signal WX10564: std_logic; attribute dont_touch of WX10564: signal is true;
	signal WX10565: std_logic; attribute dont_touch of WX10565: signal is true;
	signal WX10566: std_logic; attribute dont_touch of WX10566: signal is true;
	signal WX10567: std_logic; attribute dont_touch of WX10567: signal is true;
	signal WX10568: std_logic; attribute dont_touch of WX10568: signal is true;
	signal WX10569: std_logic; attribute dont_touch of WX10569: signal is true;
	signal WX10570: std_logic; attribute dont_touch of WX10570: signal is true;
	signal WX10571: std_logic; attribute dont_touch of WX10571: signal is true;
	signal WX10572: std_logic; attribute dont_touch of WX10572: signal is true;
	signal WX10573: std_logic; attribute dont_touch of WX10573: signal is true;
	signal WX10574: std_logic; attribute dont_touch of WX10574: signal is true;
	signal WX10575: std_logic; attribute dont_touch of WX10575: signal is true;
	signal WX10576: std_logic; attribute dont_touch of WX10576: signal is true;
	signal WX10577: std_logic; attribute dont_touch of WX10577: signal is true;
	signal WX10578: std_logic; attribute dont_touch of WX10578: signal is true;
	signal WX10579: std_logic; attribute dont_touch of WX10579: signal is true;
	signal WX10580: std_logic; attribute dont_touch of WX10580: signal is true;
	signal WX10581: std_logic; attribute dont_touch of WX10581: signal is true;
	signal WX10582: std_logic; attribute dont_touch of WX10582: signal is true;
	signal WX10583: std_logic; attribute dont_touch of WX10583: signal is true;
	signal WX10584: std_logic; attribute dont_touch of WX10584: signal is true;
	signal WX10585: std_logic; attribute dont_touch of WX10585: signal is true;
	signal WX10586: std_logic; attribute dont_touch of WX10586: signal is true;
	signal WX10587: std_logic; attribute dont_touch of WX10587: signal is true;
	signal WX10588: std_logic; attribute dont_touch of WX10588: signal is true;
	signal WX10589: std_logic; attribute dont_touch of WX10589: signal is true;
	signal WX10590: std_logic; attribute dont_touch of WX10590: signal is true;
	signal WX10591: std_logic; attribute dont_touch of WX10591: signal is true;
	signal WX10592: std_logic; attribute dont_touch of WX10592: signal is true;
	signal WX10593: std_logic; attribute dont_touch of WX10593: signal is true;
	signal WX10594: std_logic; attribute dont_touch of WX10594: signal is true;
	signal WX10595: std_logic; attribute dont_touch of WX10595: signal is true;
	signal WX10596: std_logic; attribute dont_touch of WX10596: signal is true;
	signal WX10597: std_logic; attribute dont_touch of WX10597: signal is true;
	signal WX10598: std_logic; attribute dont_touch of WX10598: signal is true;
	signal WX10599: std_logic; attribute dont_touch of WX10599: signal is true;
	signal WX10600: std_logic; attribute dont_touch of WX10600: signal is true;
	signal WX10601: std_logic; attribute dont_touch of WX10601: signal is true;
	signal WX10602: std_logic; attribute dont_touch of WX10602: signal is true;
	signal WX10603: std_logic; attribute dont_touch of WX10603: signal is true;
	signal WX10604: std_logic; attribute dont_touch of WX10604: signal is true;
	signal WX10605: std_logic; attribute dont_touch of WX10605: signal is true;
	signal WX10606: std_logic; attribute dont_touch of WX10606: signal is true;
	signal WX10607: std_logic; attribute dont_touch of WX10607: signal is true;
	signal WX10608: std_logic; attribute dont_touch of WX10608: signal is true;
	signal WX10609: std_logic; attribute dont_touch of WX10609: signal is true;
	signal WX10610: std_logic; attribute dont_touch of WX10610: signal is true;
	signal WX10611: std_logic; attribute dont_touch of WX10611: signal is true;
	signal WX10612: std_logic; attribute dont_touch of WX10612: signal is true;
	signal WX10613: std_logic; attribute dont_touch of WX10613: signal is true;
	signal WX10614: std_logic; attribute dont_touch of WX10614: signal is true;
	signal WX10615: std_logic; attribute dont_touch of WX10615: signal is true;
	signal WX10616: std_logic; attribute dont_touch of WX10616: signal is true;
	signal WX10617: std_logic; attribute dont_touch of WX10617: signal is true;
	signal WX10618: std_logic; attribute dont_touch of WX10618: signal is true;
	signal WX10619: std_logic; attribute dont_touch of WX10619: signal is true;
	signal WX10620: std_logic; attribute dont_touch of WX10620: signal is true;
	signal WX10621: std_logic; attribute dont_touch of WX10621: signal is true;
	signal WX10622: std_logic; attribute dont_touch of WX10622: signal is true;
	signal WX10623: std_logic; attribute dont_touch of WX10623: signal is true;
	signal WX10624: std_logic; attribute dont_touch of WX10624: signal is true;
	signal WX10625: std_logic; attribute dont_touch of WX10625: signal is true;
	signal WX10626: std_logic; attribute dont_touch of WX10626: signal is true;
	signal WX10627: std_logic; attribute dont_touch of WX10627: signal is true;
	signal WX10628: std_logic; attribute dont_touch of WX10628: signal is true;
	signal WX10629: std_logic; attribute dont_touch of WX10629: signal is true;
	signal WX10630: std_logic; attribute dont_touch of WX10630: signal is true;
	signal WX10631: std_logic; attribute dont_touch of WX10631: signal is true;
	signal WX10632: std_logic; attribute dont_touch of WX10632: signal is true;
	signal WX10633: std_logic; attribute dont_touch of WX10633: signal is true;
	signal WX10634: std_logic; attribute dont_touch of WX10634: signal is true;
	signal WX10635: std_logic; attribute dont_touch of WX10635: signal is true;
	signal WX10636: std_logic; attribute dont_touch of WX10636: signal is true;
	signal WX10637: std_logic; attribute dont_touch of WX10637: signal is true;
	signal WX10638: std_logic; attribute dont_touch of WX10638: signal is true;
	signal WX10639: std_logic; attribute dont_touch of WX10639: signal is true;
	signal WX10640: std_logic; attribute dont_touch of WX10640: signal is true;
	signal WX10641: std_logic; attribute dont_touch of WX10641: signal is true;
	signal WX10642: std_logic; attribute dont_touch of WX10642: signal is true;
	signal WX10643: std_logic; attribute dont_touch of WX10643: signal is true;
	signal WX10644: std_logic; attribute dont_touch of WX10644: signal is true;
	signal WX10645: std_logic; attribute dont_touch of WX10645: signal is true;
	signal WX10646: std_logic; attribute dont_touch of WX10646: signal is true;
	signal WX10647: std_logic; attribute dont_touch of WX10647: signal is true;
	signal WX10648: std_logic; attribute dont_touch of WX10648: signal is true;
	signal WX10649: std_logic; attribute dont_touch of WX10649: signal is true;
	signal WX10650: std_logic; attribute dont_touch of WX10650: signal is true;
	signal WX10651: std_logic; attribute dont_touch of WX10651: signal is true;
	signal WX10652: std_logic; attribute dont_touch of WX10652: signal is true;
	signal WX10653: std_logic; attribute dont_touch of WX10653: signal is true;
	signal WX10654: std_logic; attribute dont_touch of WX10654: signal is true;
	signal WX10655: std_logic; attribute dont_touch of WX10655: signal is true;
	signal WX10656: std_logic; attribute dont_touch of WX10656: signal is true;
	signal WX10657: std_logic; attribute dont_touch of WX10657: signal is true;
	signal WX10658: std_logic; attribute dont_touch of WX10658: signal is true;
	signal WX10659: std_logic; attribute dont_touch of WX10659: signal is true;
	signal WX10660: std_logic; attribute dont_touch of WX10660: signal is true;
	signal WX10661: std_logic; attribute dont_touch of WX10661: signal is true;
	signal WX10662: std_logic; attribute dont_touch of WX10662: signal is true;
	signal WX10663: std_logic; attribute dont_touch of WX10663: signal is true;
	signal WX10664: std_logic; attribute dont_touch of WX10664: signal is true;
	signal WX10665: std_logic; attribute dont_touch of WX10665: signal is true;
	signal WX10666: std_logic; attribute dont_touch of WX10666: signal is true;
	signal WX10667: std_logic; attribute dont_touch of WX10667: signal is true;
	signal WX10668: std_logic; attribute dont_touch of WX10668: signal is true;
	signal WX10669: std_logic; attribute dont_touch of WX10669: signal is true;
	signal WX10670: std_logic; attribute dont_touch of WX10670: signal is true;
	signal WX10671: std_logic; attribute dont_touch of WX10671: signal is true;
	signal WX10672: std_logic; attribute dont_touch of WX10672: signal is true;
	signal WX10673: std_logic; attribute dont_touch of WX10673: signal is true;
	signal WX10674: std_logic; attribute dont_touch of WX10674: signal is true;
	signal WX10675: std_logic; attribute dont_touch of WX10675: signal is true;
	signal WX10676: std_logic; attribute dont_touch of WX10676: signal is true;
	signal WX10677: std_logic; attribute dont_touch of WX10677: signal is true;
	signal WX10678: std_logic; attribute dont_touch of WX10678: signal is true;
	signal WX10679: std_logic; attribute dont_touch of WX10679: signal is true;
	signal WX10680: std_logic; attribute dont_touch of WX10680: signal is true;
	signal WX10681: std_logic; attribute dont_touch of WX10681: signal is true;
	signal WX10682: std_logic; attribute dont_touch of WX10682: signal is true;
	signal WX10683: std_logic; attribute dont_touch of WX10683: signal is true;
	signal WX10684: std_logic; attribute dont_touch of WX10684: signal is true;
	signal WX10685: std_logic; attribute dont_touch of WX10685: signal is true;
	signal WX10686: std_logic; attribute dont_touch of WX10686: signal is true;
	signal WX10687: std_logic; attribute dont_touch of WX10687: signal is true;
	signal WX10688: std_logic; attribute dont_touch of WX10688: signal is true;
	signal WX10689: std_logic; attribute dont_touch of WX10689: signal is true;
	signal WX10690: std_logic; attribute dont_touch of WX10690: signal is true;
	signal WX10691: std_logic; attribute dont_touch of WX10691: signal is true;
	signal WX10692: std_logic; attribute dont_touch of WX10692: signal is true;
	signal WX10693: std_logic; attribute dont_touch of WX10693: signal is true;
	signal WX10694: std_logic; attribute dont_touch of WX10694: signal is true;
	signal WX10695: std_logic; attribute dont_touch of WX10695: signal is true;
	signal WX10696: std_logic; attribute dont_touch of WX10696: signal is true;
	signal WX10697: std_logic; attribute dont_touch of WX10697: signal is true;
	signal WX10698: std_logic; attribute dont_touch of WX10698: signal is true;
	signal WX10699: std_logic; attribute dont_touch of WX10699: signal is true;
	signal WX10700: std_logic; attribute dont_touch of WX10700: signal is true;
	signal WX10701: std_logic; attribute dont_touch of WX10701: signal is true;
	signal WX10702: std_logic; attribute dont_touch of WX10702: signal is true;
	signal WX10703: std_logic; attribute dont_touch of WX10703: signal is true;
	signal WX10704: std_logic; attribute dont_touch of WX10704: signal is true;
	signal WX10705: std_logic; attribute dont_touch of WX10705: signal is true;
	signal WX10706: std_logic; attribute dont_touch of WX10706: signal is true;
	signal WX10707: std_logic; attribute dont_touch of WX10707: signal is true;
	signal WX10708: std_logic; attribute dont_touch of WX10708: signal is true;
	signal WX10709: std_logic; attribute dont_touch of WX10709: signal is true;
	signal WX10710: std_logic; attribute dont_touch of WX10710: signal is true;
	signal WX10711: std_logic; attribute dont_touch of WX10711: signal is true;
	signal WX10712: std_logic; attribute dont_touch of WX10712: signal is true;
	signal WX10713: std_logic; attribute dont_touch of WX10713: signal is true;
	signal WX10714: std_logic; attribute dont_touch of WX10714: signal is true;
	signal WX10715: std_logic; attribute dont_touch of WX10715: signal is true;
	signal WX10716: std_logic; attribute dont_touch of WX10716: signal is true;
	signal WX10717: std_logic; attribute dont_touch of WX10717: signal is true;
	signal WX10718: std_logic; attribute dont_touch of WX10718: signal is true;
	signal WX10719: std_logic; attribute dont_touch of WX10719: signal is true;
	signal WX10720: std_logic; attribute dont_touch of WX10720: signal is true;
	signal WX10721: std_logic; attribute dont_touch of WX10721: signal is true;
	signal WX10722: std_logic; attribute dont_touch of WX10722: signal is true;
	signal WX10723: std_logic; attribute dont_touch of WX10723: signal is true;
	signal WX10724: std_logic; attribute dont_touch of WX10724: signal is true;
	signal WX10725: std_logic; attribute dont_touch of WX10725: signal is true;
	signal WX10726: std_logic; attribute dont_touch of WX10726: signal is true;
	signal WX10727: std_logic; attribute dont_touch of WX10727: signal is true;
	signal WX10728: std_logic; attribute dont_touch of WX10728: signal is true;
	signal WX10729: std_logic; attribute dont_touch of WX10729: signal is true;
	signal WX10730: std_logic; attribute dont_touch of WX10730: signal is true;
	signal WX10731: std_logic; attribute dont_touch of WX10731: signal is true;
	signal WX10732: std_logic; attribute dont_touch of WX10732: signal is true;
	signal WX10733: std_logic; attribute dont_touch of WX10733: signal is true;
	signal WX10734: std_logic; attribute dont_touch of WX10734: signal is true;
	signal WX10735: std_logic; attribute dont_touch of WX10735: signal is true;
	signal WX10736: std_logic; attribute dont_touch of WX10736: signal is true;
	signal WX10737: std_logic; attribute dont_touch of WX10737: signal is true;
	signal WX10738: std_logic; attribute dont_touch of WX10738: signal is true;
	signal WX10739: std_logic; attribute dont_touch of WX10739: signal is true;
	signal WX10740: std_logic; attribute dont_touch of WX10740: signal is true;
	signal WX10741: std_logic; attribute dont_touch of WX10741: signal is true;
	signal WX10742: std_logic; attribute dont_touch of WX10742: signal is true;
	signal WX10743: std_logic; attribute dont_touch of WX10743: signal is true;
	signal WX10744: std_logic; attribute dont_touch of WX10744: signal is true;
	signal WX10745: std_logic; attribute dont_touch of WX10745: signal is true;
	signal WX10746: std_logic; attribute dont_touch of WX10746: signal is true;
	signal WX10747: std_logic; attribute dont_touch of WX10747: signal is true;
	signal WX10748: std_logic; attribute dont_touch of WX10748: signal is true;
	signal WX10749: std_logic; attribute dont_touch of WX10749: signal is true;
	signal WX10750: std_logic; attribute dont_touch of WX10750: signal is true;
	signal WX10751: std_logic; attribute dont_touch of WX10751: signal is true;
	signal WX10752: std_logic; attribute dont_touch of WX10752: signal is true;
	signal WX10753: std_logic; attribute dont_touch of WX10753: signal is true;
	signal WX10754: std_logic; attribute dont_touch of WX10754: signal is true;
	signal WX10755: std_logic; attribute dont_touch of WX10755: signal is true;
	signal WX10756: std_logic; attribute dont_touch of WX10756: signal is true;
	signal WX10757: std_logic; attribute dont_touch of WX10757: signal is true;
	signal WX10758: std_logic; attribute dont_touch of WX10758: signal is true;
	signal WX10759: std_logic; attribute dont_touch of WX10759: signal is true;
	signal WX10760: std_logic; attribute dont_touch of WX10760: signal is true;
	signal WX10761: std_logic; attribute dont_touch of WX10761: signal is true;
	signal WX10762: std_logic; attribute dont_touch of WX10762: signal is true;
	signal WX10763: std_logic; attribute dont_touch of WX10763: signal is true;
	signal WX10764: std_logic; attribute dont_touch of WX10764: signal is true;
	signal WX10765: std_logic; attribute dont_touch of WX10765: signal is true;
	signal WX10766: std_logic; attribute dont_touch of WX10766: signal is true;
	signal WX10767: std_logic; attribute dont_touch of WX10767: signal is true;
	signal WX10768: std_logic; attribute dont_touch of WX10768: signal is true;
	signal WX10769: std_logic; attribute dont_touch of WX10769: signal is true;
	signal WX10770: std_logic; attribute dont_touch of WX10770: signal is true;
	signal WX10771: std_logic; attribute dont_touch of WX10771: signal is true;
	signal WX10772: std_logic; attribute dont_touch of WX10772: signal is true;
	signal WX10773: std_logic; attribute dont_touch of WX10773: signal is true;
	signal WX10774: std_logic; attribute dont_touch of WX10774: signal is true;
	signal WX10775: std_logic; attribute dont_touch of WX10775: signal is true;
	signal WX10776: std_logic; attribute dont_touch of WX10776: signal is true;
	signal WX10777: std_logic; attribute dont_touch of WX10777: signal is true;
	signal WX10778: std_logic; attribute dont_touch of WX10778: signal is true;
	signal WX10779: std_logic; attribute dont_touch of WX10779: signal is true;
	signal WX10780: std_logic; attribute dont_touch of WX10780: signal is true;
	signal WX10781: std_logic; attribute dont_touch of WX10781: signal is true;
	signal WX10782: std_logic; attribute dont_touch of WX10782: signal is true;
	signal WX10783: std_logic; attribute dont_touch of WX10783: signal is true;
	signal WX10784: std_logic; attribute dont_touch of WX10784: signal is true;
	signal WX10785: std_logic; attribute dont_touch of WX10785: signal is true;
	signal WX10786: std_logic; attribute dont_touch of WX10786: signal is true;
	signal WX10787: std_logic; attribute dont_touch of WX10787: signal is true;
	signal WX10788: std_logic; attribute dont_touch of WX10788: signal is true;
	signal WX10789: std_logic; attribute dont_touch of WX10789: signal is true;
	signal WX10790: std_logic; attribute dont_touch of WX10790: signal is true;
	signal WX10791: std_logic; attribute dont_touch of WX10791: signal is true;
	signal WX10792: std_logic; attribute dont_touch of WX10792: signal is true;
	signal WX10793: std_logic; attribute dont_touch of WX10793: signal is true;
	signal WX10794: std_logic; attribute dont_touch of WX10794: signal is true;
	signal WX10795: std_logic; attribute dont_touch of WX10795: signal is true;
	signal WX10796: std_logic; attribute dont_touch of WX10796: signal is true;
	signal WX10797: std_logic; attribute dont_touch of WX10797: signal is true;
	signal WX10798: std_logic; attribute dont_touch of WX10798: signal is true;
	signal WX10799: std_logic; attribute dont_touch of WX10799: signal is true;
	signal WX10800: std_logic; attribute dont_touch of WX10800: signal is true;
	signal WX10801: std_logic; attribute dont_touch of WX10801: signal is true;
	signal WX10802: std_logic; attribute dont_touch of WX10802: signal is true;
	signal WX10803: std_logic; attribute dont_touch of WX10803: signal is true;
	signal WX10804: std_logic; attribute dont_touch of WX10804: signal is true;
	signal WX10805: std_logic; attribute dont_touch of WX10805: signal is true;
	signal WX10806: std_logic; attribute dont_touch of WX10806: signal is true;
	signal WX10807: std_logic; attribute dont_touch of WX10807: signal is true;
	signal WX10808: std_logic; attribute dont_touch of WX10808: signal is true;
	signal WX10809: std_logic; attribute dont_touch of WX10809: signal is true;
	signal WX10810: std_logic; attribute dont_touch of WX10810: signal is true;
	signal WX10811: std_logic; attribute dont_touch of WX10811: signal is true;
	signal WX10812: std_logic; attribute dont_touch of WX10812: signal is true;
	signal WX10813: std_logic; attribute dont_touch of WX10813: signal is true;
	signal WX10814: std_logic; attribute dont_touch of WX10814: signal is true;
	signal WX10815: std_logic; attribute dont_touch of WX10815: signal is true;
	signal WX10816: std_logic; attribute dont_touch of WX10816: signal is true;
	signal WX10817: std_logic; attribute dont_touch of WX10817: signal is true;
	signal WX10818: std_logic; attribute dont_touch of WX10818: signal is true;
	signal WX10819: std_logic; attribute dont_touch of WX10819: signal is true;
	signal WX10820: std_logic; attribute dont_touch of WX10820: signal is true;
	signal WX10821: std_logic; attribute dont_touch of WX10821: signal is true;
	signal WX10822: std_logic; attribute dont_touch of WX10822: signal is true;
	signal WX10823: std_logic; attribute dont_touch of WX10823: signal is true;
	signal WX10824: std_logic; attribute dont_touch of WX10824: signal is true;
	signal WX10825: std_logic; attribute dont_touch of WX10825: signal is true;
	signal WX10826: std_logic; attribute dont_touch of WX10826: signal is true;
	signal WX10827: std_logic; attribute dont_touch of WX10827: signal is true;
	signal WX10828: std_logic; attribute dont_touch of WX10828: signal is true;
	signal WX10829: std_logic; attribute dont_touch of WX10829: signal is true;
	signal WX10830: std_logic; attribute dont_touch of WX10830: signal is true;
	signal WX10831: std_logic; attribute dont_touch of WX10831: signal is true;
	signal WX10832: std_logic; attribute dont_touch of WX10832: signal is true;
	signal WX10833: std_logic; attribute dont_touch of WX10833: signal is true;
	signal WX10834: std_logic; attribute dont_touch of WX10834: signal is true;
	signal WX10835: std_logic; attribute dont_touch of WX10835: signal is true;
	signal WX10836: std_logic; attribute dont_touch of WX10836: signal is true;
	signal WX10837: std_logic; attribute dont_touch of WX10837: signal is true;
	signal WX10838: std_logic; attribute dont_touch of WX10838: signal is true;
	signal WX10839: std_logic; attribute dont_touch of WX10839: signal is true;
	signal WX10840: std_logic; attribute dont_touch of WX10840: signal is true;
	signal WX10841: std_logic; attribute dont_touch of WX10841: signal is true;
	signal WX10842: std_logic; attribute dont_touch of WX10842: signal is true;
	signal WX10843: std_logic; attribute dont_touch of WX10843: signal is true;
	signal WX10844: std_logic; attribute dont_touch of WX10844: signal is true;
	signal WX10845: std_logic; attribute dont_touch of WX10845: signal is true;
	signal WX10846: std_logic; attribute dont_touch of WX10846: signal is true;
	signal WX10847: std_logic; attribute dont_touch of WX10847: signal is true;
	signal WX10848: std_logic; attribute dont_touch of WX10848: signal is true;
	signal WX10849: std_logic; attribute dont_touch of WX10849: signal is true;
	signal WX10850: std_logic; attribute dont_touch of WX10850: signal is true;
	signal WX10851: std_logic; attribute dont_touch of WX10851: signal is true;
	signal WX10852: std_logic; attribute dont_touch of WX10852: signal is true;
	signal WX10853: std_logic; attribute dont_touch of WX10853: signal is true;
	signal WX10854: std_logic; attribute dont_touch of WX10854: signal is true;
	signal WX10855: std_logic; attribute dont_touch of WX10855: signal is true;
	signal WX10856: std_logic; attribute dont_touch of WX10856: signal is true;
	signal WX10857: std_logic; attribute dont_touch of WX10857: signal is true;
	signal WX10858: std_logic; attribute dont_touch of WX10858: signal is true;
	signal WX10859: std_logic; attribute dont_touch of WX10859: signal is true;
	signal WX10860: std_logic; attribute dont_touch of WX10860: signal is true;
	signal WX10861: std_logic; attribute dont_touch of WX10861: signal is true;
	signal WX10862: std_logic; attribute dont_touch of WX10862: signal is true;
	signal WX10863: std_logic; attribute dont_touch of WX10863: signal is true;
	signal WX10864: std_logic; attribute dont_touch of WX10864: signal is true;
	signal WX10865: std_logic; attribute dont_touch of WX10865: signal is true;
	signal WX10866: std_logic; attribute dont_touch of WX10866: signal is true;
	signal WX10867: std_logic; attribute dont_touch of WX10867: signal is true;
	signal WX10868: std_logic; attribute dont_touch of WX10868: signal is true;
	signal WX10869: std_logic; attribute dont_touch of WX10869: signal is true;
	signal WX10870: std_logic; attribute dont_touch of WX10870: signal is true;
	signal WX10871: std_logic; attribute dont_touch of WX10871: signal is true;
	signal WX10872: std_logic; attribute dont_touch of WX10872: signal is true;
	signal WX10873: std_logic; attribute dont_touch of WX10873: signal is true;
	signal WX10874: std_logic; attribute dont_touch of WX10874: signal is true;
	signal WX10875: std_logic; attribute dont_touch of WX10875: signal is true;
	signal WX10876: std_logic; attribute dont_touch of WX10876: signal is true;
	signal WX10877: std_logic; attribute dont_touch of WX10877: signal is true;
	signal WX10878: std_logic; attribute dont_touch of WX10878: signal is true;
	signal WX10879: std_logic; attribute dont_touch of WX10879: signal is true;
	signal WX10880: std_logic; attribute dont_touch of WX10880: signal is true;
	signal WX10881: std_logic; attribute dont_touch of WX10881: signal is true;
	signal WX10882: std_logic; attribute dont_touch of WX10882: signal is true;
	signal WX10883: std_logic; attribute dont_touch of WX10883: signal is true;
	signal WX10884: std_logic; attribute dont_touch of WX10884: signal is true;
	signal WX10885: std_logic; attribute dont_touch of WX10885: signal is true;
	signal WX10886: std_logic; attribute dont_touch of WX10886: signal is true;
	signal WX10887: std_logic; attribute dont_touch of WX10887: signal is true;
	signal WX10888: std_logic; attribute dont_touch of WX10888: signal is true;
	signal WX10889: std_logic; attribute dont_touch of WX10889: signal is true;
	signal WX10890: std_logic; attribute dont_touch of WX10890: signal is true;
	signal WX10891: std_logic; attribute dont_touch of WX10891: signal is true;
	signal WX10892: std_logic; attribute dont_touch of WX10892: signal is true;
	signal WX10893: std_logic; attribute dont_touch of WX10893: signal is true;
	signal WX10894: std_logic; attribute dont_touch of WX10894: signal is true;
	signal WX10895: std_logic; attribute dont_touch of WX10895: signal is true;
	signal WX10896: std_logic; attribute dont_touch of WX10896: signal is true;
	signal WX10897: std_logic; attribute dont_touch of WX10897: signal is true;
	signal WX10898: std_logic; attribute dont_touch of WX10898: signal is true;
	signal WX10899: std_logic; attribute dont_touch of WX10899: signal is true;
	signal WX10900: std_logic; attribute dont_touch of WX10900: signal is true;
	signal WX10901: std_logic; attribute dont_touch of WX10901: signal is true;
	signal WX10902: std_logic; attribute dont_touch of WX10902: signal is true;
	signal WX10903: std_logic; attribute dont_touch of WX10903: signal is true;
	signal WX10904: std_logic; attribute dont_touch of WX10904: signal is true;
	signal WX10905: std_logic; attribute dont_touch of WX10905: signal is true;
	signal WX10906: std_logic; attribute dont_touch of WX10906: signal is true;
	signal WX10907: std_logic; attribute dont_touch of WX10907: signal is true;
	signal WX10908: std_logic; attribute dont_touch of WX10908: signal is true;
	signal WX10909: std_logic; attribute dont_touch of WX10909: signal is true;
	signal WX10910: std_logic; attribute dont_touch of WX10910: signal is true;
	signal WX10911: std_logic; attribute dont_touch of WX10911: signal is true;
	signal WX10912: std_logic; attribute dont_touch of WX10912: signal is true;
	signal WX10913: std_logic; attribute dont_touch of WX10913: signal is true;
	signal WX10914: std_logic; attribute dont_touch of WX10914: signal is true;
	signal WX10915: std_logic; attribute dont_touch of WX10915: signal is true;
	signal WX10916: std_logic; attribute dont_touch of WX10916: signal is true;
	signal WX10917: std_logic; attribute dont_touch of WX10917: signal is true;
	signal WX10918: std_logic; attribute dont_touch of WX10918: signal is true;
	signal WX10919: std_logic; attribute dont_touch of WX10919: signal is true;
	signal WX10920: std_logic; attribute dont_touch of WX10920: signal is true;
	signal WX10921: std_logic; attribute dont_touch of WX10921: signal is true;
	signal WX10922: std_logic; attribute dont_touch of WX10922: signal is true;
	signal WX10923: std_logic; attribute dont_touch of WX10923: signal is true;
	signal WX10924: std_logic; attribute dont_touch of WX10924: signal is true;
	signal WX10925: std_logic; attribute dont_touch of WX10925: signal is true;
	signal WX10926: std_logic; attribute dont_touch of WX10926: signal is true;
	signal WX10927: std_logic; attribute dont_touch of WX10927: signal is true;
	signal WX10928: std_logic; attribute dont_touch of WX10928: signal is true;
	signal WX10929: std_logic; attribute dont_touch of WX10929: signal is true;
	signal WX10930: std_logic; attribute dont_touch of WX10930: signal is true;
	signal WX10931: std_logic; attribute dont_touch of WX10931: signal is true;
	signal WX10932: std_logic; attribute dont_touch of WX10932: signal is true;
	signal WX10933: std_logic; attribute dont_touch of WX10933: signal is true;
	signal WX10934: std_logic; attribute dont_touch of WX10934: signal is true;
	signal WX10935: std_logic; attribute dont_touch of WX10935: signal is true;
	signal WX10936: std_logic; attribute dont_touch of WX10936: signal is true;
	signal WX10937: std_logic; attribute dont_touch of WX10937: signal is true;
	signal WX10938: std_logic; attribute dont_touch of WX10938: signal is true;
	signal WX10939: std_logic; attribute dont_touch of WX10939: signal is true;
	signal WX10940: std_logic; attribute dont_touch of WX10940: signal is true;
	signal WX10941: std_logic; attribute dont_touch of WX10941: signal is true;
	signal WX10942: std_logic; attribute dont_touch of WX10942: signal is true;
	signal WX10943: std_logic; attribute dont_touch of WX10943: signal is true;
	signal WX10944: std_logic; attribute dont_touch of WX10944: signal is true;
	signal WX10945: std_logic; attribute dont_touch of WX10945: signal is true;
	signal WX10946: std_logic; attribute dont_touch of WX10946: signal is true;
	signal WX10947: std_logic; attribute dont_touch of WX10947: signal is true;
	signal WX10948: std_logic; attribute dont_touch of WX10948: signal is true;
	signal WX10949: std_logic; attribute dont_touch of WX10949: signal is true;
	signal WX10950: std_logic; attribute dont_touch of WX10950: signal is true;
	signal WX10951: std_logic; attribute dont_touch of WX10951: signal is true;
	signal WX10952: std_logic; attribute dont_touch of WX10952: signal is true;
	signal WX10953: std_logic; attribute dont_touch of WX10953: signal is true;
	signal WX10954: std_logic; attribute dont_touch of WX10954: signal is true;
	signal WX10955: std_logic; attribute dont_touch of WX10955: signal is true;
	signal WX10956: std_logic; attribute dont_touch of WX10956: signal is true;
	signal WX10957: std_logic; attribute dont_touch of WX10957: signal is true;
	signal WX10958: std_logic; attribute dont_touch of WX10958: signal is true;
	signal WX10959: std_logic; attribute dont_touch of WX10959: signal is true;
	signal WX10960: std_logic; attribute dont_touch of WX10960: signal is true;
	signal WX10961: std_logic; attribute dont_touch of WX10961: signal is true;
	signal WX10962: std_logic; attribute dont_touch of WX10962: signal is true;
	signal WX10963: std_logic; attribute dont_touch of WX10963: signal is true;
	signal WX10964: std_logic; attribute dont_touch of WX10964: signal is true;
	signal WX10965: std_logic; attribute dont_touch of WX10965: signal is true;
	signal WX10966: std_logic; attribute dont_touch of WX10966: signal is true;
	signal WX10967: std_logic; attribute dont_touch of WX10967: signal is true;
	signal WX10968: std_logic; attribute dont_touch of WX10968: signal is true;
	signal WX10969: std_logic; attribute dont_touch of WX10969: signal is true;
	signal WX10970: std_logic; attribute dont_touch of WX10970: signal is true;
	signal WX10971: std_logic; attribute dont_touch of WX10971: signal is true;
	signal WX10972: std_logic; attribute dont_touch of WX10972: signal is true;
	signal WX10973: std_logic; attribute dont_touch of WX10973: signal is true;
	signal WX10974: std_logic; attribute dont_touch of WX10974: signal is true;
	signal WX10975: std_logic; attribute dont_touch of WX10975: signal is true;
	signal WX10976: std_logic; attribute dont_touch of WX10976: signal is true;
	signal WX10977: std_logic; attribute dont_touch of WX10977: signal is true;
	signal WX10978: std_logic; attribute dont_touch of WX10978: signal is true;
	signal WX10979: std_logic; attribute dont_touch of WX10979: signal is true;
	signal WX10980: std_logic; attribute dont_touch of WX10980: signal is true;
	signal WX10981: std_logic; attribute dont_touch of WX10981: signal is true;
	signal WX10982: std_logic; attribute dont_touch of WX10982: signal is true;
	signal WX10983: std_logic; attribute dont_touch of WX10983: signal is true;
	signal WX10984: std_logic; attribute dont_touch of WX10984: signal is true;
	signal WX10985: std_logic; attribute dont_touch of WX10985: signal is true;
	signal WX10986: std_logic; attribute dont_touch of WX10986: signal is true;
	signal WX10987: std_logic; attribute dont_touch of WX10987: signal is true;
	signal WX10988: std_logic; attribute dont_touch of WX10988: signal is true;
	signal WX10989: std_logic; attribute dont_touch of WX10989: signal is true;
	signal WX10990: std_logic; attribute dont_touch of WX10990: signal is true;
	signal WX10991: std_logic; attribute dont_touch of WX10991: signal is true;
	signal WX10992: std_logic; attribute dont_touch of WX10992: signal is true;
	signal WX10993: std_logic; attribute dont_touch of WX10993: signal is true;
	signal WX10994: std_logic; attribute dont_touch of WX10994: signal is true;
	signal WX10995: std_logic; attribute dont_touch of WX10995: signal is true;
	signal WX10996: std_logic; attribute dont_touch of WX10996: signal is true;
	signal WX10997: std_logic; attribute dont_touch of WX10997: signal is true;
	signal WX10998: std_logic; attribute dont_touch of WX10998: signal is true;
	signal WX10999: std_logic; attribute dont_touch of WX10999: signal is true;
	signal WX11000: std_logic; attribute dont_touch of WX11000: signal is true;
	signal WX11001: std_logic; attribute dont_touch of WX11001: signal is true;
	signal WX11002: std_logic; attribute dont_touch of WX11002: signal is true;
	signal WX11003: std_logic; attribute dont_touch of WX11003: signal is true;
	signal WX11004: std_logic; attribute dont_touch of WX11004: signal is true;
	signal WX11005: std_logic; attribute dont_touch of WX11005: signal is true;
	signal WX11006: std_logic; attribute dont_touch of WX11006: signal is true;
	signal WX11007: std_logic; attribute dont_touch of WX11007: signal is true;
	signal WX11008: std_logic; attribute dont_touch of WX11008: signal is true;
	signal WX11009: std_logic; attribute dont_touch of WX11009: signal is true;
	signal WX11010: std_logic; attribute dont_touch of WX11010: signal is true;
	signal WX11011: std_logic; attribute dont_touch of WX11011: signal is true;
	signal WX11012: std_logic; attribute dont_touch of WX11012: signal is true;
	signal WX11013: std_logic; attribute dont_touch of WX11013: signal is true;
	signal WX11014: std_logic; attribute dont_touch of WX11014: signal is true;
	signal WX11015: std_logic; attribute dont_touch of WX11015: signal is true;
	signal WX11016: std_logic; attribute dont_touch of WX11016: signal is true;
	signal WX11017: std_logic; attribute dont_touch of WX11017: signal is true;
	signal WX11018: std_logic; attribute dont_touch of WX11018: signal is true;
	signal WX11019: std_logic; attribute dont_touch of WX11019: signal is true;
	signal WX11020: std_logic; attribute dont_touch of WX11020: signal is true;
	signal WX11021: std_logic; attribute dont_touch of WX11021: signal is true;
	signal WX11022: std_logic; attribute dont_touch of WX11022: signal is true;
	signal WX11023: std_logic; attribute dont_touch of WX11023: signal is true;
	signal WX11024: std_logic; attribute dont_touch of WX11024: signal is true;
	signal WX11025: std_logic; attribute dont_touch of WX11025: signal is true;
	signal WX11026: std_logic; attribute dont_touch of WX11026: signal is true;
	signal WX11027: std_logic; attribute dont_touch of WX11027: signal is true;
	signal WX11028: std_logic; attribute dont_touch of WX11028: signal is true;
	signal WX11029: std_logic; attribute dont_touch of WX11029: signal is true;
	signal WX11030: std_logic; attribute dont_touch of WX11030: signal is true;
	signal WX11031: std_logic; attribute dont_touch of WX11031: signal is true;
	signal WX11032: std_logic; attribute dont_touch of WX11032: signal is true;
	signal WX11033: std_logic; attribute dont_touch of WX11033: signal is true;
	signal WX11034: std_logic; attribute dont_touch of WX11034: signal is true;
	signal WX11035: std_logic; attribute dont_touch of WX11035: signal is true;
	signal WX11036: std_logic; attribute dont_touch of WX11036: signal is true;
	signal WX11037: std_logic; attribute dont_touch of WX11037: signal is true;
	signal WX11038: std_logic; attribute dont_touch of WX11038: signal is true;
	signal WX11039: std_logic; attribute dont_touch of WX11039: signal is true;
	signal WX11040: std_logic; attribute dont_touch of WX11040: signal is true;
	signal WX11041: std_logic; attribute dont_touch of WX11041: signal is true;
	signal WX11042: std_logic; attribute dont_touch of WX11042: signal is true;
	signal WX11043: std_logic; attribute dont_touch of WX11043: signal is true;
	signal WX11044: std_logic; attribute dont_touch of WX11044: signal is true;
	signal WX11045: std_logic; attribute dont_touch of WX11045: signal is true;
	signal WX11046: std_logic; attribute dont_touch of WX11046: signal is true;
	signal WX11047: std_logic; attribute dont_touch of WX11047: signal is true;
	signal WX11048: std_logic; attribute dont_touch of WX11048: signal is true;
	signal WX11049: std_logic; attribute dont_touch of WX11049: signal is true;
	signal WX11050: std_logic; attribute dont_touch of WX11050: signal is true;
	signal WX11051: std_logic; attribute dont_touch of WX11051: signal is true;
	signal WX11052: std_logic; attribute dont_touch of WX11052: signal is true;
	signal WX11053: std_logic; attribute dont_touch of WX11053: signal is true;
	signal WX11054: std_logic; attribute dont_touch of WX11054: signal is true;
	signal WX11055: std_logic; attribute dont_touch of WX11055: signal is true;
	signal WX11056: std_logic; attribute dont_touch of WX11056: signal is true;
	signal WX11057: std_logic; attribute dont_touch of WX11057: signal is true;
	signal WX11058: std_logic; attribute dont_touch of WX11058: signal is true;
	signal WX11059: std_logic; attribute dont_touch of WX11059: signal is true;
	signal WX11060: std_logic; attribute dont_touch of WX11060: signal is true;
	signal WX11061: std_logic; attribute dont_touch of WX11061: signal is true;
	signal WX11062: std_logic; attribute dont_touch of WX11062: signal is true;
	signal WX11063: std_logic; attribute dont_touch of WX11063: signal is true;
	signal WX11064: std_logic; attribute dont_touch of WX11064: signal is true;
	signal WX11065: std_logic; attribute dont_touch of WX11065: signal is true;
	signal WX11066: std_logic; attribute dont_touch of WX11066: signal is true;
	signal WX11067: std_logic; attribute dont_touch of WX11067: signal is true;
	signal WX11068: std_logic; attribute dont_touch of WX11068: signal is true;
	signal WX11069: std_logic; attribute dont_touch of WX11069: signal is true;
	signal WX11070: std_logic; attribute dont_touch of WX11070: signal is true;
	signal WX11071: std_logic; attribute dont_touch of WX11071: signal is true;
	signal WX11072: std_logic; attribute dont_touch of WX11072: signal is true;
	signal WX11073: std_logic; attribute dont_touch of WX11073: signal is true;
	signal WX11074: std_logic; attribute dont_touch of WX11074: signal is true;
	signal WX11075: std_logic; attribute dont_touch of WX11075: signal is true;
	signal WX11076: std_logic; attribute dont_touch of WX11076: signal is true;
	signal WX11077: std_logic; attribute dont_touch of WX11077: signal is true;
	signal WX11078: std_logic; attribute dont_touch of WX11078: signal is true;
	signal WX11079: std_logic; attribute dont_touch of WX11079: signal is true;
	signal WX11080: std_logic; attribute dont_touch of WX11080: signal is true;
	signal WX11081: std_logic; attribute dont_touch of WX11081: signal is true;
	signal WX11082: std_logic; attribute dont_touch of WX11082: signal is true;
	signal WX11083: std_logic; attribute dont_touch of WX11083: signal is true;
	signal WX11084: std_logic; attribute dont_touch of WX11084: signal is true;
	signal WX11085: std_logic; attribute dont_touch of WX11085: signal is true;
	signal WX11086: std_logic; attribute dont_touch of WX11086: signal is true;
	signal WX11087: std_logic; attribute dont_touch of WX11087: signal is true;
	signal WX11088: std_logic; attribute dont_touch of WX11088: signal is true;
	signal WX11089: std_logic; attribute dont_touch of WX11089: signal is true;
	signal WX11090: std_logic; attribute dont_touch of WX11090: signal is true;
	signal WX11091: std_logic; attribute dont_touch of WX11091: signal is true;
	signal WX11092: std_logic; attribute dont_touch of WX11092: signal is true;
	signal WX11093: std_logic; attribute dont_touch of WX11093: signal is true;
	signal WX11094: std_logic; attribute dont_touch of WX11094: signal is true;
	signal WX11095: std_logic; attribute dont_touch of WX11095: signal is true;
	signal WX11096: std_logic; attribute dont_touch of WX11096: signal is true;
	signal WX11097: std_logic; attribute dont_touch of WX11097: signal is true;
	signal WX11098: std_logic; attribute dont_touch of WX11098: signal is true;
	signal WX11099: std_logic; attribute dont_touch of WX11099: signal is true;
	signal WX11100: std_logic; attribute dont_touch of WX11100: signal is true;
	signal WX11101: std_logic; attribute dont_touch of WX11101: signal is true;
	signal WX11102: std_logic; attribute dont_touch of WX11102: signal is true;
	signal WX11103: std_logic; attribute dont_touch of WX11103: signal is true;
	signal WX11104: std_logic; attribute dont_touch of WX11104: signal is true;
	signal WX11105: std_logic; attribute dont_touch of WX11105: signal is true;
	signal WX11106: std_logic; attribute dont_touch of WX11106: signal is true;
	signal WX11107: std_logic; attribute dont_touch of WX11107: signal is true;
	signal WX11108: std_logic; attribute dont_touch of WX11108: signal is true;
	signal WX11109: std_logic; attribute dont_touch of WX11109: signal is true;
	signal WX11110: std_logic; attribute dont_touch of WX11110: signal is true;
	signal WX11111: std_logic; attribute dont_touch of WX11111: signal is true;
	signal WX11112: std_logic; attribute dont_touch of WX11112: signal is true;
	signal WX11113: std_logic; attribute dont_touch of WX11113: signal is true;
	signal WX11114: std_logic; attribute dont_touch of WX11114: signal is true;
	signal WX11115: std_logic; attribute dont_touch of WX11115: signal is true;
	signal WX11116: std_logic; attribute dont_touch of WX11116: signal is true;
	signal WX11117: std_logic; attribute dont_touch of WX11117: signal is true;
	signal WX11118: std_logic; attribute dont_touch of WX11118: signal is true;
	signal WX11119: std_logic; attribute dont_touch of WX11119: signal is true;
	signal WX11120: std_logic; attribute dont_touch of WX11120: signal is true;
	signal WX11121: std_logic; attribute dont_touch of WX11121: signal is true;
	signal WX11122: std_logic; attribute dont_touch of WX11122: signal is true;
	signal WX11123: std_logic; attribute dont_touch of WX11123: signal is true;
	signal WX11124: std_logic; attribute dont_touch of WX11124: signal is true;
	signal WX11125: std_logic; attribute dont_touch of WX11125: signal is true;
	signal WX11126: std_logic; attribute dont_touch of WX11126: signal is true;
	signal WX11127: std_logic; attribute dont_touch of WX11127: signal is true;
	signal WX11128: std_logic; attribute dont_touch of WX11128: signal is true;
	signal WX11129: std_logic; attribute dont_touch of WX11129: signal is true;
	signal WX11130: std_logic; attribute dont_touch of WX11130: signal is true;
	signal WX11131: std_logic; attribute dont_touch of WX11131: signal is true;
	signal WX11132: std_logic; attribute dont_touch of WX11132: signal is true;
	signal WX11133: std_logic; attribute dont_touch of WX11133: signal is true;
	signal WX11134: std_logic; attribute dont_touch of WX11134: signal is true;
	signal WX11135: std_logic; attribute dont_touch of WX11135: signal is true;
	signal WX11136: std_logic; attribute dont_touch of WX11136: signal is true;
	signal WX11137: std_logic; attribute dont_touch of WX11137: signal is true;
	signal WX11138: std_logic; attribute dont_touch of WX11138: signal is true;
	signal WX11139: std_logic; attribute dont_touch of WX11139: signal is true;
	signal WX11140: std_logic; attribute dont_touch of WX11140: signal is true;
	signal WX11141: std_logic; attribute dont_touch of WX11141: signal is true;
	signal WX11142: std_logic; attribute dont_touch of WX11142: signal is true;
	signal WX11143: std_logic; attribute dont_touch of WX11143: signal is true;
	signal WX11144: std_logic; attribute dont_touch of WX11144: signal is true;
	signal WX11145: std_logic; attribute dont_touch of WX11145: signal is true;
	signal WX11146: std_logic; attribute dont_touch of WX11146: signal is true;
	signal WX11147: std_logic; attribute dont_touch of WX11147: signal is true;
	signal WX11148: std_logic; attribute dont_touch of WX11148: signal is true;
	signal WX11149: std_logic; attribute dont_touch of WX11149: signal is true;
	signal WX11150: std_logic; attribute dont_touch of WX11150: signal is true;
	signal WX11151: std_logic; attribute dont_touch of WX11151: signal is true;
	signal WX11152: std_logic; attribute dont_touch of WX11152: signal is true;
	signal WX11153: std_logic; attribute dont_touch of WX11153: signal is true;
	signal WX11154: std_logic; attribute dont_touch of WX11154: signal is true;
	signal WX11155: std_logic; attribute dont_touch of WX11155: signal is true;
	signal WX11156: std_logic; attribute dont_touch of WX11156: signal is true;
	signal WX11157: std_logic; attribute dont_touch of WX11157: signal is true;
	signal WX11158: std_logic; attribute dont_touch of WX11158: signal is true;
	signal WX11159: std_logic; attribute dont_touch of WX11159: signal is true;
	signal WX11160: std_logic; attribute dont_touch of WX11160: signal is true;
	signal WX11161: std_logic; attribute dont_touch of WX11161: signal is true;
	signal WX11162: std_logic; attribute dont_touch of WX11162: signal is true;
	signal WX11163: std_logic; attribute dont_touch of WX11163: signal is true;
	signal WX11164: std_logic; attribute dont_touch of WX11164: signal is true;
	signal WX11165: std_logic; attribute dont_touch of WX11165: signal is true;
	signal WX11166: std_logic; attribute dont_touch of WX11166: signal is true;
	signal WX11167: std_logic; attribute dont_touch of WX11167: signal is true;
	signal WX11168: std_logic; attribute dont_touch of WX11168: signal is true;
	signal WX11169: std_logic; attribute dont_touch of WX11169: signal is true;
	signal WX11170: std_logic; attribute dont_touch of WX11170: signal is true;
	signal WX11171: std_logic; attribute dont_touch of WX11171: signal is true;
	signal WX11172: std_logic; attribute dont_touch of WX11172: signal is true;
	signal WX11173: std_logic; attribute dont_touch of WX11173: signal is true;
	signal WX11174: std_logic; attribute dont_touch of WX11174: signal is true;
	signal WX11175: std_logic; attribute dont_touch of WX11175: signal is true;
	signal WX11176: std_logic; attribute dont_touch of WX11176: signal is true;
	signal WX11177: std_logic; attribute dont_touch of WX11177: signal is true;
	signal WX11178: std_logic; attribute dont_touch of WX11178: signal is true;
	signal WX11179: std_logic; attribute dont_touch of WX11179: signal is true;
	signal WX11180: std_logic; attribute dont_touch of WX11180: signal is true;
	signal WX11181: std_logic; attribute dont_touch of WX11181: signal is true;
	signal WX11182: std_logic; attribute dont_touch of WX11182: signal is true;
	signal WX11183: std_logic; attribute dont_touch of WX11183: signal is true;
	signal WX11184: std_logic; attribute dont_touch of WX11184: signal is true;
	signal WX11185: std_logic; attribute dont_touch of WX11185: signal is true;
	signal WX11186: std_logic; attribute dont_touch of WX11186: signal is true;
	signal WX11187: std_logic; attribute dont_touch of WX11187: signal is true;
	signal WX11188: std_logic; attribute dont_touch of WX11188: signal is true;
	signal WX11189: std_logic; attribute dont_touch of WX11189: signal is true;
	signal WX11190: std_logic; attribute dont_touch of WX11190: signal is true;
	signal WX11191: std_logic; attribute dont_touch of WX11191: signal is true;
	signal WX11192: std_logic; attribute dont_touch of WX11192: signal is true;
	signal WX11193: std_logic; attribute dont_touch of WX11193: signal is true;
	signal WX11194: std_logic; attribute dont_touch of WX11194: signal is true;
	signal WX11195: std_logic; attribute dont_touch of WX11195: signal is true;
	signal WX11196: std_logic; attribute dont_touch of WX11196: signal is true;
	signal WX11197: std_logic; attribute dont_touch of WX11197: signal is true;
	signal WX11198: std_logic; attribute dont_touch of WX11198: signal is true;
	signal WX11199: std_logic; attribute dont_touch of WX11199: signal is true;
	signal WX11200: std_logic; attribute dont_touch of WX11200: signal is true;
	signal WX11201: std_logic; attribute dont_touch of WX11201: signal is true;
	signal WX11202: std_logic; attribute dont_touch of WX11202: signal is true;
	signal WX11203: std_logic; attribute dont_touch of WX11203: signal is true;
	signal WX11204: std_logic; attribute dont_touch of WX11204: signal is true;
	signal WX11205: std_logic; attribute dont_touch of WX11205: signal is true;
	signal WX11206: std_logic; attribute dont_touch of WX11206: signal is true;
	signal WX11207: std_logic; attribute dont_touch of WX11207: signal is true;
	signal WX11208: std_logic; attribute dont_touch of WX11208: signal is true;
	signal WX11209: std_logic; attribute dont_touch of WX11209: signal is true;
	signal WX11210: std_logic; attribute dont_touch of WX11210: signal is true;
	signal WX11211: std_logic; attribute dont_touch of WX11211: signal is true;
	signal WX11212: std_logic; attribute dont_touch of WX11212: signal is true;
	signal WX11213: std_logic; attribute dont_touch of WX11213: signal is true;
	signal WX11214: std_logic; attribute dont_touch of WX11214: signal is true;
	signal WX11215: std_logic; attribute dont_touch of WX11215: signal is true;
	signal WX11216: std_logic; attribute dont_touch of WX11216: signal is true;
	signal WX11217: std_logic; attribute dont_touch of WX11217: signal is true;
	signal WX11218: std_logic; attribute dont_touch of WX11218: signal is true;
	signal WX11219: std_logic; attribute dont_touch of WX11219: signal is true;
	signal WX11220: std_logic; attribute dont_touch of WX11220: signal is true;
	signal WX11221: std_logic; attribute dont_touch of WX11221: signal is true;
	signal WX11222: std_logic; attribute dont_touch of WX11222: signal is true;
	signal WX11223: std_logic; attribute dont_touch of WX11223: signal is true;
	signal WX11224: std_logic; attribute dont_touch of WX11224: signal is true;
	signal WX11225: std_logic; attribute dont_touch of WX11225: signal is true;
	signal WX11226: std_logic; attribute dont_touch of WX11226: signal is true;
	signal WX11227: std_logic; attribute dont_touch of WX11227: signal is true;
	signal WX11228: std_logic; attribute dont_touch of WX11228: signal is true;
	signal WX11229: std_logic; attribute dont_touch of WX11229: signal is true;
	signal WX11230: std_logic; attribute dont_touch of WX11230: signal is true;
	signal WX11231: std_logic; attribute dont_touch of WX11231: signal is true;
	signal WX11232: std_logic; attribute dont_touch of WX11232: signal is true;
	signal WX11233: std_logic; attribute dont_touch of WX11233: signal is true;
	signal WX11234: std_logic; attribute dont_touch of WX11234: signal is true;
	signal WX11235: std_logic; attribute dont_touch of WX11235: signal is true;
	signal WX11236: std_logic; attribute dont_touch of WX11236: signal is true;
	signal WX11237: std_logic; attribute dont_touch of WX11237: signal is true;
	signal WX11238: std_logic; attribute dont_touch of WX11238: signal is true;
	signal WX11239: std_logic; attribute dont_touch of WX11239: signal is true;
	signal WX11240: std_logic; attribute dont_touch of WX11240: signal is true;
	signal WX11241: std_logic; attribute dont_touch of WX11241: signal is true;
	signal WX11242: std_logic; attribute dont_touch of WX11242: signal is true;
	signal WX11243: std_logic; attribute dont_touch of WX11243: signal is true;
	signal WX11244: std_logic; attribute dont_touch of WX11244: signal is true;
	signal WX11245: std_logic; attribute dont_touch of WX11245: signal is true;
	signal WX11246: std_logic; attribute dont_touch of WX11246: signal is true;
	signal WX11247: std_logic; attribute dont_touch of WX11247: signal is true;
	signal WX11248: std_logic; attribute dont_touch of WX11248: signal is true;
	signal WX11249: std_logic; attribute dont_touch of WX11249: signal is true;
	signal WX11250: std_logic; attribute dont_touch of WX11250: signal is true;
	signal WX11251: std_logic; attribute dont_touch of WX11251: signal is true;
	signal WX11252: std_logic; attribute dont_touch of WX11252: signal is true;
	signal WX11253: std_logic; attribute dont_touch of WX11253: signal is true;
	signal WX11254: std_logic; attribute dont_touch of WX11254: signal is true;
	signal WX11255: std_logic; attribute dont_touch of WX11255: signal is true;
	signal WX11256: std_logic; attribute dont_touch of WX11256: signal is true;
	signal WX11257: std_logic; attribute dont_touch of WX11257: signal is true;
	signal WX11258: std_logic; attribute dont_touch of WX11258: signal is true;
	signal WX11259: std_logic; attribute dont_touch of WX11259: signal is true;
	signal WX11260: std_logic; attribute dont_touch of WX11260: signal is true;
	signal WX11261: std_logic; attribute dont_touch of WX11261: signal is true;
	signal WX11262: std_logic; attribute dont_touch of WX11262: signal is true;
	signal WX11263: std_logic; attribute dont_touch of WX11263: signal is true;
	signal WX11264: std_logic; attribute dont_touch of WX11264: signal is true;
	signal WX11265: std_logic; attribute dont_touch of WX11265: signal is true;
	signal WX11266: std_logic; attribute dont_touch of WX11266: signal is true;
	signal WX11267: std_logic; attribute dont_touch of WX11267: signal is true;
	signal WX11268: std_logic; attribute dont_touch of WX11268: signal is true;
	signal WX11269: std_logic; attribute dont_touch of WX11269: signal is true;
	signal WX11270: std_logic; attribute dont_touch of WX11270: signal is true;
	signal WX11271: std_logic; attribute dont_touch of WX11271: signal is true;
	signal WX11272: std_logic; attribute dont_touch of WX11272: signal is true;
	signal WX11273: std_logic; attribute dont_touch of WX11273: signal is true;
	signal WX11274: std_logic; attribute dont_touch of WX11274: signal is true;
	signal WX11275: std_logic; attribute dont_touch of WX11275: signal is true;
	signal WX11276: std_logic; attribute dont_touch of WX11276: signal is true;
	signal WX11277: std_logic; attribute dont_touch of WX11277: signal is true;
	signal WX11278: std_logic; attribute dont_touch of WX11278: signal is true;
	signal WX11279: std_logic; attribute dont_touch of WX11279: signal is true;
	signal WX11280: std_logic; attribute dont_touch of WX11280: signal is true;
	signal WX11281: std_logic; attribute dont_touch of WX11281: signal is true;
	signal WX11282: std_logic; attribute dont_touch of WX11282: signal is true;
	signal WX11283: std_logic; attribute dont_touch of WX11283: signal is true;
	signal WX11284: std_logic; attribute dont_touch of WX11284: signal is true;
	signal WX11285: std_logic; attribute dont_touch of WX11285: signal is true;
	signal WX11286: std_logic; attribute dont_touch of WX11286: signal is true;
	signal WX11287: std_logic; attribute dont_touch of WX11287: signal is true;
	signal WX11288: std_logic; attribute dont_touch of WX11288: signal is true;
	signal WX11289: std_logic; attribute dont_touch of WX11289: signal is true;
	signal WX11290: std_logic; attribute dont_touch of WX11290: signal is true;
	signal WX11291: std_logic; attribute dont_touch of WX11291: signal is true;
	signal WX11292: std_logic; attribute dont_touch of WX11292: signal is true;
	signal WX11293: std_logic; attribute dont_touch of WX11293: signal is true;
	signal WX11294: std_logic; attribute dont_touch of WX11294: signal is true;
	signal WX11295: std_logic; attribute dont_touch of WX11295: signal is true;
	signal WX11296: std_logic; attribute dont_touch of WX11296: signal is true;
	signal WX11297: std_logic; attribute dont_touch of WX11297: signal is true;
	signal WX11298: std_logic; attribute dont_touch of WX11298: signal is true;
	signal WX11299: std_logic; attribute dont_touch of WX11299: signal is true;
	signal WX11300: std_logic; attribute dont_touch of WX11300: signal is true;
	signal WX11301: std_logic; attribute dont_touch of WX11301: signal is true;
	signal WX11302: std_logic; attribute dont_touch of WX11302: signal is true;
	signal WX11303: std_logic; attribute dont_touch of WX11303: signal is true;
	signal WX11304: std_logic; attribute dont_touch of WX11304: signal is true;
	signal WX11305: std_logic; attribute dont_touch of WX11305: signal is true;
	signal WX11306: std_logic; attribute dont_touch of WX11306: signal is true;
	signal WX11307: std_logic; attribute dont_touch of WX11307: signal is true;
	signal WX11308: std_logic; attribute dont_touch of WX11308: signal is true;
	signal WX11309: std_logic; attribute dont_touch of WX11309: signal is true;
	signal WX11310: std_logic; attribute dont_touch of WX11310: signal is true;
	signal WX11311: std_logic; attribute dont_touch of WX11311: signal is true;
	signal WX11312: std_logic; attribute dont_touch of WX11312: signal is true;
	signal WX11313: std_logic; attribute dont_touch of WX11313: signal is true;
	signal WX11314: std_logic; attribute dont_touch of WX11314: signal is true;
	signal WX11315: std_logic; attribute dont_touch of WX11315: signal is true;
	signal WX11316: std_logic; attribute dont_touch of WX11316: signal is true;
	signal WX11317: std_logic; attribute dont_touch of WX11317: signal is true;
	signal WX11318: std_logic; attribute dont_touch of WX11318: signal is true;
	signal WX11319: std_logic; attribute dont_touch of WX11319: signal is true;
	signal WX11320: std_logic; attribute dont_touch of WX11320: signal is true;
	signal WX11321: std_logic; attribute dont_touch of WX11321: signal is true;
	signal WX11322: std_logic; attribute dont_touch of WX11322: signal is true;
	signal WX11323: std_logic; attribute dont_touch of WX11323: signal is true;
	signal WX11324: std_logic; attribute dont_touch of WX11324: signal is true;
	signal WX11325: std_logic; attribute dont_touch of WX11325: signal is true;
	signal WX11326: std_logic; attribute dont_touch of WX11326: signal is true;
	signal WX11327: std_logic; attribute dont_touch of WX11327: signal is true;
	signal WX11328: std_logic; attribute dont_touch of WX11328: signal is true;
	signal WX11329: std_logic; attribute dont_touch of WX11329: signal is true;
	signal WX11330: std_logic; attribute dont_touch of WX11330: signal is true;
	signal WX11331: std_logic; attribute dont_touch of WX11331: signal is true;
	signal WX11332: std_logic; attribute dont_touch of WX11332: signal is true;
	signal WX11333: std_logic; attribute dont_touch of WX11333: signal is true;
	signal WX11334: std_logic; attribute dont_touch of WX11334: signal is true;
	signal WX11335: std_logic; attribute dont_touch of WX11335: signal is true;
	signal WX11336: std_logic; attribute dont_touch of WX11336: signal is true;
	signal WX11337: std_logic; attribute dont_touch of WX11337: signal is true;
	signal WX11338: std_logic; attribute dont_touch of WX11338: signal is true;
	signal WX11339: std_logic; attribute dont_touch of WX11339: signal is true;
	signal WX11340: std_logic; attribute dont_touch of WX11340: signal is true;
	signal WX11341: std_logic; attribute dont_touch of WX11341: signal is true;
	signal WX11342: std_logic; attribute dont_touch of WX11342: signal is true;
	signal WX11343: std_logic; attribute dont_touch of WX11343: signal is true;
	signal WX11344: std_logic; attribute dont_touch of WX11344: signal is true;
	signal WX11345: std_logic; attribute dont_touch of WX11345: signal is true;
	signal WX11346: std_logic; attribute dont_touch of WX11346: signal is true;
	signal WX11347: std_logic; attribute dont_touch of WX11347: signal is true;
	signal WX11348: std_logic; attribute dont_touch of WX11348: signal is true;
	signal WX11349: std_logic; attribute dont_touch of WX11349: signal is true;
	signal WX11350: std_logic; attribute dont_touch of WX11350: signal is true;
	signal WX11351: std_logic; attribute dont_touch of WX11351: signal is true;
	signal WX11352: std_logic; attribute dont_touch of WX11352: signal is true;
	signal WX11353: std_logic; attribute dont_touch of WX11353: signal is true;
	signal WX11354: std_logic; attribute dont_touch of WX11354: signal is true;
	signal WX11355: std_logic; attribute dont_touch of WX11355: signal is true;
	signal WX11356: std_logic; attribute dont_touch of WX11356: signal is true;
	signal WX11357: std_logic; attribute dont_touch of WX11357: signal is true;
	signal WX11358: std_logic; attribute dont_touch of WX11358: signal is true;
	signal WX11359: std_logic; attribute dont_touch of WX11359: signal is true;
	signal WX11360: std_logic; attribute dont_touch of WX11360: signal is true;
	signal WX11361: std_logic; attribute dont_touch of WX11361: signal is true;
	signal WX11362: std_logic; attribute dont_touch of WX11362: signal is true;
	signal WX11363: std_logic; attribute dont_touch of WX11363: signal is true;
	signal WX11364: std_logic; attribute dont_touch of WX11364: signal is true;
	signal WX11365: std_logic; attribute dont_touch of WX11365: signal is true;
	signal WX11366: std_logic; attribute dont_touch of WX11366: signal is true;
	signal WX11367: std_logic; attribute dont_touch of WX11367: signal is true;
	signal WX11368: std_logic; attribute dont_touch of WX11368: signal is true;
	signal WX11369: std_logic; attribute dont_touch of WX11369: signal is true;
	signal WX11370: std_logic; attribute dont_touch of WX11370: signal is true;
	signal WX11371: std_logic; attribute dont_touch of WX11371: signal is true;
	signal WX11372: std_logic; attribute dont_touch of WX11372: signal is true;
	signal WX11373: std_logic; attribute dont_touch of WX11373: signal is true;
	signal WX11374: std_logic; attribute dont_touch of WX11374: signal is true;
	signal WX11375: std_logic; attribute dont_touch of WX11375: signal is true;
	signal WX11376: std_logic; attribute dont_touch of WX11376: signal is true;
	signal WX11377: std_logic; attribute dont_touch of WX11377: signal is true;
	signal WX11378: std_logic; attribute dont_touch of WX11378: signal is true;
	signal WX11379: std_logic; attribute dont_touch of WX11379: signal is true;
	signal WX11380: std_logic; attribute dont_touch of WX11380: signal is true;
	signal WX11381: std_logic; attribute dont_touch of WX11381: signal is true;
	signal WX11382: std_logic; attribute dont_touch of WX11382: signal is true;
	signal WX11383: std_logic; attribute dont_touch of WX11383: signal is true;
	signal WX11384: std_logic; attribute dont_touch of WX11384: signal is true;
	signal WX11385: std_logic; attribute dont_touch of WX11385: signal is true;
	signal WX11386: std_logic; attribute dont_touch of WX11386: signal is true;
	signal WX11387: std_logic; attribute dont_touch of WX11387: signal is true;
	signal WX11388: std_logic; attribute dont_touch of WX11388: signal is true;
	signal WX11389: std_logic; attribute dont_touch of WX11389: signal is true;
	signal WX11390: std_logic; attribute dont_touch of WX11390: signal is true;
	signal WX11391: std_logic; attribute dont_touch of WX11391: signal is true;
	signal WX11392: std_logic; attribute dont_touch of WX11392: signal is true;
	signal WX11393: std_logic; attribute dont_touch of WX11393: signal is true;
	signal WX11394: std_logic; attribute dont_touch of WX11394: signal is true;
	signal WX11395: std_logic; attribute dont_touch of WX11395: signal is true;
	signal WX11396: std_logic; attribute dont_touch of WX11396: signal is true;
	signal WX11397: std_logic; attribute dont_touch of WX11397: signal is true;
	signal WX11398: std_logic; attribute dont_touch of WX11398: signal is true;
	signal WX11399: std_logic; attribute dont_touch of WX11399: signal is true;
	signal WX11400: std_logic; attribute dont_touch of WX11400: signal is true;
	signal WX11401: std_logic; attribute dont_touch of WX11401: signal is true;
	signal WX11402: std_logic; attribute dont_touch of WX11402: signal is true;
	signal WX11403: std_logic; attribute dont_touch of WX11403: signal is true;
	signal WX11404: std_logic; attribute dont_touch of WX11404: signal is true;
	signal WX11405: std_logic; attribute dont_touch of WX11405: signal is true;
	signal WX11406: std_logic; attribute dont_touch of WX11406: signal is true;
	signal WX11407: std_logic; attribute dont_touch of WX11407: signal is true;
	signal WX11408: std_logic; attribute dont_touch of WX11408: signal is true;
	signal WX11409: std_logic; attribute dont_touch of WX11409: signal is true;
	signal WX11410: std_logic; attribute dont_touch of WX11410: signal is true;
	signal WX11411: std_logic; attribute dont_touch of WX11411: signal is true;
	signal WX11412: std_logic; attribute dont_touch of WX11412: signal is true;
	signal WX11413: std_logic; attribute dont_touch of WX11413: signal is true;
	signal WX11414: std_logic; attribute dont_touch of WX11414: signal is true;
	signal WX11415: std_logic; attribute dont_touch of WX11415: signal is true;
	signal WX11416: std_logic; attribute dont_touch of WX11416: signal is true;
	signal WX11417: std_logic; attribute dont_touch of WX11417: signal is true;
	signal WX11418: std_logic; attribute dont_touch of WX11418: signal is true;
	signal WX11419: std_logic; attribute dont_touch of WX11419: signal is true;
	signal WX11420: std_logic; attribute dont_touch of WX11420: signal is true;
	signal WX11421: std_logic; attribute dont_touch of WX11421: signal is true;
	signal WX11422: std_logic; attribute dont_touch of WX11422: signal is true;
	signal WX11423: std_logic; attribute dont_touch of WX11423: signal is true;
	signal WX11424: std_logic; attribute dont_touch of WX11424: signal is true;
	signal WX11425: std_logic; attribute dont_touch of WX11425: signal is true;
	signal WX11426: std_logic; attribute dont_touch of WX11426: signal is true;
	signal WX11427: std_logic; attribute dont_touch of WX11427: signal is true;
	signal WX11428: std_logic; attribute dont_touch of WX11428: signal is true;
	signal WX11429: std_logic; attribute dont_touch of WX11429: signal is true;
	signal WX11430: std_logic; attribute dont_touch of WX11430: signal is true;
	signal WX11431: std_logic; attribute dont_touch of WX11431: signal is true;
	signal WX11432: std_logic; attribute dont_touch of WX11432: signal is true;
	signal WX11433: std_logic; attribute dont_touch of WX11433: signal is true;
	signal WX11434: std_logic; attribute dont_touch of WX11434: signal is true;
	signal WX11435: std_logic; attribute dont_touch of WX11435: signal is true;
	signal WX11436: std_logic; attribute dont_touch of WX11436: signal is true;
	signal WX11437: std_logic; attribute dont_touch of WX11437: signal is true;
	signal WX11438: std_logic; attribute dont_touch of WX11438: signal is true;
	signal WX11439: std_logic; attribute dont_touch of WX11439: signal is true;
	signal WX11440: std_logic; attribute dont_touch of WX11440: signal is true;
	signal WX11441: std_logic; attribute dont_touch of WX11441: signal is true;
	signal WX11442: std_logic; attribute dont_touch of WX11442: signal is true;
	signal WX11443: std_logic; attribute dont_touch of WX11443: signal is true;
	signal WX11444: std_logic; attribute dont_touch of WX11444: signal is true;
	signal WX11445: std_logic; attribute dont_touch of WX11445: signal is true;
	signal WX11446: std_logic; attribute dont_touch of WX11446: signal is true;
	signal WX11447: std_logic; attribute dont_touch of WX11447: signal is true;
	signal WX11448: std_logic; attribute dont_touch of WX11448: signal is true;
	signal WX11449: std_logic; attribute dont_touch of WX11449: signal is true;
	signal WX11450: std_logic; attribute dont_touch of WX11450: signal is true;
	signal WX11451: std_logic; attribute dont_touch of WX11451: signal is true;
	signal WX11452: std_logic; attribute dont_touch of WX11452: signal is true;
	signal WX11453: std_logic; attribute dont_touch of WX11453: signal is true;
	signal WX11454: std_logic; attribute dont_touch of WX11454: signal is true;
	signal WX11455: std_logic; attribute dont_touch of WX11455: signal is true;
	signal WX11456: std_logic; attribute dont_touch of WX11456: signal is true;
	signal WX11457: std_logic; attribute dont_touch of WX11457: signal is true;
	signal WX11458: std_logic; attribute dont_touch of WX11458: signal is true;
	signal WX11459: std_logic; attribute dont_touch of WX11459: signal is true;
	signal WX11460: std_logic; attribute dont_touch of WX11460: signal is true;
	signal WX11461: std_logic; attribute dont_touch of WX11461: signal is true;
	signal WX11462: std_logic; attribute dont_touch of WX11462: signal is true;
	signal WX11463: std_logic; attribute dont_touch of WX11463: signal is true;
	signal WX11464: std_logic; attribute dont_touch of WX11464: signal is true;
	signal WX11465: std_logic; attribute dont_touch of WX11465: signal is true;
	signal WX11466: std_logic; attribute dont_touch of WX11466: signal is true;
	signal WX11467: std_logic; attribute dont_touch of WX11467: signal is true;
	signal WX11468: std_logic; attribute dont_touch of WX11468: signal is true;
	signal WX11469: std_logic; attribute dont_touch of WX11469: signal is true;
	signal WX11470: std_logic; attribute dont_touch of WX11470: signal is true;
	signal WX11471: std_logic; attribute dont_touch of WX11471: signal is true;
	signal WX11472: std_logic; attribute dont_touch of WX11472: signal is true;
	signal WX11473: std_logic; attribute dont_touch of WX11473: signal is true;
	signal WX11474: std_logic; attribute dont_touch of WX11474: signal is true;
	signal WX11475: std_logic; attribute dont_touch of WX11475: signal is true;
	signal WX11476: std_logic; attribute dont_touch of WX11476: signal is true;
	signal WX11477: std_logic; attribute dont_touch of WX11477: signal is true;
	signal WX11478: std_logic; attribute dont_touch of WX11478: signal is true;
	signal WX11479: std_logic; attribute dont_touch of WX11479: signal is true;
	signal WX11480: std_logic; attribute dont_touch of WX11480: signal is true;
	signal WX11481: std_logic; attribute dont_touch of WX11481: signal is true;
	signal WX11482: std_logic; attribute dont_touch of WX11482: signal is true;
	signal WX11483: std_logic; attribute dont_touch of WX11483: signal is true;
	signal WX11484: std_logic; attribute dont_touch of WX11484: signal is true;
	signal WX11485: std_logic; attribute dont_touch of WX11485: signal is true;
	signal WX11486: std_logic; attribute dont_touch of WX11486: signal is true;
	signal WX11487: std_logic; attribute dont_touch of WX11487: signal is true;
	signal WX11488: std_logic; attribute dont_touch of WX11488: signal is true;
	signal WX11489: std_logic; attribute dont_touch of WX11489: signal is true;
	signal WX11490: std_logic; attribute dont_touch of WX11490: signal is true;
	signal WX11491: std_logic; attribute dont_touch of WX11491: signal is true;
	signal WX11492: std_logic; attribute dont_touch of WX11492: signal is true;
	signal WX11493: std_logic; attribute dont_touch of WX11493: signal is true;
	signal WX11494: std_logic; attribute dont_touch of WX11494: signal is true;
	signal WX11495: std_logic; attribute dont_touch of WX11495: signal is true;
	signal WX11496: std_logic; attribute dont_touch of WX11496: signal is true;
	signal WX11497: std_logic; attribute dont_touch of WX11497: signal is true;
	signal WX11498: std_logic; attribute dont_touch of WX11498: signal is true;
	signal WX11499: std_logic; attribute dont_touch of WX11499: signal is true;
	signal WX11500: std_logic; attribute dont_touch of WX11500: signal is true;
	signal WX11501: std_logic; attribute dont_touch of WX11501: signal is true;
	signal WX11502: std_logic; attribute dont_touch of WX11502: signal is true;
	signal WX11503: std_logic; attribute dont_touch of WX11503: signal is true;
	signal WX11504: std_logic; attribute dont_touch of WX11504: signal is true;
	signal WX11505: std_logic; attribute dont_touch of WX11505: signal is true;
	signal WX11506: std_logic; attribute dont_touch of WX11506: signal is true;
	signal WX11507: std_logic; attribute dont_touch of WX11507: signal is true;
	signal WX11508: std_logic; attribute dont_touch of WX11508: signal is true;
	signal WX11509: std_logic; attribute dont_touch of WX11509: signal is true;
	signal WX11510: std_logic; attribute dont_touch of WX11510: signal is true;
	signal WX11511: std_logic; attribute dont_touch of WX11511: signal is true;
	signal WX11512: std_logic; attribute dont_touch of WX11512: signal is true;
	signal WX11513: std_logic; attribute dont_touch of WX11513: signal is true;
	signal WX11514: std_logic; attribute dont_touch of WX11514: signal is true;
	signal WX11515: std_logic; attribute dont_touch of WX11515: signal is true;
	signal WX11516: std_logic; attribute dont_touch of WX11516: signal is true;
	signal WX11517: std_logic; attribute dont_touch of WX11517: signal is true;
	signal WX11518: std_logic; attribute dont_touch of WX11518: signal is true;
	signal WX11519: std_logic; attribute dont_touch of WX11519: signal is true;
	signal WX11520: std_logic; attribute dont_touch of WX11520: signal is true;
	signal WX11521: std_logic; attribute dont_touch of WX11521: signal is true;
	signal WX11522: std_logic; attribute dont_touch of WX11522: signal is true;
	signal WX11523: std_logic; attribute dont_touch of WX11523: signal is true;
	signal WX11524: std_logic; attribute dont_touch of WX11524: signal is true;
	signal WX11525: std_logic; attribute dont_touch of WX11525: signal is true;
	signal WX11526: std_logic; attribute dont_touch of WX11526: signal is true;
	signal WX11527: std_logic; attribute dont_touch of WX11527: signal is true;
	signal WX11528: std_logic; attribute dont_touch of WX11528: signal is true;
	signal WX11529: std_logic; attribute dont_touch of WX11529: signal is true;
	signal WX11530: std_logic; attribute dont_touch of WX11530: signal is true;
	signal WX11531: std_logic; attribute dont_touch of WX11531: signal is true;
	signal WX11532: std_logic; attribute dont_touch of WX11532: signal is true;
	signal WX11533: std_logic; attribute dont_touch of WX11533: signal is true;
	signal WX11534: std_logic; attribute dont_touch of WX11534: signal is true;
	signal WX11535: std_logic; attribute dont_touch of WX11535: signal is true;
	signal WX11536: std_logic; attribute dont_touch of WX11536: signal is true;
	signal WX11537: std_logic; attribute dont_touch of WX11537: signal is true;
	signal WX11538: std_logic; attribute dont_touch of WX11538: signal is true;
	signal WX11539: std_logic; attribute dont_touch of WX11539: signal is true;
	signal WX11540: std_logic; attribute dont_touch of WX11540: signal is true;
	signal WX11541: std_logic; attribute dont_touch of WX11541: signal is true;
	signal WX11542: std_logic; attribute dont_touch of WX11542: signal is true;
	signal WX11543: std_logic; attribute dont_touch of WX11543: signal is true;
	signal WX11544: std_logic; attribute dont_touch of WX11544: signal is true;
	signal WX11545: std_logic; attribute dont_touch of WX11545: signal is true;
	signal WX11546: std_logic; attribute dont_touch of WX11546: signal is true;
	signal WX11547: std_logic; attribute dont_touch of WX11547: signal is true;
	signal WX11548: std_logic; attribute dont_touch of WX11548: signal is true;
	signal WX11549: std_logic; attribute dont_touch of WX11549: signal is true;
	signal WX11550: std_logic; attribute dont_touch of WX11550: signal is true;
	signal WX11551: std_logic; attribute dont_touch of WX11551: signal is true;
	signal WX11552: std_logic; attribute dont_touch of WX11552: signal is true;
	signal WX11553: std_logic; attribute dont_touch of WX11553: signal is true;
	signal WX11554: std_logic; attribute dont_touch of WX11554: signal is true;
	signal WX11555: std_logic; attribute dont_touch of WX11555: signal is true;
	signal WX11556: std_logic; attribute dont_touch of WX11556: signal is true;
	signal WX11557: std_logic; attribute dont_touch of WX11557: signal is true;
	signal WX11558: std_logic; attribute dont_touch of WX11558: signal is true;
	signal WX11559: std_logic; attribute dont_touch of WX11559: signal is true;
	signal WX11560: std_logic; attribute dont_touch of WX11560: signal is true;
	signal WX11561: std_logic; attribute dont_touch of WX11561: signal is true;
	signal WX11562: std_logic; attribute dont_touch of WX11562: signal is true;
	signal WX11563: std_logic; attribute dont_touch of WX11563: signal is true;
	signal WX11564: std_logic; attribute dont_touch of WX11564: signal is true;
	signal WX11565: std_logic; attribute dont_touch of WX11565: signal is true;
	signal WX11566: std_logic; attribute dont_touch of WX11566: signal is true;
	signal WX11567: std_logic; attribute dont_touch of WX11567: signal is true;
	signal WX11568: std_logic; attribute dont_touch of WX11568: signal is true;
	signal WX11569: std_logic; attribute dont_touch of WX11569: signal is true;
	signal WX11570: std_logic; attribute dont_touch of WX11570: signal is true;
	signal WX11571: std_logic; attribute dont_touch of WX11571: signal is true;
	signal WX11572: std_logic; attribute dont_touch of WX11572: signal is true;
	signal WX11573: std_logic; attribute dont_touch of WX11573: signal is true;
	signal WX11574: std_logic; attribute dont_touch of WX11574: signal is true;
	signal WX11575: std_logic; attribute dont_touch of WX11575: signal is true;
	signal WX11576: std_logic; attribute dont_touch of WX11576: signal is true;
	signal WX11577: std_logic; attribute dont_touch of WX11577: signal is true;
	signal WX11578: std_logic; attribute dont_touch of WX11578: signal is true;
	signal WX11579: std_logic; attribute dont_touch of WX11579: signal is true;
	signal WX11580: std_logic; attribute dont_touch of WX11580: signal is true;
	signal WX11581: std_logic; attribute dont_touch of WX11581: signal is true;
	signal WX11582: std_logic; attribute dont_touch of WX11582: signal is true;
	signal WX11583: std_logic; attribute dont_touch of WX11583: signal is true;
	signal WX11584: std_logic; attribute dont_touch of WX11584: signal is true;
	signal WX11585: std_logic; attribute dont_touch of WX11585: signal is true;
	signal WX11586: std_logic; attribute dont_touch of WX11586: signal is true;
	signal WX11587: std_logic; attribute dont_touch of WX11587: signal is true;
	signal WX11588: std_logic; attribute dont_touch of WX11588: signal is true;
	signal WX11589: std_logic; attribute dont_touch of WX11589: signal is true;
	signal WX11590: std_logic; attribute dont_touch of WX11590: signal is true;
	signal WX11591: std_logic; attribute dont_touch of WX11591: signal is true;
	signal WX11592: std_logic; attribute dont_touch of WX11592: signal is true;
	signal WX11593: std_logic; attribute dont_touch of WX11593: signal is true;
	signal WX11594: std_logic; attribute dont_touch of WX11594: signal is true;
	signal WX11595: std_logic; attribute dont_touch of WX11595: signal is true;
	signal WX11596: std_logic; attribute dont_touch of WX11596: signal is true;
	signal WX11597: std_logic; attribute dont_touch of WX11597: signal is true;
	signal WX11598: std_logic; attribute dont_touch of WX11598: signal is true;
	signal WX11599: std_logic; attribute dont_touch of WX11599: signal is true;
	signal WX11600: std_logic; attribute dont_touch of WX11600: signal is true;
	signal WX11601: std_logic; attribute dont_touch of WX11601: signal is true;
	signal WX11602: std_logic; attribute dont_touch of WX11602: signal is true;
	signal WX11603: std_logic; attribute dont_touch of WX11603: signal is true;
	signal WX11604: std_logic; attribute dont_touch of WX11604: signal is true;
	signal WX11605: std_logic; attribute dont_touch of WX11605: signal is true;
	signal WX11606: std_logic; attribute dont_touch of WX11606: signal is true;
	signal WX11607: std_logic; attribute dont_touch of WX11607: signal is true;
	signal WX11608: std_logic; attribute dont_touch of WX11608: signal is true;
	signal WX11610: std_logic; attribute dont_touch of WX11610: signal is true;
	signal WX11612: std_logic; attribute dont_touch of WX11612: signal is true;
	signal WX11614: std_logic; attribute dont_touch of WX11614: signal is true;
	signal WX11616: std_logic; attribute dont_touch of WX11616: signal is true;
	signal WX11618: std_logic; attribute dont_touch of WX11618: signal is true;
	signal WX11620: std_logic; attribute dont_touch of WX11620: signal is true;
	signal WX11622: std_logic; attribute dont_touch of WX11622: signal is true;
	signal WX11624: std_logic; attribute dont_touch of WX11624: signal is true;
	signal WX11626: std_logic; attribute dont_touch of WX11626: signal is true;
	signal WX11628: std_logic; attribute dont_touch of WX11628: signal is true;
	signal WX11630: std_logic; attribute dont_touch of WX11630: signal is true;
	signal WX11632: std_logic; attribute dont_touch of WX11632: signal is true;
	signal WX11634: std_logic; attribute dont_touch of WX11634: signal is true;
	signal WX11636: std_logic; attribute dont_touch of WX11636: signal is true;
	signal WX11638: std_logic; attribute dont_touch of WX11638: signal is true;
	signal WX11640: std_logic; attribute dont_touch of WX11640: signal is true;
	signal WX11642: std_logic; attribute dont_touch of WX11642: signal is true;
	signal WX11644: std_logic; attribute dont_touch of WX11644: signal is true;
	signal WX11646: std_logic; attribute dont_touch of WX11646: signal is true;
	signal WX11648: std_logic; attribute dont_touch of WX11648: signal is true;
	signal WX11650: std_logic; attribute dont_touch of WX11650: signal is true;
	signal WX11652: std_logic; attribute dont_touch of WX11652: signal is true;
	signal WX11654: std_logic; attribute dont_touch of WX11654: signal is true;
	signal WX11656: std_logic; attribute dont_touch of WX11656: signal is true;
	signal WX11658: std_logic; attribute dont_touch of WX11658: signal is true;
	signal WX11660: std_logic; attribute dont_touch of WX11660: signal is true;
	signal WX11662: std_logic; attribute dont_touch of WX11662: signal is true;
	signal WX11664: std_logic; attribute dont_touch of WX11664: signal is true;
	signal WX11666: std_logic; attribute dont_touch of WX11666: signal is true;
	signal WX11668: std_logic; attribute dont_touch of WX11668: signal is true;
	signal WX11670: std_logic; attribute dont_touch of WX11670: signal is true;
begin
	process(CLK)
	begin
		if(rising_edge(CLK)) then
			CRC_OUT_1_0<=WX11608;
			CRC_OUT_1_1<=WX11610;
			CRC_OUT_1_2<=WX11612;
			CRC_OUT_1_3<=WX11614;
			CRC_OUT_1_4<=WX11616;
			CRC_OUT_1_5<=WX11618;
			CRC_OUT_1_6<=WX11620;
			CRC_OUT_1_7<=WX11622;
			CRC_OUT_1_8<=WX11624;
			CRC_OUT_1_9<=WX11626;
			CRC_OUT_1_10<=WX11628;
			CRC_OUT_1_11<=WX11630;
			CRC_OUT_1_12<=WX11632;
			CRC_OUT_1_13<=WX11634;
			CRC_OUT_1_14<=WX11636;
			CRC_OUT_1_15<=WX11638;
			CRC_OUT_1_16<=WX11640;
			CRC_OUT_1_17<=WX11642;
			CRC_OUT_1_18<=WX11644;
			CRC_OUT_1_19<=WX11646;
			CRC_OUT_1_20<=WX11648;
			CRC_OUT_1_21<=WX11650;
			CRC_OUT_1_22<=WX11652;
			CRC_OUT_1_23<=WX11654;
			CRC_OUT_1_24<=WX11656;
			CRC_OUT_1_25<=WX11658;
			CRC_OUT_1_26<=WX11660;
			CRC_OUT_1_27<=WX11662;
			CRC_OUT_1_28<=WX11664;
			CRC_OUT_1_29<=WX11666;
			CRC_OUT_1_30<=WX11668;
			CRC_OUT_1_31<=WX11670;
			CRC_OUT_2_0<=WX10315;
			CRC_OUT_2_1<=WX10317;
			CRC_OUT_2_2<=WX10319;
			CRC_OUT_2_3<=WX10321;
			CRC_OUT_2_4<=WX10323;
			CRC_OUT_2_5<=WX10325;
			CRC_OUT_2_6<=WX10327;
			CRC_OUT_2_7<=WX10329;
			CRC_OUT_2_8<=WX10331;
			CRC_OUT_2_9<=WX10333;
			CRC_OUT_2_10<=WX10335;
			CRC_OUT_2_11<=WX10337;
			CRC_OUT_2_12<=WX10339;
			CRC_OUT_2_13<=WX10341;
			CRC_OUT_2_14<=WX10343;
			CRC_OUT_2_15<=WX10345;
			CRC_OUT_2_16<=WX10347;
			CRC_OUT_2_17<=WX10349;
			CRC_OUT_2_18<=WX10351;
			CRC_OUT_2_19<=WX10353;
			CRC_OUT_2_20<=WX10355;
			CRC_OUT_2_21<=WX10357;
			CRC_OUT_2_22<=WX10359;
			CRC_OUT_2_23<=WX10361;
			CRC_OUT_2_24<=WX10363;
			CRC_OUT_2_25<=WX10365;
			CRC_OUT_2_26<=WX10367;
			CRC_OUT_2_27<=WX10369;
			CRC_OUT_2_28<=WX10371;
			CRC_OUT_2_29<=WX10373;
			CRC_OUT_2_30<=WX10375;
			CRC_OUT_2_31<=WX10377;
			CRC_OUT_3_0<=WX9022;
			CRC_OUT_3_1<=WX9024;
			CRC_OUT_3_2<=WX9026;
			CRC_OUT_3_3<=WX9028;
			CRC_OUT_3_4<=WX9030;
			CRC_OUT_3_5<=WX9032;
			CRC_OUT_3_6<=WX9034;
			CRC_OUT_3_7<=WX9036;
			CRC_OUT_3_8<=WX9038;
			CRC_OUT_3_9<=WX9040;
			CRC_OUT_3_10<=WX9042;
			CRC_OUT_3_11<=WX9044;
			CRC_OUT_3_12<=WX9046;
			CRC_OUT_3_13<=WX9048;
			CRC_OUT_3_14<=WX9050;
			CRC_OUT_3_15<=WX9052;
			CRC_OUT_3_16<=WX9054;
			CRC_OUT_3_17<=WX9056;
			CRC_OUT_3_18<=WX9058;
			CRC_OUT_3_19<=WX9060;
			CRC_OUT_3_20<=WX9062;
			CRC_OUT_3_21<=WX9064;
			CRC_OUT_3_22<=WX9066;
			CRC_OUT_3_23<=WX9068;
			CRC_OUT_3_24<=WX9070;
			CRC_OUT_3_25<=WX9072;
			CRC_OUT_3_26<=WX9074;
			CRC_OUT_3_27<=WX9076;
			CRC_OUT_3_28<=WX9078;
			CRC_OUT_3_29<=WX9080;
			CRC_OUT_3_30<=WX9082;
			CRC_OUT_3_31<=WX9084;
			CRC_OUT_4_0<=WX7729;
			CRC_OUT_4_1<=WX7731;
			CRC_OUT_4_2<=WX7733;
			CRC_OUT_4_3<=WX7735;
			CRC_OUT_4_4<=WX7737;
			CRC_OUT_4_5<=WX7739;
			CRC_OUT_4_6<=WX7741;
			CRC_OUT_4_7<=WX7743;
			CRC_OUT_4_8<=WX7745;
			CRC_OUT_4_9<=WX7747;
			CRC_OUT_4_10<=WX7749;
			CRC_OUT_4_11<=WX7751;
			CRC_OUT_4_12<=WX7753;
			CRC_OUT_4_13<=WX7755;
			CRC_OUT_4_14<=WX7757;
			CRC_OUT_4_15<=WX7759;
			CRC_OUT_4_16<=WX7761;
			CRC_OUT_4_17<=WX7763;
			CRC_OUT_4_18<=WX7765;
			CRC_OUT_4_19<=WX7767;
			CRC_OUT_4_20<=WX7769;
			CRC_OUT_4_21<=WX7771;
			CRC_OUT_4_22<=WX7773;
			CRC_OUT_4_23<=WX7775;
			CRC_OUT_4_24<=WX7777;
			CRC_OUT_4_25<=WX7779;
			CRC_OUT_4_26<=WX7781;
			CRC_OUT_4_27<=WX7783;
			CRC_OUT_4_28<=WX7785;
			CRC_OUT_4_29<=WX7787;
			CRC_OUT_4_30<=WX7789;
			CRC_OUT_4_31<=WX7791;
			CRC_OUT_5_0<=WX6436;
			CRC_OUT_5_1<=WX6438;
			CRC_OUT_5_2<=WX6440;
			CRC_OUT_5_3<=WX6442;
			CRC_OUT_5_4<=WX6444;
			CRC_OUT_5_5<=WX6446;
			CRC_OUT_5_6<=WX6448;
			CRC_OUT_5_7<=WX6450;
			CRC_OUT_5_8<=WX6452;
			CRC_OUT_5_9<=WX6454;
			CRC_OUT_5_10<=WX6456;
			CRC_OUT_5_11<=WX6458;
			CRC_OUT_5_12<=WX6460;
			CRC_OUT_5_13<=WX6462;
			CRC_OUT_5_14<=WX6464;
			CRC_OUT_5_15<=WX6466;
			CRC_OUT_5_16<=WX6468;
			CRC_OUT_5_17<=WX6470;
			CRC_OUT_5_18<=WX6472;
			CRC_OUT_5_19<=WX6474;
			CRC_OUT_5_20<=WX6476;
			CRC_OUT_5_21<=WX6478;
			CRC_OUT_5_22<=WX6480;
			CRC_OUT_5_23<=WX6482;
			CRC_OUT_5_24<=WX6484;
			CRC_OUT_5_25<=WX6486;
			CRC_OUT_5_26<=WX6488;
			CRC_OUT_5_27<=WX6490;
			CRC_OUT_5_28<=WX6492;
			CRC_OUT_5_29<=WX6494;
			CRC_OUT_5_30<=WX6496;
			CRC_OUT_5_31<=WX6498;
			CRC_OUT_6_0<=WX5143;
			CRC_OUT_6_1<=WX5145;
			CRC_OUT_6_2<=WX5147;
			CRC_OUT_6_3<=WX5149;
			CRC_OUT_6_4<=WX5151;
			CRC_OUT_6_5<=WX5153;
			CRC_OUT_6_6<=WX5155;
			CRC_OUT_6_7<=WX5157;
			CRC_OUT_6_8<=WX5159;
			CRC_OUT_6_9<=WX5161;
			CRC_OUT_6_10<=WX5163;
			CRC_OUT_6_11<=WX5165;
			CRC_OUT_6_12<=WX5167;
			CRC_OUT_6_13<=WX5169;
			CRC_OUT_6_14<=WX5171;
			CRC_OUT_6_15<=WX5173;
			CRC_OUT_6_16<=WX5175;
			CRC_OUT_6_17<=WX5177;
			CRC_OUT_6_18<=WX5179;
			CRC_OUT_6_19<=WX5181;
			CRC_OUT_6_20<=WX5183;
			CRC_OUT_6_21<=WX5185;
			CRC_OUT_6_22<=WX5187;
			CRC_OUT_6_23<=WX5189;
			CRC_OUT_6_24<=WX5191;
			CRC_OUT_6_25<=WX5193;
			CRC_OUT_6_26<=WX5195;
			CRC_OUT_6_27<=WX5197;
			CRC_OUT_6_28<=WX5199;
			CRC_OUT_6_29<=WX5201;
			CRC_OUT_6_30<=WX5203;
			CRC_OUT_6_31<=WX5205;
			CRC_OUT_7_0<=WX3850;
			CRC_OUT_7_1<=WX3852;
			CRC_OUT_7_2<=WX3854;
			CRC_OUT_7_3<=WX3856;
			CRC_OUT_7_4<=WX3858;
			CRC_OUT_7_5<=WX3860;
			CRC_OUT_7_6<=WX3862;
			CRC_OUT_7_7<=WX3864;
			CRC_OUT_7_8<=WX3866;
			CRC_OUT_7_9<=WX3868;
			CRC_OUT_7_10<=WX3870;
			CRC_OUT_7_11<=WX3872;
			CRC_OUT_7_12<=WX3874;
			CRC_OUT_7_13<=WX3876;
			CRC_OUT_7_14<=WX3878;
			CRC_OUT_7_15<=WX3880;
			CRC_OUT_7_16<=WX3882;
			CRC_OUT_7_17<=WX3884;
			CRC_OUT_7_18<=WX3886;
			CRC_OUT_7_19<=WX3888;
			CRC_OUT_7_20<=WX3890;
			CRC_OUT_7_21<=WX3892;
			CRC_OUT_7_22<=WX3894;
			CRC_OUT_7_23<=WX3896;
			CRC_OUT_7_24<=WX3898;
			CRC_OUT_7_25<=WX3900;
			CRC_OUT_7_26<=WX3902;
			CRC_OUT_7_27<=WX3904;
			CRC_OUT_7_28<=WX3906;
			CRC_OUT_7_29<=WX3908;
			CRC_OUT_7_30<=WX3910;
			CRC_OUT_7_31<=WX3912;
			CRC_OUT_8_0<=WX2557;
			CRC_OUT_8_1<=WX2559;
			CRC_OUT_8_2<=WX2561;
			CRC_OUT_8_3<=WX2563;
			CRC_OUT_8_4<=WX2565;
			CRC_OUT_8_5<=WX2567;
			CRC_OUT_8_6<=WX2569;
			CRC_OUT_8_7<=WX2571;
			CRC_OUT_8_8<=WX2573;
			CRC_OUT_8_9<=WX2575;
			CRC_OUT_8_10<=WX2577;
			CRC_OUT_8_11<=WX2579;
			CRC_OUT_8_12<=WX2581;
			CRC_OUT_8_13<=WX2583;
			CRC_OUT_8_14<=WX2585;
			CRC_OUT_8_15<=WX2587;
			CRC_OUT_8_16<=WX2589;
			CRC_OUT_8_17<=WX2591;
			CRC_OUT_8_18<=WX2593;
			CRC_OUT_8_19<=WX2595;
			CRC_OUT_8_20<=WX2597;
			CRC_OUT_8_21<=WX2599;
			CRC_OUT_8_22<=WX2601;
			CRC_OUT_8_23<=WX2603;
			CRC_OUT_8_24<=WX2605;
			CRC_OUT_8_25<=WX2607;
			CRC_OUT_8_26<=WX2609;
			CRC_OUT_8_27<=WX2611;
			CRC_OUT_8_28<=WX2613;
			CRC_OUT_8_29<=WX2615;
			CRC_OUT_8_30<=WX2617;
			CRC_OUT_8_31<=WX2619;
			CRC_OUT_9_0<=WX1264;
			CRC_OUT_9_1<=WX1266;
			CRC_OUT_9_2<=WX1268;
			CRC_OUT_9_3<=WX1270;
			CRC_OUT_9_4<=WX1272;
			CRC_OUT_9_5<=WX1274;
			CRC_OUT_9_6<=WX1276;
			CRC_OUT_9_7<=WX1278;
			CRC_OUT_9_8<=WX1280;
			CRC_OUT_9_9<=WX1282;
			CRC_OUT_9_10<=WX1284;
			CRC_OUT_9_11<=WX1286;
			CRC_OUT_9_12<=WX1288;
			CRC_OUT_9_13<=WX1290;
			CRC_OUT_9_14<=WX1292;
			CRC_OUT_9_15<=WX1294;
			CRC_OUT_9_16<=WX1296;
			CRC_OUT_9_17<=WX1298;
			CRC_OUT_9_18<=WX1300;
			CRC_OUT_9_19<=WX1302;
			CRC_OUT_9_20<=WX1304;
			CRC_OUT_9_21<=WX1306;
			CRC_OUT_9_22<=WX1308;
			CRC_OUT_9_23<=WX1310;
			CRC_OUT_9_24<=WX1312;
			CRC_OUT_9_25<=WX1314;
			CRC_OUT_9_26<=WX1316;
			CRC_OUT_9_27<=WX1318;
			CRC_OUT_9_28<=WX1320;
			CRC_OUT_9_29<=WX1322;
			CRC_OUT_9_30<=WX1324;
			CRC_OUT_9_31<=WX1326;
			WX485<=WX484;
			WX487<=WX486;
			WX489<=WX488;
			WX491<=WX490;
			WX493<=WX492;
			WX495<=WX494;
			WX497<=WX496;
			WX499<=WX498;
			WX501<=WX500;
			WX503<=WX502;
			WX505<=WX504;
			WX507<=WX506;
			WX509<=WX508;
			WX511<=WX510;
			WX513<=WX512;
			WX515<=WX514;
			WX517<=WX516;
			WX519<=WX518;
			WX521<=WX520;
			WX523<=WX522;
			WX525<=WX524;
			WX527<=WX526;
			WX529<=WX528;
			WX531<=WX530;
			WX533<=WX532;
			WX535<=WX534;
			WX537<=WX536;
			WX539<=WX538;
			WX541<=WX540;
			WX543<=WX542;
			WX545<=WX544;
			WX547<=WX546;
			WX645<=WX644;
			WX647<=WX646;
			WX649<=WX648;
			WX651<=WX650;
			WX653<=WX652;
			WX655<=WX654;
			WX657<=WX656;
			WX659<=WX658;
			WX661<=WX660;
			WX663<=WX662;
			WX665<=WX664;
			WX667<=WX666;
			WX669<=WX668;
			WX671<=WX670;
			WX673<=WX672;
			WX675<=WX674;
			WX677<=WX676;
			WX679<=WX678;
			WX681<=WX680;
			WX683<=WX682;
			WX685<=WX684;
			WX687<=WX686;
			WX689<=WX688;
			WX691<=WX690;
			WX693<=WX692;
			WX695<=WX694;
			WX697<=WX696;
			WX699<=WX698;
			WX701<=WX700;
			WX703<=WX702;
			WX705<=WX704;
			WX707<=WX706;
			WX709<=WX708;
			WX711<=WX710;
			WX713<=WX712;
			WX715<=WX714;
			WX717<=WX716;
			WX719<=WX718;
			WX721<=WX720;
			WX723<=WX722;
			WX725<=WX724;
			WX727<=WX726;
			WX729<=WX728;
			WX731<=WX730;
			WX733<=WX732;
			WX735<=WX734;
			WX737<=WX736;
			WX739<=WX738;
			WX741<=WX740;
			WX743<=WX742;
			WX745<=WX744;
			WX747<=WX746;
			WX749<=WX748;
			WX751<=WX750;
			WX753<=WX752;
			WX755<=WX754;
			WX757<=WX756;
			WX759<=WX758;
			WX761<=WX760;
			WX763<=WX762;
			WX765<=WX764;
			WX767<=WX766;
			WX769<=WX768;
			WX771<=WX770;
			WX773<=WX772;
			WX775<=WX774;
			WX777<=WX776;
			WX779<=WX778;
			WX781<=WX780;
			WX783<=WX782;
			WX785<=WX784;
			WX787<=WX786;
			WX789<=WX788;
			WX791<=WX790;
			WX793<=WX792;
			WX795<=WX794;
			WX797<=WX796;
			WX799<=WX798;
			WX801<=WX800;
			WX803<=WX802;
			WX805<=WX804;
			WX807<=WX806;
			WX809<=WX808;
			WX811<=WX810;
			WX813<=WX812;
			WX815<=WX814;
			WX817<=WX816;
			WX819<=WX818;
			WX821<=WX820;
			WX823<=WX822;
			WX825<=WX824;
			WX827<=WX826;
			WX829<=WX828;
			WX831<=WX830;
			WX833<=WX832;
			WX835<=WX834;
			WX837<=WX836;
			WX839<=WX838;
			WX841<=WX840;
			WX843<=WX842;
			WX845<=WX844;
			WX847<=WX846;
			WX849<=WX848;
			WX851<=WX850;
			WX853<=WX852;
			WX855<=WX854;
			WX857<=WX856;
			WX859<=WX858;
			WX861<=WX860;
			WX863<=WX862;
			WX865<=WX864;
			WX867<=WX866;
			WX869<=WX868;
			WX871<=WX870;
			WX873<=WX872;
			WX875<=WX874;
			WX877<=WX876;
			WX879<=WX878;
			WX881<=WX880;
			WX883<=WX882;
			WX885<=WX884;
			WX887<=WX886;
			WX889<=WX888;
			WX891<=WX890;
			WX893<=WX892;
			WX895<=WX894;
			WX897<=WX896;
			WX899<=WX898;
			WX1778<=WX1777;
			WX1780<=WX1779;
			WX1782<=WX1781;
			WX1784<=WX1783;
			WX1786<=WX1785;
			WX1788<=WX1787;
			WX1790<=WX1789;
			WX1792<=WX1791;
			WX1794<=WX1793;
			WX1796<=WX1795;
			WX1798<=WX1797;
			WX1800<=WX1799;
			WX1802<=WX1801;
			WX1804<=WX1803;
			WX1806<=WX1805;
			WX1808<=WX1807;
			WX1810<=WX1809;
			WX1812<=WX1811;
			WX1814<=WX1813;
			WX1816<=WX1815;
			WX1818<=WX1817;
			WX1820<=WX1819;
			WX1822<=WX1821;
			WX1824<=WX1823;
			WX1826<=WX1825;
			WX1828<=WX1827;
			WX1830<=WX1829;
			WX1832<=WX1831;
			WX1834<=WX1833;
			WX1836<=WX1835;
			WX1838<=WX1837;
			WX1840<=WX1839;
			WX1938<=WX1937;
			WX1940<=WX1939;
			WX1942<=WX1941;
			WX1944<=WX1943;
			WX1946<=WX1945;
			WX1948<=WX1947;
			WX1950<=WX1949;
			WX1952<=WX1951;
			WX1954<=WX1953;
			WX1956<=WX1955;
			WX1958<=WX1957;
			WX1960<=WX1959;
			WX1962<=WX1961;
			WX1964<=WX1963;
			WX1966<=WX1965;
			WX1968<=WX1967;
			WX1970<=WX1969;
			WX1972<=WX1971;
			WX1974<=WX1973;
			WX1976<=WX1975;
			WX1978<=WX1977;
			WX1980<=WX1979;
			WX1982<=WX1981;
			WX1984<=WX1983;
			WX1986<=WX1985;
			WX1988<=WX1987;
			WX1990<=WX1989;
			WX1992<=WX1991;
			WX1994<=WX1993;
			WX1996<=WX1995;
			WX1998<=WX1997;
			WX2000<=WX1999;
			WX2002<=WX2001;
			WX2004<=WX2003;
			WX2006<=WX2005;
			WX2008<=WX2007;
			WX2010<=WX2009;
			WX2012<=WX2011;
			WX2014<=WX2013;
			WX2016<=WX2015;
			WX2018<=WX2017;
			WX2020<=WX2019;
			WX2022<=WX2021;
			WX2024<=WX2023;
			WX2026<=WX2025;
			WX2028<=WX2027;
			WX2030<=WX2029;
			WX2032<=WX2031;
			WX2034<=WX2033;
			WX2036<=WX2035;
			WX2038<=WX2037;
			WX2040<=WX2039;
			WX2042<=WX2041;
			WX2044<=WX2043;
			WX2046<=WX2045;
			WX2048<=WX2047;
			WX2050<=WX2049;
			WX2052<=WX2051;
			WX2054<=WX2053;
			WX2056<=WX2055;
			WX2058<=WX2057;
			WX2060<=WX2059;
			WX2062<=WX2061;
			WX2064<=WX2063;
			WX2066<=WX2065;
			WX2068<=WX2067;
			WX2070<=WX2069;
			WX2072<=WX2071;
			WX2074<=WX2073;
			WX2076<=WX2075;
			WX2078<=WX2077;
			WX2080<=WX2079;
			WX2082<=WX2081;
			WX2084<=WX2083;
			WX2086<=WX2085;
			WX2088<=WX2087;
			WX2090<=WX2089;
			WX2092<=WX2091;
			WX2094<=WX2093;
			WX2096<=WX2095;
			WX2098<=WX2097;
			WX2100<=WX2099;
			WX2102<=WX2101;
			WX2104<=WX2103;
			WX2106<=WX2105;
			WX2108<=WX2107;
			WX2110<=WX2109;
			WX2112<=WX2111;
			WX2114<=WX2113;
			WX2116<=WX2115;
			WX2118<=WX2117;
			WX2120<=WX2119;
			WX2122<=WX2121;
			WX2124<=WX2123;
			WX2126<=WX2125;
			WX2128<=WX2127;
			WX2130<=WX2129;
			WX2132<=WX2131;
			WX2134<=WX2133;
			WX2136<=WX2135;
			WX2138<=WX2137;
			WX2140<=WX2139;
			WX2142<=WX2141;
			WX2144<=WX2143;
			WX2146<=WX2145;
			WX2148<=WX2147;
			WX2150<=WX2149;
			WX2152<=WX2151;
			WX2154<=WX2153;
			WX2156<=WX2155;
			WX2158<=WX2157;
			WX2160<=WX2159;
			WX2162<=WX2161;
			WX2164<=WX2163;
			WX2166<=WX2165;
			WX2168<=WX2167;
			WX2170<=WX2169;
			WX2172<=WX2171;
			WX2174<=WX2173;
			WX2176<=WX2175;
			WX2178<=WX2177;
			WX2180<=WX2179;
			WX2182<=WX2181;
			WX2184<=WX2183;
			WX2186<=WX2185;
			WX2188<=WX2187;
			WX2190<=WX2189;
			WX2192<=WX2191;
			WX3071<=WX3070;
			WX3073<=WX3072;
			WX3075<=WX3074;
			WX3077<=WX3076;
			WX3079<=WX3078;
			WX3081<=WX3080;
			WX3083<=WX3082;
			WX3085<=WX3084;
			WX3087<=WX3086;
			WX3089<=WX3088;
			WX3091<=WX3090;
			WX3093<=WX3092;
			WX3095<=WX3094;
			WX3097<=WX3096;
			WX3099<=WX3098;
			WX3101<=WX3100;
			WX3103<=WX3102;
			WX3105<=WX3104;
			WX3107<=WX3106;
			WX3109<=WX3108;
			WX3111<=WX3110;
			WX3113<=WX3112;
			WX3115<=WX3114;
			WX3117<=WX3116;
			WX3119<=WX3118;
			WX3121<=WX3120;
			WX3123<=WX3122;
			WX3125<=WX3124;
			WX3127<=WX3126;
			WX3129<=WX3128;
			WX3131<=WX3130;
			WX3133<=WX3132;
			WX3231<=WX3230;
			WX3233<=WX3232;
			WX3235<=WX3234;
			WX3237<=WX3236;
			WX3239<=WX3238;
			WX3241<=WX3240;
			WX3243<=WX3242;
			WX3245<=WX3244;
			WX3247<=WX3246;
			WX3249<=WX3248;
			WX3251<=WX3250;
			WX3253<=WX3252;
			WX3255<=WX3254;
			WX3257<=WX3256;
			WX3259<=WX3258;
			WX3261<=WX3260;
			WX3263<=WX3262;
			WX3265<=WX3264;
			WX3267<=WX3266;
			WX3269<=WX3268;
			WX3271<=WX3270;
			WX3273<=WX3272;
			WX3275<=WX3274;
			WX3277<=WX3276;
			WX3279<=WX3278;
			WX3281<=WX3280;
			WX3283<=WX3282;
			WX3285<=WX3284;
			WX3287<=WX3286;
			WX3289<=WX3288;
			WX3291<=WX3290;
			WX3293<=WX3292;
			WX3295<=WX3294;
			WX3297<=WX3296;
			WX3299<=WX3298;
			WX3301<=WX3300;
			WX3303<=WX3302;
			WX3305<=WX3304;
			WX3307<=WX3306;
			WX3309<=WX3308;
			WX3311<=WX3310;
			WX3313<=WX3312;
			WX3315<=WX3314;
			WX3317<=WX3316;
			WX3319<=WX3318;
			WX3321<=WX3320;
			WX3323<=WX3322;
			WX3325<=WX3324;
			WX3327<=WX3326;
			WX3329<=WX3328;
			WX3331<=WX3330;
			WX3333<=WX3332;
			WX3335<=WX3334;
			WX3337<=WX3336;
			WX3339<=WX3338;
			WX3341<=WX3340;
			WX3343<=WX3342;
			WX3345<=WX3344;
			WX3347<=WX3346;
			WX3349<=WX3348;
			WX3351<=WX3350;
			WX3353<=WX3352;
			WX3355<=WX3354;
			WX3357<=WX3356;
			WX3359<=WX3358;
			WX3361<=WX3360;
			WX3363<=WX3362;
			WX3365<=WX3364;
			WX3367<=WX3366;
			WX3369<=WX3368;
			WX3371<=WX3370;
			WX3373<=WX3372;
			WX3375<=WX3374;
			WX3377<=WX3376;
			WX3379<=WX3378;
			WX3381<=WX3380;
			WX3383<=WX3382;
			WX3385<=WX3384;
			WX3387<=WX3386;
			WX3389<=WX3388;
			WX3391<=WX3390;
			WX3393<=WX3392;
			WX3395<=WX3394;
			WX3397<=WX3396;
			WX3399<=WX3398;
			WX3401<=WX3400;
			WX3403<=WX3402;
			WX3405<=WX3404;
			WX3407<=WX3406;
			WX3409<=WX3408;
			WX3411<=WX3410;
			WX3413<=WX3412;
			WX3415<=WX3414;
			WX3417<=WX3416;
			WX3419<=WX3418;
			WX3421<=WX3420;
			WX3423<=WX3422;
			WX3425<=WX3424;
			WX3427<=WX3426;
			WX3429<=WX3428;
			WX3431<=WX3430;
			WX3433<=WX3432;
			WX3435<=WX3434;
			WX3437<=WX3436;
			WX3439<=WX3438;
			WX3441<=WX3440;
			WX3443<=WX3442;
			WX3445<=WX3444;
			WX3447<=WX3446;
			WX3449<=WX3448;
			WX3451<=WX3450;
			WX3453<=WX3452;
			WX3455<=WX3454;
			WX3457<=WX3456;
			WX3459<=WX3458;
			WX3461<=WX3460;
			WX3463<=WX3462;
			WX3465<=WX3464;
			WX3467<=WX3466;
			WX3469<=WX3468;
			WX3471<=WX3470;
			WX3473<=WX3472;
			WX3475<=WX3474;
			WX3477<=WX3476;
			WX3479<=WX3478;
			WX3481<=WX3480;
			WX3483<=WX3482;
			WX3485<=WX3484;
			WX4364<=WX4363;
			WX4366<=WX4365;
			WX4368<=WX4367;
			WX4370<=WX4369;
			WX4372<=WX4371;
			WX4374<=WX4373;
			WX4376<=WX4375;
			WX4378<=WX4377;
			WX4380<=WX4379;
			WX4382<=WX4381;
			WX4384<=WX4383;
			WX4386<=WX4385;
			WX4388<=WX4387;
			WX4390<=WX4389;
			WX4392<=WX4391;
			WX4394<=WX4393;
			WX4396<=WX4395;
			WX4398<=WX4397;
			WX4400<=WX4399;
			WX4402<=WX4401;
			WX4404<=WX4403;
			WX4406<=WX4405;
			WX4408<=WX4407;
			WX4410<=WX4409;
			WX4412<=WX4411;
			WX4414<=WX4413;
			WX4416<=WX4415;
			WX4418<=WX4417;
			WX4420<=WX4419;
			WX4422<=WX4421;
			WX4424<=WX4423;
			WX4426<=WX4425;
			WX4524<=WX4523;
			WX4526<=WX4525;
			WX4528<=WX4527;
			WX4530<=WX4529;
			WX4532<=WX4531;
			WX4534<=WX4533;
			WX4536<=WX4535;
			WX4538<=WX4537;
			WX4540<=WX4539;
			WX4542<=WX4541;
			WX4544<=WX4543;
			WX4546<=WX4545;
			WX4548<=WX4547;
			WX4550<=WX4549;
			WX4552<=WX4551;
			WX4554<=WX4553;
			WX4556<=WX4555;
			WX4558<=WX4557;
			WX4560<=WX4559;
			WX4562<=WX4561;
			WX4564<=WX4563;
			WX4566<=WX4565;
			WX4568<=WX4567;
			WX4570<=WX4569;
			WX4572<=WX4571;
			WX4574<=WX4573;
			WX4576<=WX4575;
			WX4578<=WX4577;
			WX4580<=WX4579;
			WX4582<=WX4581;
			WX4584<=WX4583;
			WX4586<=WX4585;
			WX4588<=WX4587;
			WX4590<=WX4589;
			WX4592<=WX4591;
			WX4594<=WX4593;
			WX4596<=WX4595;
			WX4598<=WX4597;
			WX4600<=WX4599;
			WX4602<=WX4601;
			WX4604<=WX4603;
			WX4606<=WX4605;
			WX4608<=WX4607;
			WX4610<=WX4609;
			WX4612<=WX4611;
			WX4614<=WX4613;
			WX4616<=WX4615;
			WX4618<=WX4617;
			WX4620<=WX4619;
			WX4622<=WX4621;
			WX4624<=WX4623;
			WX4626<=WX4625;
			WX4628<=WX4627;
			WX4630<=WX4629;
			WX4632<=WX4631;
			WX4634<=WX4633;
			WX4636<=WX4635;
			WX4638<=WX4637;
			WX4640<=WX4639;
			WX4642<=WX4641;
			WX4644<=WX4643;
			WX4646<=WX4645;
			WX4648<=WX4647;
			WX4650<=WX4649;
			WX4652<=WX4651;
			WX4654<=WX4653;
			WX4656<=WX4655;
			WX4658<=WX4657;
			WX4660<=WX4659;
			WX4662<=WX4661;
			WX4664<=WX4663;
			WX4666<=WX4665;
			WX4668<=WX4667;
			WX4670<=WX4669;
			WX4672<=WX4671;
			WX4674<=WX4673;
			WX4676<=WX4675;
			WX4678<=WX4677;
			WX4680<=WX4679;
			WX4682<=WX4681;
			WX4684<=WX4683;
			WX4686<=WX4685;
			WX4688<=WX4687;
			WX4690<=WX4689;
			WX4692<=WX4691;
			WX4694<=WX4693;
			WX4696<=WX4695;
			WX4698<=WX4697;
			WX4700<=WX4699;
			WX4702<=WX4701;
			WX4704<=WX4703;
			WX4706<=WX4705;
			WX4708<=WX4707;
			WX4710<=WX4709;
			WX4712<=WX4711;
			WX4714<=WX4713;
			WX4716<=WX4715;
			WX4718<=WX4717;
			WX4720<=WX4719;
			WX4722<=WX4721;
			WX4724<=WX4723;
			WX4726<=WX4725;
			WX4728<=WX4727;
			WX4730<=WX4729;
			WX4732<=WX4731;
			WX4734<=WX4733;
			WX4736<=WX4735;
			WX4738<=WX4737;
			WX4740<=WX4739;
			WX4742<=WX4741;
			WX4744<=WX4743;
			WX4746<=WX4745;
			WX4748<=WX4747;
			WX4750<=WX4749;
			WX4752<=WX4751;
			WX4754<=WX4753;
			WX4756<=WX4755;
			WX4758<=WX4757;
			WX4760<=WX4759;
			WX4762<=WX4761;
			WX4764<=WX4763;
			WX4766<=WX4765;
			WX4768<=WX4767;
			WX4770<=WX4769;
			WX4772<=WX4771;
			WX4774<=WX4773;
			WX4776<=WX4775;
			WX4778<=WX4777;
			WX5657<=WX5656;
			WX5659<=WX5658;
			WX5661<=WX5660;
			WX5663<=WX5662;
			WX5665<=WX5664;
			WX5667<=WX5666;
			WX5669<=WX5668;
			WX5671<=WX5670;
			WX5673<=WX5672;
			WX5675<=WX5674;
			WX5677<=WX5676;
			WX5679<=WX5678;
			WX5681<=WX5680;
			WX5683<=WX5682;
			WX5685<=WX5684;
			WX5687<=WX5686;
			WX5689<=WX5688;
			WX5691<=WX5690;
			WX5693<=WX5692;
			WX5695<=WX5694;
			WX5697<=WX5696;
			WX5699<=WX5698;
			WX5701<=WX5700;
			WX5703<=WX5702;
			WX5705<=WX5704;
			WX5707<=WX5706;
			WX5709<=WX5708;
			WX5711<=WX5710;
			WX5713<=WX5712;
			WX5715<=WX5714;
			WX5717<=WX5716;
			WX5719<=WX5718;
			WX5817<=WX5816;
			WX5819<=WX5818;
			WX5821<=WX5820;
			WX5823<=WX5822;
			WX5825<=WX5824;
			WX5827<=WX5826;
			WX5829<=WX5828;
			WX5831<=WX5830;
			WX5833<=WX5832;
			WX5835<=WX5834;
			WX5837<=WX5836;
			WX5839<=WX5838;
			WX5841<=WX5840;
			WX5843<=WX5842;
			WX5845<=WX5844;
			WX5847<=WX5846;
			WX5849<=WX5848;
			WX5851<=WX5850;
			WX5853<=WX5852;
			WX5855<=WX5854;
			WX5857<=WX5856;
			WX5859<=WX5858;
			WX5861<=WX5860;
			WX5863<=WX5862;
			WX5865<=WX5864;
			WX5867<=WX5866;
			WX5869<=WX5868;
			WX5871<=WX5870;
			WX5873<=WX5872;
			WX5875<=WX5874;
			WX5877<=WX5876;
			WX5879<=WX5878;
			WX5881<=WX5880;
			WX5883<=WX5882;
			WX5885<=WX5884;
			WX5887<=WX5886;
			WX5889<=WX5888;
			WX5891<=WX5890;
			WX5893<=WX5892;
			WX5895<=WX5894;
			WX5897<=WX5896;
			WX5899<=WX5898;
			WX5901<=WX5900;
			WX5903<=WX5902;
			WX5905<=WX5904;
			WX5907<=WX5906;
			WX5909<=WX5908;
			WX5911<=WX5910;
			WX5913<=WX5912;
			WX5915<=WX5914;
			WX5917<=WX5916;
			WX5919<=WX5918;
			WX5921<=WX5920;
			WX5923<=WX5922;
			WX5925<=WX5924;
			WX5927<=WX5926;
			WX5929<=WX5928;
			WX5931<=WX5930;
			WX5933<=WX5932;
			WX5935<=WX5934;
			WX5937<=WX5936;
			WX5939<=WX5938;
			WX5941<=WX5940;
			WX5943<=WX5942;
			WX5945<=WX5944;
			WX5947<=WX5946;
			WX5949<=WX5948;
			WX5951<=WX5950;
			WX5953<=WX5952;
			WX5955<=WX5954;
			WX5957<=WX5956;
			WX5959<=WX5958;
			WX5961<=WX5960;
			WX5963<=WX5962;
			WX5965<=WX5964;
			WX5967<=WX5966;
			WX5969<=WX5968;
			WX5971<=WX5970;
			WX5973<=WX5972;
			WX5975<=WX5974;
			WX5977<=WX5976;
			WX5979<=WX5978;
			WX5981<=WX5980;
			WX5983<=WX5982;
			WX5985<=WX5984;
			WX5987<=WX5986;
			WX5989<=WX5988;
			WX5991<=WX5990;
			WX5993<=WX5992;
			WX5995<=WX5994;
			WX5997<=WX5996;
			WX5999<=WX5998;
			WX6001<=WX6000;
			WX6003<=WX6002;
			WX6005<=WX6004;
			WX6007<=WX6006;
			WX6009<=WX6008;
			WX6011<=WX6010;
			WX6013<=WX6012;
			WX6015<=WX6014;
			WX6017<=WX6016;
			WX6019<=WX6018;
			WX6021<=WX6020;
			WX6023<=WX6022;
			WX6025<=WX6024;
			WX6027<=WX6026;
			WX6029<=WX6028;
			WX6031<=WX6030;
			WX6033<=WX6032;
			WX6035<=WX6034;
			WX6037<=WX6036;
			WX6039<=WX6038;
			WX6041<=WX6040;
			WX6043<=WX6042;
			WX6045<=WX6044;
			WX6047<=WX6046;
			WX6049<=WX6048;
			WX6051<=WX6050;
			WX6053<=WX6052;
			WX6055<=WX6054;
			WX6057<=WX6056;
			WX6059<=WX6058;
			WX6061<=WX6060;
			WX6063<=WX6062;
			WX6065<=WX6064;
			WX6067<=WX6066;
			WX6069<=WX6068;
			WX6071<=WX6070;
			WX6950<=WX6949;
			WX6952<=WX6951;
			WX6954<=WX6953;
			WX6956<=WX6955;
			WX6958<=WX6957;
			WX6960<=WX6959;
			WX6962<=WX6961;
			WX6964<=WX6963;
			WX6966<=WX6965;
			WX6968<=WX6967;
			WX6970<=WX6969;
			WX6972<=WX6971;
			WX6974<=WX6973;
			WX6976<=WX6975;
			WX6978<=WX6977;
			WX6980<=WX6979;
			WX6982<=WX6981;
			WX6984<=WX6983;
			WX6986<=WX6985;
			WX6988<=WX6987;
			WX6990<=WX6989;
			WX6992<=WX6991;
			WX6994<=WX6993;
			WX6996<=WX6995;
			WX6998<=WX6997;
			WX7000<=WX6999;
			WX7002<=WX7001;
			WX7004<=WX7003;
			WX7006<=WX7005;
			WX7008<=WX7007;
			WX7010<=WX7009;
			WX7012<=WX7011;
			WX7110<=WX7109;
			WX7112<=WX7111;
			WX7114<=WX7113;
			WX7116<=WX7115;
			WX7118<=WX7117;
			WX7120<=WX7119;
			WX7122<=WX7121;
			WX7124<=WX7123;
			WX7126<=WX7125;
			WX7128<=WX7127;
			WX7130<=WX7129;
			WX7132<=WX7131;
			WX7134<=WX7133;
			WX7136<=WX7135;
			WX7138<=WX7137;
			WX7140<=WX7139;
			WX7142<=WX7141;
			WX7144<=WX7143;
			WX7146<=WX7145;
			WX7148<=WX7147;
			WX7150<=WX7149;
			WX7152<=WX7151;
			WX7154<=WX7153;
			WX7156<=WX7155;
			WX7158<=WX7157;
			WX7160<=WX7159;
			WX7162<=WX7161;
			WX7164<=WX7163;
			WX7166<=WX7165;
			WX7168<=WX7167;
			WX7170<=WX7169;
			WX7172<=WX7171;
			WX7174<=WX7173;
			WX7176<=WX7175;
			WX7178<=WX7177;
			WX7180<=WX7179;
			WX7182<=WX7181;
			WX7184<=WX7183;
			WX7186<=WX7185;
			WX7188<=WX7187;
			WX7190<=WX7189;
			WX7192<=WX7191;
			WX7194<=WX7193;
			WX7196<=WX7195;
			WX7198<=WX7197;
			WX7200<=WX7199;
			WX7202<=WX7201;
			WX7204<=WX7203;
			WX7206<=WX7205;
			WX7208<=WX7207;
			WX7210<=WX7209;
			WX7212<=WX7211;
			WX7214<=WX7213;
			WX7216<=WX7215;
			WX7218<=WX7217;
			WX7220<=WX7219;
			WX7222<=WX7221;
			WX7224<=WX7223;
			WX7226<=WX7225;
			WX7228<=WX7227;
			WX7230<=WX7229;
			WX7232<=WX7231;
			WX7234<=WX7233;
			WX7236<=WX7235;
			WX7238<=WX7237;
			WX7240<=WX7239;
			WX7242<=WX7241;
			WX7244<=WX7243;
			WX7246<=WX7245;
			WX7248<=WX7247;
			WX7250<=WX7249;
			WX7252<=WX7251;
			WX7254<=WX7253;
			WX7256<=WX7255;
			WX7258<=WX7257;
			WX7260<=WX7259;
			WX7262<=WX7261;
			WX7264<=WX7263;
			WX7266<=WX7265;
			WX7268<=WX7267;
			WX7270<=WX7269;
			WX7272<=WX7271;
			WX7274<=WX7273;
			WX7276<=WX7275;
			WX7278<=WX7277;
			WX7280<=WX7279;
			WX7282<=WX7281;
			WX7284<=WX7283;
			WX7286<=WX7285;
			WX7288<=WX7287;
			WX7290<=WX7289;
			WX7292<=WX7291;
			WX7294<=WX7293;
			WX7296<=WX7295;
			WX7298<=WX7297;
			WX7300<=WX7299;
			WX7302<=WX7301;
			WX7304<=WX7303;
			WX7306<=WX7305;
			WX7308<=WX7307;
			WX7310<=WX7309;
			WX7312<=WX7311;
			WX7314<=WX7313;
			WX7316<=WX7315;
			WX7318<=WX7317;
			WX7320<=WX7319;
			WX7322<=WX7321;
			WX7324<=WX7323;
			WX7326<=WX7325;
			WX7328<=WX7327;
			WX7330<=WX7329;
			WX7332<=WX7331;
			WX7334<=WX7333;
			WX7336<=WX7335;
			WX7338<=WX7337;
			WX7340<=WX7339;
			WX7342<=WX7341;
			WX7344<=WX7343;
			WX7346<=WX7345;
			WX7348<=WX7347;
			WX7350<=WX7349;
			WX7352<=WX7351;
			WX7354<=WX7353;
			WX7356<=WX7355;
			WX7358<=WX7357;
			WX7360<=WX7359;
			WX7362<=WX7361;
			WX7364<=WX7363;
			WX8243<=WX8242;
			WX8245<=WX8244;
			WX8247<=WX8246;
			WX8249<=WX8248;
			WX8251<=WX8250;
			WX8253<=WX8252;
			WX8255<=WX8254;
			WX8257<=WX8256;
			WX8259<=WX8258;
			WX8261<=WX8260;
			WX8263<=WX8262;
			WX8265<=WX8264;
			WX8267<=WX8266;
			WX8269<=WX8268;
			WX8271<=WX8270;
			WX8273<=WX8272;
			WX8275<=WX8274;
			WX8277<=WX8276;
			WX8279<=WX8278;
			WX8281<=WX8280;
			WX8283<=WX8282;
			WX8285<=WX8284;
			WX8287<=WX8286;
			WX8289<=WX8288;
			WX8291<=WX8290;
			WX8293<=WX8292;
			WX8295<=WX8294;
			WX8297<=WX8296;
			WX8299<=WX8298;
			WX8301<=WX8300;
			WX8303<=WX8302;
			WX8305<=WX8304;
			WX8403<=WX8402;
			WX8405<=WX8404;
			WX8407<=WX8406;
			WX8409<=WX8408;
			WX8411<=WX8410;
			WX8413<=WX8412;
			WX8415<=WX8414;
			WX8417<=WX8416;
			WX8419<=WX8418;
			WX8421<=WX8420;
			WX8423<=WX8422;
			WX8425<=WX8424;
			WX8427<=WX8426;
			WX8429<=WX8428;
			WX8431<=WX8430;
			WX8433<=WX8432;
			WX8435<=WX8434;
			WX8437<=WX8436;
			WX8439<=WX8438;
			WX8441<=WX8440;
			WX8443<=WX8442;
			WX8445<=WX8444;
			WX8447<=WX8446;
			WX8449<=WX8448;
			WX8451<=WX8450;
			WX8453<=WX8452;
			WX8455<=WX8454;
			WX8457<=WX8456;
			WX8459<=WX8458;
			WX8461<=WX8460;
			WX8463<=WX8462;
			WX8465<=WX8464;
			WX8467<=WX8466;
			WX8469<=WX8468;
			WX8471<=WX8470;
			WX8473<=WX8472;
			WX8475<=WX8474;
			WX8477<=WX8476;
			WX8479<=WX8478;
			WX8481<=WX8480;
			WX8483<=WX8482;
			WX8485<=WX8484;
			WX8487<=WX8486;
			WX8489<=WX8488;
			WX8491<=WX8490;
			WX8493<=WX8492;
			WX8495<=WX8494;
			WX8497<=WX8496;
			WX8499<=WX8498;
			WX8501<=WX8500;
			WX8503<=WX8502;
			WX8505<=WX8504;
			WX8507<=WX8506;
			WX8509<=WX8508;
			WX8511<=WX8510;
			WX8513<=WX8512;
			WX8515<=WX8514;
			WX8517<=WX8516;
			WX8519<=WX8518;
			WX8521<=WX8520;
			WX8523<=WX8522;
			WX8525<=WX8524;
			WX8527<=WX8526;
			WX8529<=WX8528;
			WX8531<=WX8530;
			WX8533<=WX8532;
			WX8535<=WX8534;
			WX8537<=WX8536;
			WX8539<=WX8538;
			WX8541<=WX8540;
			WX8543<=WX8542;
			WX8545<=WX8544;
			WX8547<=WX8546;
			WX8549<=WX8548;
			WX8551<=WX8550;
			WX8553<=WX8552;
			WX8555<=WX8554;
			WX8557<=WX8556;
			WX8559<=WX8558;
			WX8561<=WX8560;
			WX8563<=WX8562;
			WX8565<=WX8564;
			WX8567<=WX8566;
			WX8569<=WX8568;
			WX8571<=WX8570;
			WX8573<=WX8572;
			WX8575<=WX8574;
			WX8577<=WX8576;
			WX8579<=WX8578;
			WX8581<=WX8580;
			WX8583<=WX8582;
			WX8585<=WX8584;
			WX8587<=WX8586;
			WX8589<=WX8588;
			WX8591<=WX8590;
			WX8593<=WX8592;
			WX8595<=WX8594;
			WX8597<=WX8596;
			WX8599<=WX8598;
			WX8601<=WX8600;
			WX8603<=WX8602;
			WX8605<=WX8604;
			WX8607<=WX8606;
			WX8609<=WX8608;
			WX8611<=WX8610;
			WX8613<=WX8612;
			WX8615<=WX8614;
			WX8617<=WX8616;
			WX8619<=WX8618;
			WX8621<=WX8620;
			WX8623<=WX8622;
			WX8625<=WX8624;
			WX8627<=WX8626;
			WX8629<=WX8628;
			WX8631<=WX8630;
			WX8633<=WX8632;
			WX8635<=WX8634;
			WX8637<=WX8636;
			WX8639<=WX8638;
			WX8641<=WX8640;
			WX8643<=WX8642;
			WX8645<=WX8644;
			WX8647<=WX8646;
			WX8649<=WX8648;
			WX8651<=WX8650;
			WX8653<=WX8652;
			WX8655<=WX8654;
			WX8657<=WX8656;
			WX9536<=WX9535;
			WX9538<=WX9537;
			WX9540<=WX9539;
			WX9542<=WX9541;
			WX9544<=WX9543;
			WX9546<=WX9545;
			WX9548<=WX9547;
			WX9550<=WX9549;
			WX9552<=WX9551;
			WX9554<=WX9553;
			WX9556<=WX9555;
			WX9558<=WX9557;
			WX9560<=WX9559;
			WX9562<=WX9561;
			WX9564<=WX9563;
			WX9566<=WX9565;
			WX9568<=WX9567;
			WX9570<=WX9569;
			WX9572<=WX9571;
			WX9574<=WX9573;
			WX9576<=WX9575;
			WX9578<=WX9577;
			WX9580<=WX9579;
			WX9582<=WX9581;
			WX9584<=WX9583;
			WX9586<=WX9585;
			WX9588<=WX9587;
			WX9590<=WX9589;
			WX9592<=WX9591;
			WX9594<=WX9593;
			WX9596<=WX9595;
			WX9598<=WX9597;
			WX9696<=WX9695;
			WX9698<=WX9697;
			WX9700<=WX9699;
			WX9702<=WX9701;
			WX9704<=WX9703;
			WX9706<=WX9705;
			WX9708<=WX9707;
			WX9710<=WX9709;
			WX9712<=WX9711;
			WX9714<=WX9713;
			WX9716<=WX9715;
			WX9718<=WX9717;
			WX9720<=WX9719;
			WX9722<=WX9721;
			WX9724<=WX9723;
			WX9726<=WX9725;
			WX9728<=WX9727;
			WX9730<=WX9729;
			WX9732<=WX9731;
			WX9734<=WX9733;
			WX9736<=WX9735;
			WX9738<=WX9737;
			WX9740<=WX9739;
			WX9742<=WX9741;
			WX9744<=WX9743;
			WX9746<=WX9745;
			WX9748<=WX9747;
			WX9750<=WX9749;
			WX9752<=WX9751;
			WX9754<=WX9753;
			WX9756<=WX9755;
			WX9758<=WX9757;
			WX9760<=WX9759;
			WX9762<=WX9761;
			WX9764<=WX9763;
			WX9766<=WX9765;
			WX9768<=WX9767;
			WX9770<=WX9769;
			WX9772<=WX9771;
			WX9774<=WX9773;
			WX9776<=WX9775;
			WX9778<=WX9777;
			WX9780<=WX9779;
			WX9782<=WX9781;
			WX9784<=WX9783;
			WX9786<=WX9785;
			WX9788<=WX9787;
			WX9790<=WX9789;
			WX9792<=WX9791;
			WX9794<=WX9793;
			WX9796<=WX9795;
			WX9798<=WX9797;
			WX9800<=WX9799;
			WX9802<=WX9801;
			WX9804<=WX9803;
			WX9806<=WX9805;
			WX9808<=WX9807;
			WX9810<=WX9809;
			WX9812<=WX9811;
			WX9814<=WX9813;
			WX9816<=WX9815;
			WX9818<=WX9817;
			WX9820<=WX9819;
			WX9822<=WX9821;
			WX9824<=WX9823;
			WX9826<=WX9825;
			WX9828<=WX9827;
			WX9830<=WX9829;
			WX9832<=WX9831;
			WX9834<=WX9833;
			WX9836<=WX9835;
			WX9838<=WX9837;
			WX9840<=WX9839;
			WX9842<=WX9841;
			WX9844<=WX9843;
			WX9846<=WX9845;
			WX9848<=WX9847;
			WX9850<=WX9849;
			WX9852<=WX9851;
			WX9854<=WX9853;
			WX9856<=WX9855;
			WX9858<=WX9857;
			WX9860<=WX9859;
			WX9862<=WX9861;
			WX9864<=WX9863;
			WX9866<=WX9865;
			WX9868<=WX9867;
			WX9870<=WX9869;
			WX9872<=WX9871;
			WX9874<=WX9873;
			WX9876<=WX9875;
			WX9878<=WX9877;
			WX9880<=WX9879;
			WX9882<=WX9881;
			WX9884<=WX9883;
			WX9886<=WX9885;
			WX9888<=WX9887;
			WX9890<=WX9889;
			WX9892<=WX9891;
			WX9894<=WX9893;
			WX9896<=WX9895;
			WX9898<=WX9897;
			WX9900<=WX9899;
			WX9902<=WX9901;
			WX9904<=WX9903;
			WX9906<=WX9905;
			WX9908<=WX9907;
			WX9910<=WX9909;
			WX9912<=WX9911;
			WX9914<=WX9913;
			WX9916<=WX9915;
			WX9918<=WX9917;
			WX9920<=WX9919;
			WX9922<=WX9921;
			WX9924<=WX9923;
			WX9926<=WX9925;
			WX9928<=WX9927;
			WX9930<=WX9929;
			WX9932<=WX9931;
			WX9934<=WX9933;
			WX9936<=WX9935;
			WX9938<=WX9937;
			WX9940<=WX9939;
			WX9942<=WX9941;
			WX9944<=WX9943;
			WX9946<=WX9945;
			WX9948<=WX9947;
			WX9950<=WX9949;
			WX10829<=WX10828;
			WX10831<=WX10830;
			WX10833<=WX10832;
			WX10835<=WX10834;
			WX10837<=WX10836;
			WX10839<=WX10838;
			WX10841<=WX10840;
			WX10843<=WX10842;
			WX10845<=WX10844;
			WX10847<=WX10846;
			WX10849<=WX10848;
			WX10851<=WX10850;
			WX10853<=WX10852;
			WX10855<=WX10854;
			WX10857<=WX10856;
			WX10859<=WX10858;
			WX10861<=WX10860;
			WX10863<=WX10862;
			WX10865<=WX10864;
			WX10867<=WX10866;
			WX10869<=WX10868;
			WX10871<=WX10870;
			WX10873<=WX10872;
			WX10875<=WX10874;
			WX10877<=WX10876;
			WX10879<=WX10878;
			WX10881<=WX10880;
			WX10883<=WX10882;
			WX10885<=WX10884;
			WX10887<=WX10886;
			WX10889<=WX10888;
			WX10891<=WX10890;
			WX10989<=WX10988;
			WX10991<=WX10990;
			WX10993<=WX10992;
			WX10995<=WX10994;
			WX10997<=WX10996;
			WX10999<=WX10998;
			WX11001<=WX11000;
			WX11003<=WX11002;
			WX11005<=WX11004;
			WX11007<=WX11006;
			WX11009<=WX11008;
			WX11011<=WX11010;
			WX11013<=WX11012;
			WX11015<=WX11014;
			WX11017<=WX11016;
			WX11019<=WX11018;
			WX11021<=WX11020;
			WX11023<=WX11022;
			WX11025<=WX11024;
			WX11027<=WX11026;
			WX11029<=WX11028;
			WX11031<=WX11030;
			WX11033<=WX11032;
			WX11035<=WX11034;
			WX11037<=WX11036;
			WX11039<=WX11038;
			WX11041<=WX11040;
			WX11043<=WX11042;
			WX11045<=WX11044;
			WX11047<=WX11046;
			WX11049<=WX11048;
			WX11051<=WX11050;
			WX11053<=WX11052;
			WX11055<=WX11054;
			WX11057<=WX11056;
			WX11059<=WX11058;
			WX11061<=WX11060;
			WX11063<=WX11062;
			WX11065<=WX11064;
			WX11067<=WX11066;
			WX11069<=WX11068;
			WX11071<=WX11070;
			WX11073<=WX11072;
			WX11075<=WX11074;
			WX11077<=WX11076;
			WX11079<=WX11078;
			WX11081<=WX11080;
			WX11083<=WX11082;
			WX11085<=WX11084;
			WX11087<=WX11086;
			WX11089<=WX11088;
			WX11091<=WX11090;
			WX11093<=WX11092;
			WX11095<=WX11094;
			WX11097<=WX11096;
			WX11099<=WX11098;
			WX11101<=WX11100;
			WX11103<=WX11102;
			WX11105<=WX11104;
			WX11107<=WX11106;
			WX11109<=WX11108;
			WX11111<=WX11110;
			WX11113<=WX11112;
			WX11115<=WX11114;
			WX11117<=WX11116;
			WX11119<=WX11118;
			WX11121<=WX11120;
			WX11123<=WX11122;
			WX11125<=WX11124;
			WX11127<=WX11126;
			WX11129<=WX11128;
			WX11131<=WX11130;
			WX11133<=WX11132;
			WX11135<=WX11134;
			WX11137<=WX11136;
			WX11139<=WX11138;
			WX11141<=WX11140;
			WX11143<=WX11142;
			WX11145<=WX11144;
			WX11147<=WX11146;
			WX11149<=WX11148;
			WX11151<=WX11150;
			WX11153<=WX11152;
			WX11155<=WX11154;
			WX11157<=WX11156;
			WX11159<=WX11158;
			WX11161<=WX11160;
			WX11163<=WX11162;
			WX11165<=WX11164;
			WX11167<=WX11166;
			WX11169<=WX11168;
			WX11171<=WX11170;
			WX11173<=WX11172;
			WX11175<=WX11174;
			WX11177<=WX11176;
			WX11179<=WX11178;
			WX11181<=WX11180;
			WX11183<=WX11182;
			WX11185<=WX11184;
			WX11187<=WX11186;
			WX11189<=WX11188;
			WX11191<=WX11190;
			WX11193<=WX11192;
			WX11195<=WX11194;
			WX11197<=WX11196;
			WX11199<=WX11198;
			WX11201<=WX11200;
			WX11203<=WX11202;
			WX11205<=WX11204;
			WX11207<=WX11206;
			WX11209<=WX11208;
			WX11211<=WX11210;
			WX11213<=WX11212;
			WX11215<=WX11214;
			WX11217<=WX11216;
			WX11219<=WX11218;
			WX11221<=WX11220;
			WX11223<=WX11222;
			WX11225<=WX11224;
			WX11227<=WX11226;
			WX11229<=WX11228;
			WX11231<=WX11230;
			WX11233<=WX11232;
			WX11235<=WX11234;
			WX11237<=WX11236;
			WX11239<=WX11238;
			WX11241<=WX11240;
			WX11243<=WX11242;
		end if;
	end process;
	DATA_9_0<= not WX1228;
	DATA_9_1<= not WX1221;
	DATA_9_2<= not WX1214;
	DATA_9_3<= not WX1207;
	DATA_9_4<= not WX1200;
	DATA_9_5<= not WX1193;
	DATA_9_6<= not WX1186;
	DATA_9_7<= not WX1179;
	DATA_9_8<= not WX1172;
	DATA_9_9<= not WX1165;
	DATA_9_10<= not WX1158;
	DATA_9_11<= not WX1151;
	DATA_9_12<= not WX1144;
	DATA_9_13<= not WX1137;
	DATA_9_14<= not WX1130;
	DATA_9_15<= not WX1123;
	DATA_9_16<= not WX1116;
	DATA_9_17<= not WX1109;
	DATA_9_18<= not WX1102;
	DATA_9_19<= not WX1095;
	DATA_9_20<= not WX1088;
	DATA_9_21<= not WX1081;
	DATA_9_22<= not WX1074;
	DATA_9_23<= not WX1067;
	DATA_9_24<= not WX1060;
	DATA_9_25<= not WX1053;
	DATA_9_26<= not WX1046;
	DATA_9_27<= not WX1039;
	DATA_9_28<= not WX1032;
	DATA_9_29<= not WX1025;
	DATA_9_30<= not WX1018;
	DATA_9_31<= not WX1011;
	WX37<= not WX1003;
	WX41<= not WX1004;
	WX45<= not WX1004;
	WX47<= not WX38;
	WX48<= not WX47;
	WX51<= not WX1003;
	WX55<= not WX1004;
	WX59<= not WX1004;
	WX61<= not WX52;
	WX62<= not WX61;
	WX65<= not WX1003;
	WX69<= not WX1004;
	WX73<= not WX1004;
	WX75<= not WX66;
	WX76<= not WX75;
	WX79<= not WX1003;
	WX83<= not WX1004;
	WX87<= not WX1004;
	WX89<= not WX80;
	WX90<= not WX89;
	WX93<= not WX1003;
	WX97<= not WX1004;
	WX101<= not WX1004;
	WX103<= not WX94;
	WX104<= not WX103;
	WX107<= not WX1003;
	WX111<= not WX1004;
	WX115<= not WX1004;
	WX117<= not WX108;
	WX118<= not WX117;
	WX121<= not WX1003;
	WX125<= not WX1004;
	WX129<= not WX1004;
	WX131<= not WX122;
	WX132<= not WX131;
	WX135<= not WX1003;
	WX139<= not WX1004;
	WX143<= not WX1004;
	WX145<= not WX136;
	WX146<= not WX145;
	WX149<= not WX1003;
	WX153<= not WX1004;
	WX157<= not WX1004;
	WX159<= not WX150;
	WX160<= not WX159;
	WX163<= not WX1003;
	WX167<= not WX1004;
	WX171<= not WX1004;
	WX173<= not WX164;
	WX174<= not WX173;
	WX177<= not WX1003;
	WX181<= not WX1004;
	WX185<= not WX1004;
	WX187<= not WX178;
	WX188<= not WX187;
	WX191<= not WX1003;
	WX195<= not WX1004;
	WX199<= not WX1004;
	WX201<= not WX192;
	WX202<= not WX201;
	WX205<= not WX1003;
	WX209<= not WX1004;
	WX213<= not WX1004;
	WX215<= not WX206;
	WX216<= not WX215;
	WX219<= not WX1003;
	WX223<= not WX1004;
	WX227<= not WX1004;
	WX229<= not WX220;
	WX230<= not WX229;
	WX233<= not WX1003;
	WX237<= not WX1004;
	WX241<= not WX1004;
	WX243<= not WX234;
	WX244<= not WX243;
	WX247<= not WX1003;
	WX251<= not WX1004;
	WX255<= not WX1004;
	WX257<= not WX248;
	WX258<= not WX257;
	WX261<= not WX1003;
	WX265<= not WX1004;
	WX269<= not WX1004;
	WX271<= not WX262;
	WX272<= not WX271;
	WX275<= not WX1003;
	WX279<= not WX1004;
	WX283<= not WX1004;
	WX285<= not WX276;
	WX286<= not WX285;
	WX289<= not WX1003;
	WX293<= not WX1004;
	WX297<= not WX1004;
	WX299<= not WX290;
	WX300<= not WX299;
	WX303<= not WX1003;
	WX307<= not WX1004;
	WX311<= not WX1004;
	WX313<= not WX304;
	WX314<= not WX313;
	WX317<= not WX1003;
	WX321<= not WX1004;
	WX325<= not WX1004;
	WX327<= not WX318;
	WX328<= not WX327;
	WX331<= not WX1003;
	WX335<= not WX1004;
	WX339<= not WX1004;
	WX341<= not WX332;
	WX342<= not WX341;
	WX345<= not WX1003;
	WX349<= not WX1004;
	WX353<= not WX1004;
	WX355<= not WX346;
	WX356<= not WX355;
	WX359<= not WX1003;
	WX363<= not WX1004;
	WX367<= not WX1004;
	WX369<= not WX360;
	WX370<= not WX369;
	WX373<= not WX1003;
	WX377<= not WX1004;
	WX381<= not WX1004;
	WX383<= not WX374;
	WX384<= not WX383;
	WX387<= not WX1003;
	WX391<= not WX1004;
	WX395<= not WX1004;
	WX397<= not WX388;
	WX398<= not WX397;
	WX401<= not WX1003;
	WX405<= not WX1004;
	WX409<= not WX1004;
	WX411<= not WX402;
	WX412<= not WX411;
	WX415<= not WX1003;
	WX419<= not WX1004;
	WX423<= not WX1004;
	WX425<= not WX416;
	WX426<= not WX425;
	WX429<= not WX1003;
	WX433<= not WX1004;
	WX437<= not WX1004;
	WX439<= not WX430;
	WX440<= not WX439;
	WX443<= not WX1003;
	WX447<= not WX1004;
	WX451<= not WX1004;
	WX453<= not WX444;
	WX454<= not WX453;
	WX457<= not WX1003;
	WX461<= not WX1004;
	WX465<= not WX1004;
	WX467<= not WX458;
	WX468<= not WX467;
	WX471<= not WX1003;
	WX475<= not WX1004;
	WX479<= not WX1004;
	WX481<= not WX472;
	WX482<= not WX481;
	WX483<= not WX485;
	WX548<= not WX965;
	WX549<= not WX967;
	WX550<= not WX969;
	WX551<= not WX971;
	WX552<= not WX973;
	WX553<= not WX975;
	WX554<= not WX977;
	WX555<= not WX979;
	WX556<= not WX981;
	WX557<= not WX983;
	WX558<= not WX985;
	WX559<= not WX987;
	WX560<= not WX989;
	WX561<= not WX991;
	WX562<= not WX993;
	WX563<= not WX995;
	WX564<= not WX933;
	WX565<= not WX935;
	WX566<= not WX937;
	WX567<= not WX939;
	WX568<= not WX941;
	WX569<= not WX943;
	WX570<= not WX945;
	WX571<= not WX947;
	WX572<= not WX949;
	WX573<= not WX951;
	WX574<= not WX953;
	WX575<= not WX955;
	WX576<= not WX957;
	WX577<= not WX959;
	WX578<= not WX961;
	WX579<= not WX963;
	WX580<= not WX548;
	WX581<= not WX549;
	WX582<= not WX550;
	WX583<= not WX551;
	WX584<= not WX552;
	WX585<= not WX553;
	WX586<= not WX554;
	WX587<= not WX555;
	WX588<= not WX556;
	WX589<= not WX557;
	WX590<= not WX558;
	WX591<= not WX559;
	WX592<= not WX560;
	WX593<= not WX561;
	WX594<= not WX562;
	WX595<= not WX563;
	WX596<= not WX564;
	WX597<= not WX565;
	WX598<= not WX566;
	WX599<= not WX567;
	WX600<= not WX568;
	WX601<= not WX569;
	WX602<= not WX570;
	WX603<= not WX571;
	WX604<= not WX572;
	WX605<= not WX573;
	WX606<= not WX574;
	WX607<= not WX575;
	WX608<= not WX576;
	WX609<= not WX577;
	WX610<= not WX578;
	WX611<= not WX579;
	WX612<= not WX837;
	WX613<= not WX839;
	WX614<= not WX841;
	WX615<= not WX843;
	WX616<= not WX845;
	WX617<= not WX847;
	WX618<= not WX849;
	WX619<= not WX851;
	WX620<= not WX853;
	WX621<= not WX855;
	WX622<= not WX857;
	WX623<= not WX859;
	WX624<= not WX861;
	WX625<= not WX863;
	WX626<= not WX865;
	WX627<= not WX867;
	WX628<= not WX869;
	WX629<= not WX871;
	WX630<= not WX873;
	WX631<= not WX875;
	WX632<= not WX877;
	WX633<= not WX879;
	WX634<= not WX881;
	WX635<= not WX883;
	WX636<= not WX885;
	WX637<= not WX887;
	WX638<= not WX889;
	WX639<= not WX891;
	WX640<= not WX893;
	WX641<= not WX895;
	WX642<= not WX897;
	WX643<= not WX899;
	WX932<= not WX916;
	WX933<= not WX932;
	WX934<= not WX917;
	WX935<= not WX934;
	WX936<= not WX918;
	WX937<= not WX936;
	WX938<= not WX919;
	WX939<= not WX938;
	WX940<= not WX920;
	WX941<= not WX940;
	WX942<= not WX921;
	WX943<= not WX942;
	WX944<= not WX922;
	WX945<= not WX944;
	WX946<= not WX923;
	WX947<= not WX946;
	WX948<= not WX924;
	WX949<= not WX948;
	WX950<= not WX925;
	WX951<= not WX950;
	WX952<= not WX926;
	WX953<= not WX952;
	WX954<= not WX927;
	WX955<= not WX954;
	WX956<= not WX928;
	WX957<= not WX956;
	WX958<= not WX929;
	WX959<= not WX958;
	WX960<= not WX930;
	WX961<= not WX960;
	WX962<= not WX931;
	WX963<= not WX962;
	WX964<= not WX900;
	WX965<= not WX964;
	WX966<= not WX901;
	WX967<= not WX966;
	WX968<= not WX902;
	WX969<= not WX968;
	WX970<= not WX903;
	WX971<= not WX970;
	WX972<= not WX904;
	WX973<= not WX972;
	WX974<= not WX905;
	WX975<= not WX974;
	WX976<= not WX906;
	WX977<= not WX976;
	WX978<= not WX907;
	WX979<= not WX978;
	WX980<= not WX908;
	WX981<= not WX980;
	WX982<= not WX909;
	WX983<= not WX982;
	WX984<= not WX910;
	WX985<= not WX984;
	WX986<= not WX911;
	WX987<= not WX986;
	WX988<= not WX912;
	WX989<= not WX988;
	WX990<= not WX913;
	WX991<= not WX990;
	WX992<= not WX914;
	WX993<= not WX992;
	WX994<= not WX915;
	WX995<= not WX994;
	WX996<= not TM0;
	WX997<= not TM0;
	WX998<= not TM0;
	WX999<= not TM1;
	WX1000<= not TM1;
	WX1001<= not WX1000;
	WX1002<= not WX998;
	WX1003<= not WX999;
	WX1004<= not WX997;
	WX1005<= not WX996;
	WX1009<= not WX1005;
	WX1011<= not WX1010;
	WX1016<= not WX1005;
	WX1018<= not WX1017;
	WX1023<= not WX1005;
	WX1025<= not WX1024;
	WX1030<= not WX1005;
	WX1032<= not WX1031;
	WX1037<= not WX1005;
	WX1039<= not WX1038;
	WX1044<= not WX1005;
	WX1046<= not WX1045;
	WX1051<= not WX1005;
	WX1053<= not WX1052;
	WX1058<= not WX1005;
	WX1060<= not WX1059;
	WX1065<= not WX1005;
	WX1067<= not WX1066;
	WX1072<= not WX1005;
	WX1074<= not WX1073;
	WX1079<= not WX1005;
	WX1081<= not WX1080;
	WX1086<= not WX1005;
	WX1088<= not WX1087;
	WX1093<= not WX1005;
	WX1095<= not WX1094;
	WX1100<= not WX1005;
	WX1102<= not WX1101;
	WX1107<= not WX1005;
	WX1109<= not WX1108;
	WX1114<= not WX1005;
	WX1116<= not WX1115;
	WX1121<= not WX1005;
	WX1123<= not WX1122;
	WX1128<= not WX1005;
	WX1130<= not WX1129;
	WX1135<= not WX1005;
	WX1137<= not WX1136;
	WX1142<= not WX1005;
	WX1144<= not WX1143;
	WX1149<= not WX1005;
	WX1151<= not WX1150;
	WX1156<= not WX1005;
	WX1158<= not WX1157;
	WX1163<= not WX1005;
	WX1165<= not WX1164;
	WX1170<= not WX1005;
	WX1172<= not WX1171;
	WX1177<= not WX1005;
	WX1179<= not WX1178;
	WX1184<= not WX1005;
	WX1186<= not WX1185;
	WX1191<= not WX1005;
	WX1193<= not WX1192;
	WX1198<= not WX1005;
	WX1200<= not WX1199;
	WX1205<= not WX1005;
	WX1207<= not WX1206;
	WX1212<= not WX1005;
	WX1214<= not WX1213;
	WX1219<= not WX1005;
	WX1221<= not WX1220;
	WX1226<= not WX1005;
	WX1228<= not WX1227;
	WX1230<= not RESET;
	WX1263<= not WX1230;
	WX1330<= not WX2296;
	WX1334<= not WX2297;
	WX1338<= not WX2297;
	WX1340<= not WX1331;
	WX1341<= not WX1340;
	WX1344<= not WX2296;
	WX1348<= not WX2297;
	WX1352<= not WX2297;
	WX1354<= not WX1345;
	WX1355<= not WX1354;
	WX1358<= not WX2296;
	WX1362<= not WX2297;
	WX1366<= not WX2297;
	WX1368<= not WX1359;
	WX1369<= not WX1368;
	WX1372<= not WX2296;
	WX1376<= not WX2297;
	WX1380<= not WX2297;
	WX1382<= not WX1373;
	WX1383<= not WX1382;
	WX1386<= not WX2296;
	WX1390<= not WX2297;
	WX1394<= not WX2297;
	WX1396<= not WX1387;
	WX1397<= not WX1396;
	WX1400<= not WX2296;
	WX1404<= not WX2297;
	WX1408<= not WX2297;
	WX1410<= not WX1401;
	WX1411<= not WX1410;
	WX1414<= not WX2296;
	WX1418<= not WX2297;
	WX1422<= not WX2297;
	WX1424<= not WX1415;
	WX1425<= not WX1424;
	WX1428<= not WX2296;
	WX1432<= not WX2297;
	WX1436<= not WX2297;
	WX1438<= not WX1429;
	WX1439<= not WX1438;
	WX1442<= not WX2296;
	WX1446<= not WX2297;
	WX1450<= not WX2297;
	WX1452<= not WX1443;
	WX1453<= not WX1452;
	WX1456<= not WX2296;
	WX1460<= not WX2297;
	WX1464<= not WX2297;
	WX1466<= not WX1457;
	WX1467<= not WX1466;
	WX1470<= not WX2296;
	WX1474<= not WX2297;
	WX1478<= not WX2297;
	WX1480<= not WX1471;
	WX1481<= not WX1480;
	WX1484<= not WX2296;
	WX1488<= not WX2297;
	WX1492<= not WX2297;
	WX1494<= not WX1485;
	WX1495<= not WX1494;
	WX1498<= not WX2296;
	WX1502<= not WX2297;
	WX1506<= not WX2297;
	WX1508<= not WX1499;
	WX1509<= not WX1508;
	WX1512<= not WX2296;
	WX1516<= not WX2297;
	WX1520<= not WX2297;
	WX1522<= not WX1513;
	WX1523<= not WX1522;
	WX1526<= not WX2296;
	WX1530<= not WX2297;
	WX1534<= not WX2297;
	WX1536<= not WX1527;
	WX1537<= not WX1536;
	WX1540<= not WX2296;
	WX1544<= not WX2297;
	WX1548<= not WX2297;
	WX1550<= not WX1541;
	WX1551<= not WX1550;
	WX1554<= not WX2296;
	WX1558<= not WX2297;
	WX1562<= not WX2297;
	WX1564<= not WX1555;
	WX1565<= not WX1564;
	WX1568<= not WX2296;
	WX1572<= not WX2297;
	WX1576<= not WX2297;
	WX1578<= not WX1569;
	WX1579<= not WX1578;
	WX1582<= not WX2296;
	WX1586<= not WX2297;
	WX1590<= not WX2297;
	WX1592<= not WX1583;
	WX1593<= not WX1592;
	WX1596<= not WX2296;
	WX1600<= not WX2297;
	WX1604<= not WX2297;
	WX1606<= not WX1597;
	WX1607<= not WX1606;
	WX1610<= not WX2296;
	WX1614<= not WX2297;
	WX1618<= not WX2297;
	WX1620<= not WX1611;
	WX1621<= not WX1620;
	WX1624<= not WX2296;
	WX1628<= not WX2297;
	WX1632<= not WX2297;
	WX1634<= not WX1625;
	WX1635<= not WX1634;
	WX1638<= not WX2296;
	WX1642<= not WX2297;
	WX1646<= not WX2297;
	WX1648<= not WX1639;
	WX1649<= not WX1648;
	WX1652<= not WX2296;
	WX1656<= not WX2297;
	WX1660<= not WX2297;
	WX1662<= not WX1653;
	WX1663<= not WX1662;
	WX1666<= not WX2296;
	WX1670<= not WX2297;
	WX1674<= not WX2297;
	WX1676<= not WX1667;
	WX1677<= not WX1676;
	WX1680<= not WX2296;
	WX1684<= not WX2297;
	WX1688<= not WX2297;
	WX1690<= not WX1681;
	WX1691<= not WX1690;
	WX1694<= not WX2296;
	WX1698<= not WX2297;
	WX1702<= not WX2297;
	WX1704<= not WX1695;
	WX1705<= not WX1704;
	WX1708<= not WX2296;
	WX1712<= not WX2297;
	WX1716<= not WX2297;
	WX1718<= not WX1709;
	WX1719<= not WX1718;
	WX1722<= not WX2296;
	WX1726<= not WX2297;
	WX1730<= not WX2297;
	WX1732<= not WX1723;
	WX1733<= not WX1732;
	WX1736<= not WX2296;
	WX1740<= not WX2297;
	WX1744<= not WX2297;
	WX1746<= not WX1737;
	WX1747<= not WX1746;
	WX1750<= not WX2296;
	WX1754<= not WX2297;
	WX1758<= not WX2297;
	WX1760<= not WX1751;
	WX1761<= not WX1760;
	WX1764<= not WX2296;
	WX1768<= not WX2297;
	WX1772<= not WX2297;
	WX1774<= not WX1765;
	WX1775<= not WX1774;
	WX1776<= not WX1778;
	WX1841<= not WX2258;
	WX1842<= not WX2260;
	WX1843<= not WX2262;
	WX1844<= not WX2264;
	WX1845<= not WX2266;
	WX1846<= not WX2268;
	WX1847<= not WX2270;
	WX1848<= not WX2272;
	WX1849<= not WX2274;
	WX1850<= not WX2276;
	WX1851<= not WX2278;
	WX1852<= not WX2280;
	WX1853<= not WX2282;
	WX1854<= not WX2284;
	WX1855<= not WX2286;
	WX1856<= not WX2288;
	WX1857<= not WX2226;
	WX1858<= not WX2228;
	WX1859<= not WX2230;
	WX1860<= not WX2232;
	WX1861<= not WX2234;
	WX1862<= not WX2236;
	WX1863<= not WX2238;
	WX1864<= not WX2240;
	WX1865<= not WX2242;
	WX1866<= not WX2244;
	WX1867<= not WX2246;
	WX1868<= not WX2248;
	WX1869<= not WX2250;
	WX1870<= not WX2252;
	WX1871<= not WX2254;
	WX1872<= not WX2256;
	WX1873<= not WX1841;
	WX1874<= not WX1842;
	WX1875<= not WX1843;
	WX1876<= not WX1844;
	WX1877<= not WX1845;
	WX1878<= not WX1846;
	WX1879<= not WX1847;
	WX1880<= not WX1848;
	WX1881<= not WX1849;
	WX1882<= not WX1850;
	WX1883<= not WX1851;
	WX1884<= not WX1852;
	WX1885<= not WX1853;
	WX1886<= not WX1854;
	WX1887<= not WX1855;
	WX1888<= not WX1856;
	WX1889<= not WX1857;
	WX1890<= not WX1858;
	WX1891<= not WX1859;
	WX1892<= not WX1860;
	WX1893<= not WX1861;
	WX1894<= not WX1862;
	WX1895<= not WX1863;
	WX1896<= not WX1864;
	WX1897<= not WX1865;
	WX1898<= not WX1866;
	WX1899<= not WX1867;
	WX1900<= not WX1868;
	WX1901<= not WX1869;
	WX1902<= not WX1870;
	WX1903<= not WX1871;
	WX1904<= not WX1872;
	WX1905<= not WX2130;
	WX1906<= not WX2132;
	WX1907<= not WX2134;
	WX1908<= not WX2136;
	WX1909<= not WX2138;
	WX1910<= not WX2140;
	WX1911<= not WX2142;
	WX1912<= not WX2144;
	WX1913<= not WX2146;
	WX1914<= not WX2148;
	WX1915<= not WX2150;
	WX1916<= not WX2152;
	WX1917<= not WX2154;
	WX1918<= not WX2156;
	WX1919<= not WX2158;
	WX1920<= not WX2160;
	WX1921<= not WX2162;
	WX1922<= not WX2164;
	WX1923<= not WX2166;
	WX1924<= not WX2168;
	WX1925<= not WX2170;
	WX1926<= not WX2172;
	WX1927<= not WX2174;
	WX1928<= not WX2176;
	WX1929<= not WX2178;
	WX1930<= not WX2180;
	WX1931<= not WX2182;
	WX1932<= not WX2184;
	WX1933<= not WX2186;
	WX1934<= not WX2188;
	WX1935<= not WX2190;
	WX1936<= not WX2192;
	WX2225<= not WX2209;
	WX2226<= not WX2225;
	WX2227<= not WX2210;
	WX2228<= not WX2227;
	WX2229<= not WX2211;
	WX2230<= not WX2229;
	WX2231<= not WX2212;
	WX2232<= not WX2231;
	WX2233<= not WX2213;
	WX2234<= not WX2233;
	WX2235<= not WX2214;
	WX2236<= not WX2235;
	WX2237<= not WX2215;
	WX2238<= not WX2237;
	WX2239<= not WX2216;
	WX2240<= not WX2239;
	WX2241<= not WX2217;
	WX2242<= not WX2241;
	WX2243<= not WX2218;
	WX2244<= not WX2243;
	WX2245<= not WX2219;
	WX2246<= not WX2245;
	WX2247<= not WX2220;
	WX2248<= not WX2247;
	WX2249<= not WX2221;
	WX2250<= not WX2249;
	WX2251<= not WX2222;
	WX2252<= not WX2251;
	WX2253<= not WX2223;
	WX2254<= not WX2253;
	WX2255<= not WX2224;
	WX2256<= not WX2255;
	WX2257<= not WX2193;
	WX2258<= not WX2257;
	WX2259<= not WX2194;
	WX2260<= not WX2259;
	WX2261<= not WX2195;
	WX2262<= not WX2261;
	WX2263<= not WX2196;
	WX2264<= not WX2263;
	WX2265<= not WX2197;
	WX2266<= not WX2265;
	WX2267<= not WX2198;
	WX2268<= not WX2267;
	WX2269<= not WX2199;
	WX2270<= not WX2269;
	WX2271<= not WX2200;
	WX2272<= not WX2271;
	WX2273<= not WX2201;
	WX2274<= not WX2273;
	WX2275<= not WX2202;
	WX2276<= not WX2275;
	WX2277<= not WX2203;
	WX2278<= not WX2277;
	WX2279<= not WX2204;
	WX2280<= not WX2279;
	WX2281<= not WX2205;
	WX2282<= not WX2281;
	WX2283<= not WX2206;
	WX2284<= not WX2283;
	WX2285<= not WX2207;
	WX2286<= not WX2285;
	WX2287<= not WX2208;
	WX2288<= not WX2287;
	WX2289<= not TM0;
	WX2290<= not TM0;
	WX2291<= not TM0;
	WX2292<= not TM1;
	WX2293<= not TM1;
	WX2294<= not WX2293;
	WX2295<= not WX2291;
	WX2296<= not WX2292;
	WX2297<= not WX2290;
	WX2298<= not WX2289;
	WX2302<= not WX2298;
	WX2304<= not WX2303;
	WX2305<= not WX2304;
	WX2309<= not WX2298;
	WX2311<= not WX2310;
	WX2312<= not WX2311;
	WX2316<= not WX2298;
	WX2318<= not WX2317;
	WX2319<= not WX2318;
	WX2323<= not WX2298;
	WX2325<= not WX2324;
	WX2326<= not WX2325;
	WX2330<= not WX2298;
	WX2332<= not WX2331;
	WX2333<= not WX2332;
	WX2337<= not WX2298;
	WX2339<= not WX2338;
	WX2340<= not WX2339;
	WX2344<= not WX2298;
	WX2346<= not WX2345;
	WX2347<= not WX2346;
	WX2351<= not WX2298;
	WX2353<= not WX2352;
	WX2354<= not WX2353;
	WX2358<= not WX2298;
	WX2360<= not WX2359;
	WX2361<= not WX2360;
	WX2365<= not WX2298;
	WX2367<= not WX2366;
	WX2368<= not WX2367;
	WX2372<= not WX2298;
	WX2374<= not WX2373;
	WX2375<= not WX2374;
	WX2379<= not WX2298;
	WX2381<= not WX2380;
	WX2382<= not WX2381;
	WX2386<= not WX2298;
	WX2388<= not WX2387;
	WX2389<= not WX2388;
	WX2393<= not WX2298;
	WX2395<= not WX2394;
	WX2396<= not WX2395;
	WX2400<= not WX2298;
	WX2402<= not WX2401;
	WX2403<= not WX2402;
	WX2407<= not WX2298;
	WX2409<= not WX2408;
	WX2410<= not WX2409;
	WX2414<= not WX2298;
	WX2416<= not WX2415;
	WX2417<= not WX2416;
	WX2421<= not WX2298;
	WX2423<= not WX2422;
	WX2424<= not WX2423;
	WX2428<= not WX2298;
	WX2430<= not WX2429;
	WX2431<= not WX2430;
	WX2435<= not WX2298;
	WX2437<= not WX2436;
	WX2438<= not WX2437;
	WX2442<= not WX2298;
	WX2444<= not WX2443;
	WX2445<= not WX2444;
	WX2449<= not WX2298;
	WX2451<= not WX2450;
	WX2452<= not WX2451;
	WX2456<= not WX2298;
	WX2458<= not WX2457;
	WX2459<= not WX2458;
	WX2463<= not WX2298;
	WX2465<= not WX2464;
	WX2466<= not WX2465;
	WX2470<= not WX2298;
	WX2472<= not WX2471;
	WX2473<= not WX2472;
	WX2477<= not WX2298;
	WX2479<= not WX2478;
	WX2480<= not WX2479;
	WX2484<= not WX2298;
	WX2486<= not WX2485;
	WX2487<= not WX2486;
	WX2491<= not WX2298;
	WX2493<= not WX2492;
	WX2494<= not WX2493;
	WX2498<= not WX2298;
	WX2500<= not WX2499;
	WX2501<= not WX2500;
	WX2505<= not WX2298;
	WX2507<= not WX2506;
	WX2508<= not WX2507;
	WX2512<= not WX2298;
	WX2514<= not WX2513;
	WX2515<= not WX2514;
	WX2519<= not WX2298;
	WX2521<= not WX2520;
	WX2522<= not WX2521;
	WX2523<= not RESET;
	WX2556<= not WX2523;
	WX2623<= not WX3589;
	WX2627<= not WX3590;
	WX2631<= not WX3590;
	WX2633<= not WX2624;
	WX2634<= not WX2633;
	WX2637<= not WX3589;
	WX2641<= not WX3590;
	WX2645<= not WX3590;
	WX2647<= not WX2638;
	WX2648<= not WX2647;
	WX2651<= not WX3589;
	WX2655<= not WX3590;
	WX2659<= not WX3590;
	WX2661<= not WX2652;
	WX2662<= not WX2661;
	WX2665<= not WX3589;
	WX2669<= not WX3590;
	WX2673<= not WX3590;
	WX2675<= not WX2666;
	WX2676<= not WX2675;
	WX2679<= not WX3589;
	WX2683<= not WX3590;
	WX2687<= not WX3590;
	WX2689<= not WX2680;
	WX2690<= not WX2689;
	WX2693<= not WX3589;
	WX2697<= not WX3590;
	WX2701<= not WX3590;
	WX2703<= not WX2694;
	WX2704<= not WX2703;
	WX2707<= not WX3589;
	WX2711<= not WX3590;
	WX2715<= not WX3590;
	WX2717<= not WX2708;
	WX2718<= not WX2717;
	WX2721<= not WX3589;
	WX2725<= not WX3590;
	WX2729<= not WX3590;
	WX2731<= not WX2722;
	WX2732<= not WX2731;
	WX2735<= not WX3589;
	WX2739<= not WX3590;
	WX2743<= not WX3590;
	WX2745<= not WX2736;
	WX2746<= not WX2745;
	WX2749<= not WX3589;
	WX2753<= not WX3590;
	WX2757<= not WX3590;
	WX2759<= not WX2750;
	WX2760<= not WX2759;
	WX2763<= not WX3589;
	WX2767<= not WX3590;
	WX2771<= not WX3590;
	WX2773<= not WX2764;
	WX2774<= not WX2773;
	WX2777<= not WX3589;
	WX2781<= not WX3590;
	WX2785<= not WX3590;
	WX2787<= not WX2778;
	WX2788<= not WX2787;
	WX2791<= not WX3589;
	WX2795<= not WX3590;
	WX2799<= not WX3590;
	WX2801<= not WX2792;
	WX2802<= not WX2801;
	WX2805<= not WX3589;
	WX2809<= not WX3590;
	WX2813<= not WX3590;
	WX2815<= not WX2806;
	WX2816<= not WX2815;
	WX2819<= not WX3589;
	WX2823<= not WX3590;
	WX2827<= not WX3590;
	WX2829<= not WX2820;
	WX2830<= not WX2829;
	WX2833<= not WX3589;
	WX2837<= not WX3590;
	WX2841<= not WX3590;
	WX2843<= not WX2834;
	WX2844<= not WX2843;
	WX2847<= not WX3589;
	WX2851<= not WX3590;
	WX2855<= not WX3590;
	WX2857<= not WX2848;
	WX2858<= not WX2857;
	WX2861<= not WX3589;
	WX2865<= not WX3590;
	WX2869<= not WX3590;
	WX2871<= not WX2862;
	WX2872<= not WX2871;
	WX2875<= not WX3589;
	WX2879<= not WX3590;
	WX2883<= not WX3590;
	WX2885<= not WX2876;
	WX2886<= not WX2885;
	WX2889<= not WX3589;
	WX2893<= not WX3590;
	WX2897<= not WX3590;
	WX2899<= not WX2890;
	WX2900<= not WX2899;
	WX2903<= not WX3589;
	WX2907<= not WX3590;
	WX2911<= not WX3590;
	WX2913<= not WX2904;
	WX2914<= not WX2913;
	WX2917<= not WX3589;
	WX2921<= not WX3590;
	WX2925<= not WX3590;
	WX2927<= not WX2918;
	WX2928<= not WX2927;
	WX2931<= not WX3589;
	WX2935<= not WX3590;
	WX2939<= not WX3590;
	WX2941<= not WX2932;
	WX2942<= not WX2941;
	WX2945<= not WX3589;
	WX2949<= not WX3590;
	WX2953<= not WX3590;
	WX2955<= not WX2946;
	WX2956<= not WX2955;
	WX2959<= not WX3589;
	WX2963<= not WX3590;
	WX2967<= not WX3590;
	WX2969<= not WX2960;
	WX2970<= not WX2969;
	WX2973<= not WX3589;
	WX2977<= not WX3590;
	WX2981<= not WX3590;
	WX2983<= not WX2974;
	WX2984<= not WX2983;
	WX2987<= not WX3589;
	WX2991<= not WX3590;
	WX2995<= not WX3590;
	WX2997<= not WX2988;
	WX2998<= not WX2997;
	WX3001<= not WX3589;
	WX3005<= not WX3590;
	WX3009<= not WX3590;
	WX3011<= not WX3002;
	WX3012<= not WX3011;
	WX3015<= not WX3589;
	WX3019<= not WX3590;
	WX3023<= not WX3590;
	WX3025<= not WX3016;
	WX3026<= not WX3025;
	WX3029<= not WX3589;
	WX3033<= not WX3590;
	WX3037<= not WX3590;
	WX3039<= not WX3030;
	WX3040<= not WX3039;
	WX3043<= not WX3589;
	WX3047<= not WX3590;
	WX3051<= not WX3590;
	WX3053<= not WX3044;
	WX3054<= not WX3053;
	WX3057<= not WX3589;
	WX3061<= not WX3590;
	WX3065<= not WX3590;
	WX3067<= not WX3058;
	WX3068<= not WX3067;
	WX3069<= not WX3071;
	WX3134<= not WX3551;
	WX3135<= not WX3553;
	WX3136<= not WX3555;
	WX3137<= not WX3557;
	WX3138<= not WX3559;
	WX3139<= not WX3561;
	WX3140<= not WX3563;
	WX3141<= not WX3565;
	WX3142<= not WX3567;
	WX3143<= not WX3569;
	WX3144<= not WX3571;
	WX3145<= not WX3573;
	WX3146<= not WX3575;
	WX3147<= not WX3577;
	WX3148<= not WX3579;
	WX3149<= not WX3581;
	WX3150<= not WX3519;
	WX3151<= not WX3521;
	WX3152<= not WX3523;
	WX3153<= not WX3525;
	WX3154<= not WX3527;
	WX3155<= not WX3529;
	WX3156<= not WX3531;
	WX3157<= not WX3533;
	WX3158<= not WX3535;
	WX3159<= not WX3537;
	WX3160<= not WX3539;
	WX3161<= not WX3541;
	WX3162<= not WX3543;
	WX3163<= not WX3545;
	WX3164<= not WX3547;
	WX3165<= not WX3549;
	WX3166<= not WX3134;
	WX3167<= not WX3135;
	WX3168<= not WX3136;
	WX3169<= not WX3137;
	WX3170<= not WX3138;
	WX3171<= not WX3139;
	WX3172<= not WX3140;
	WX3173<= not WX3141;
	WX3174<= not WX3142;
	WX3175<= not WX3143;
	WX3176<= not WX3144;
	WX3177<= not WX3145;
	WX3178<= not WX3146;
	WX3179<= not WX3147;
	WX3180<= not WX3148;
	WX3181<= not WX3149;
	WX3182<= not WX3150;
	WX3183<= not WX3151;
	WX3184<= not WX3152;
	WX3185<= not WX3153;
	WX3186<= not WX3154;
	WX3187<= not WX3155;
	WX3188<= not WX3156;
	WX3189<= not WX3157;
	WX3190<= not WX3158;
	WX3191<= not WX3159;
	WX3192<= not WX3160;
	WX3193<= not WX3161;
	WX3194<= not WX3162;
	WX3195<= not WX3163;
	WX3196<= not WX3164;
	WX3197<= not WX3165;
	WX3198<= not WX3423;
	WX3199<= not WX3425;
	WX3200<= not WX3427;
	WX3201<= not WX3429;
	WX3202<= not WX3431;
	WX3203<= not WX3433;
	WX3204<= not WX3435;
	WX3205<= not WX3437;
	WX3206<= not WX3439;
	WX3207<= not WX3441;
	WX3208<= not WX3443;
	WX3209<= not WX3445;
	WX3210<= not WX3447;
	WX3211<= not WX3449;
	WX3212<= not WX3451;
	WX3213<= not WX3453;
	WX3214<= not WX3455;
	WX3215<= not WX3457;
	WX3216<= not WX3459;
	WX3217<= not WX3461;
	WX3218<= not WX3463;
	WX3219<= not WX3465;
	WX3220<= not WX3467;
	WX3221<= not WX3469;
	WX3222<= not WX3471;
	WX3223<= not WX3473;
	WX3224<= not WX3475;
	WX3225<= not WX3477;
	WX3226<= not WX3479;
	WX3227<= not WX3481;
	WX3228<= not WX3483;
	WX3229<= not WX3485;
	WX3518<= not WX3502;
	WX3519<= not WX3518;
	WX3520<= not WX3503;
	WX3521<= not WX3520;
	WX3522<= not WX3504;
	WX3523<= not WX3522;
	WX3524<= not WX3505;
	WX3525<= not WX3524;
	WX3526<= not WX3506;
	WX3527<= not WX3526;
	WX3528<= not WX3507;
	WX3529<= not WX3528;
	WX3530<= not WX3508;
	WX3531<= not WX3530;
	WX3532<= not WX3509;
	WX3533<= not WX3532;
	WX3534<= not WX3510;
	WX3535<= not WX3534;
	WX3536<= not WX3511;
	WX3537<= not WX3536;
	WX3538<= not WX3512;
	WX3539<= not WX3538;
	WX3540<= not WX3513;
	WX3541<= not WX3540;
	WX3542<= not WX3514;
	WX3543<= not WX3542;
	WX3544<= not WX3515;
	WX3545<= not WX3544;
	WX3546<= not WX3516;
	WX3547<= not WX3546;
	WX3548<= not WX3517;
	WX3549<= not WX3548;
	WX3550<= not WX3486;
	WX3551<= not WX3550;
	WX3552<= not WX3487;
	WX3553<= not WX3552;
	WX3554<= not WX3488;
	WX3555<= not WX3554;
	WX3556<= not WX3489;
	WX3557<= not WX3556;
	WX3558<= not WX3490;
	WX3559<= not WX3558;
	WX3560<= not WX3491;
	WX3561<= not WX3560;
	WX3562<= not WX3492;
	WX3563<= not WX3562;
	WX3564<= not WX3493;
	WX3565<= not WX3564;
	WX3566<= not WX3494;
	WX3567<= not WX3566;
	WX3568<= not WX3495;
	WX3569<= not WX3568;
	WX3570<= not WX3496;
	WX3571<= not WX3570;
	WX3572<= not WX3497;
	WX3573<= not WX3572;
	WX3574<= not WX3498;
	WX3575<= not WX3574;
	WX3576<= not WX3499;
	WX3577<= not WX3576;
	WX3578<= not WX3500;
	WX3579<= not WX3578;
	WX3580<= not WX3501;
	WX3581<= not WX3580;
	WX3582<= not TM0;
	WX3583<= not TM0;
	WX3584<= not TM0;
	WX3585<= not TM1;
	WX3586<= not TM1;
	WX3587<= not WX3586;
	WX3588<= not WX3584;
	WX3589<= not WX3585;
	WX3590<= not WX3583;
	WX3591<= not WX3582;
	WX3595<= not WX3591;
	WX3597<= not WX3596;
	WX3598<= not WX3597;
	WX3602<= not WX3591;
	WX3604<= not WX3603;
	WX3605<= not WX3604;
	WX3609<= not WX3591;
	WX3611<= not WX3610;
	WX3612<= not WX3611;
	WX3616<= not WX3591;
	WX3618<= not WX3617;
	WX3619<= not WX3618;
	WX3623<= not WX3591;
	WX3625<= not WX3624;
	WX3626<= not WX3625;
	WX3630<= not WX3591;
	WX3632<= not WX3631;
	WX3633<= not WX3632;
	WX3637<= not WX3591;
	WX3639<= not WX3638;
	WX3640<= not WX3639;
	WX3644<= not WX3591;
	WX3646<= not WX3645;
	WX3647<= not WX3646;
	WX3651<= not WX3591;
	WX3653<= not WX3652;
	WX3654<= not WX3653;
	WX3658<= not WX3591;
	WX3660<= not WX3659;
	WX3661<= not WX3660;
	WX3665<= not WX3591;
	WX3667<= not WX3666;
	WX3668<= not WX3667;
	WX3672<= not WX3591;
	WX3674<= not WX3673;
	WX3675<= not WX3674;
	WX3679<= not WX3591;
	WX3681<= not WX3680;
	WX3682<= not WX3681;
	WX3686<= not WX3591;
	WX3688<= not WX3687;
	WX3689<= not WX3688;
	WX3693<= not WX3591;
	WX3695<= not WX3694;
	WX3696<= not WX3695;
	WX3700<= not WX3591;
	WX3702<= not WX3701;
	WX3703<= not WX3702;
	WX3707<= not WX3591;
	WX3709<= not WX3708;
	WX3710<= not WX3709;
	WX3714<= not WX3591;
	WX3716<= not WX3715;
	WX3717<= not WX3716;
	WX3721<= not WX3591;
	WX3723<= not WX3722;
	WX3724<= not WX3723;
	WX3728<= not WX3591;
	WX3730<= not WX3729;
	WX3731<= not WX3730;
	WX3735<= not WX3591;
	WX3737<= not WX3736;
	WX3738<= not WX3737;
	WX3742<= not WX3591;
	WX3744<= not WX3743;
	WX3745<= not WX3744;
	WX3749<= not WX3591;
	WX3751<= not WX3750;
	WX3752<= not WX3751;
	WX3756<= not WX3591;
	WX3758<= not WX3757;
	WX3759<= not WX3758;
	WX3763<= not WX3591;
	WX3765<= not WX3764;
	WX3766<= not WX3765;
	WX3770<= not WX3591;
	WX3772<= not WX3771;
	WX3773<= not WX3772;
	WX3777<= not WX3591;
	WX3779<= not WX3778;
	WX3780<= not WX3779;
	WX3784<= not WX3591;
	WX3786<= not WX3785;
	WX3787<= not WX3786;
	WX3791<= not WX3591;
	WX3793<= not WX3792;
	WX3794<= not WX3793;
	WX3798<= not WX3591;
	WX3800<= not WX3799;
	WX3801<= not WX3800;
	WX3805<= not WX3591;
	WX3807<= not WX3806;
	WX3808<= not WX3807;
	WX3812<= not WX3591;
	WX3814<= not WX3813;
	WX3815<= not WX3814;
	WX3816<= not RESET;
	WX3849<= not WX3816;
	WX3916<= not WX4882;
	WX3920<= not WX4883;
	WX3924<= not WX4883;
	WX3926<= not WX3917;
	WX3927<= not WX3926;
	WX3930<= not WX4882;
	WX3934<= not WX4883;
	WX3938<= not WX4883;
	WX3940<= not WX3931;
	WX3941<= not WX3940;
	WX3944<= not WX4882;
	WX3948<= not WX4883;
	WX3952<= not WX4883;
	WX3954<= not WX3945;
	WX3955<= not WX3954;
	WX3958<= not WX4882;
	WX3962<= not WX4883;
	WX3966<= not WX4883;
	WX3968<= not WX3959;
	WX3969<= not WX3968;
	WX3972<= not WX4882;
	WX3976<= not WX4883;
	WX3980<= not WX4883;
	WX3982<= not WX3973;
	WX3983<= not WX3982;
	WX3986<= not WX4882;
	WX3990<= not WX4883;
	WX3994<= not WX4883;
	WX3996<= not WX3987;
	WX3997<= not WX3996;
	WX4000<= not WX4882;
	WX4004<= not WX4883;
	WX4008<= not WX4883;
	WX4010<= not WX4001;
	WX4011<= not WX4010;
	WX4014<= not WX4882;
	WX4018<= not WX4883;
	WX4022<= not WX4883;
	WX4024<= not WX4015;
	WX4025<= not WX4024;
	WX4028<= not WX4882;
	WX4032<= not WX4883;
	WX4036<= not WX4883;
	WX4038<= not WX4029;
	WX4039<= not WX4038;
	WX4042<= not WX4882;
	WX4046<= not WX4883;
	WX4050<= not WX4883;
	WX4052<= not WX4043;
	WX4053<= not WX4052;
	WX4056<= not WX4882;
	WX4060<= not WX4883;
	WX4064<= not WX4883;
	WX4066<= not WX4057;
	WX4067<= not WX4066;
	WX4070<= not WX4882;
	WX4074<= not WX4883;
	WX4078<= not WX4883;
	WX4080<= not WX4071;
	WX4081<= not WX4080;
	WX4084<= not WX4882;
	WX4088<= not WX4883;
	WX4092<= not WX4883;
	WX4094<= not WX4085;
	WX4095<= not WX4094;
	WX4098<= not WX4882;
	WX4102<= not WX4883;
	WX4106<= not WX4883;
	WX4108<= not WX4099;
	WX4109<= not WX4108;
	WX4112<= not WX4882;
	WX4116<= not WX4883;
	WX4120<= not WX4883;
	WX4122<= not WX4113;
	WX4123<= not WX4122;
	WX4126<= not WX4882;
	WX4130<= not WX4883;
	WX4134<= not WX4883;
	WX4136<= not WX4127;
	WX4137<= not WX4136;
	WX4140<= not WX4882;
	WX4144<= not WX4883;
	WX4148<= not WX4883;
	WX4150<= not WX4141;
	WX4151<= not WX4150;
	WX4154<= not WX4882;
	WX4158<= not WX4883;
	WX4162<= not WX4883;
	WX4164<= not WX4155;
	WX4165<= not WX4164;
	WX4168<= not WX4882;
	WX4172<= not WX4883;
	WX4176<= not WX4883;
	WX4178<= not WX4169;
	WX4179<= not WX4178;
	WX4182<= not WX4882;
	WX4186<= not WX4883;
	WX4190<= not WX4883;
	WX4192<= not WX4183;
	WX4193<= not WX4192;
	WX4196<= not WX4882;
	WX4200<= not WX4883;
	WX4204<= not WX4883;
	WX4206<= not WX4197;
	WX4207<= not WX4206;
	WX4210<= not WX4882;
	WX4214<= not WX4883;
	WX4218<= not WX4883;
	WX4220<= not WX4211;
	WX4221<= not WX4220;
	WX4224<= not WX4882;
	WX4228<= not WX4883;
	WX4232<= not WX4883;
	WX4234<= not WX4225;
	WX4235<= not WX4234;
	WX4238<= not WX4882;
	WX4242<= not WX4883;
	WX4246<= not WX4883;
	WX4248<= not WX4239;
	WX4249<= not WX4248;
	WX4252<= not WX4882;
	WX4256<= not WX4883;
	WX4260<= not WX4883;
	WX4262<= not WX4253;
	WX4263<= not WX4262;
	WX4266<= not WX4882;
	WX4270<= not WX4883;
	WX4274<= not WX4883;
	WX4276<= not WX4267;
	WX4277<= not WX4276;
	WX4280<= not WX4882;
	WX4284<= not WX4883;
	WX4288<= not WX4883;
	WX4290<= not WX4281;
	WX4291<= not WX4290;
	WX4294<= not WX4882;
	WX4298<= not WX4883;
	WX4302<= not WX4883;
	WX4304<= not WX4295;
	WX4305<= not WX4304;
	WX4308<= not WX4882;
	WX4312<= not WX4883;
	WX4316<= not WX4883;
	WX4318<= not WX4309;
	WX4319<= not WX4318;
	WX4322<= not WX4882;
	WX4326<= not WX4883;
	WX4330<= not WX4883;
	WX4332<= not WX4323;
	WX4333<= not WX4332;
	WX4336<= not WX4882;
	WX4340<= not WX4883;
	WX4344<= not WX4883;
	WX4346<= not WX4337;
	WX4347<= not WX4346;
	WX4350<= not WX4882;
	WX4354<= not WX4883;
	WX4358<= not WX4883;
	WX4360<= not WX4351;
	WX4361<= not WX4360;
	WX4362<= not WX4364;
	WX4427<= not WX4844;
	WX4428<= not WX4846;
	WX4429<= not WX4848;
	WX4430<= not WX4850;
	WX4431<= not WX4852;
	WX4432<= not WX4854;
	WX4433<= not WX4856;
	WX4434<= not WX4858;
	WX4435<= not WX4860;
	WX4436<= not WX4862;
	WX4437<= not WX4864;
	WX4438<= not WX4866;
	WX4439<= not WX4868;
	WX4440<= not WX4870;
	WX4441<= not WX4872;
	WX4442<= not WX4874;
	WX4443<= not WX4812;
	WX4444<= not WX4814;
	WX4445<= not WX4816;
	WX4446<= not WX4818;
	WX4447<= not WX4820;
	WX4448<= not WX4822;
	WX4449<= not WX4824;
	WX4450<= not WX4826;
	WX4451<= not WX4828;
	WX4452<= not WX4830;
	WX4453<= not WX4832;
	WX4454<= not WX4834;
	WX4455<= not WX4836;
	WX4456<= not WX4838;
	WX4457<= not WX4840;
	WX4458<= not WX4842;
	WX4459<= not WX4427;
	WX4460<= not WX4428;
	WX4461<= not WX4429;
	WX4462<= not WX4430;
	WX4463<= not WX4431;
	WX4464<= not WX4432;
	WX4465<= not WX4433;
	WX4466<= not WX4434;
	WX4467<= not WX4435;
	WX4468<= not WX4436;
	WX4469<= not WX4437;
	WX4470<= not WX4438;
	WX4471<= not WX4439;
	WX4472<= not WX4440;
	WX4473<= not WX4441;
	WX4474<= not WX4442;
	WX4475<= not WX4443;
	WX4476<= not WX4444;
	WX4477<= not WX4445;
	WX4478<= not WX4446;
	WX4479<= not WX4447;
	WX4480<= not WX4448;
	WX4481<= not WX4449;
	WX4482<= not WX4450;
	WX4483<= not WX4451;
	WX4484<= not WX4452;
	WX4485<= not WX4453;
	WX4486<= not WX4454;
	WX4487<= not WX4455;
	WX4488<= not WX4456;
	WX4489<= not WX4457;
	WX4490<= not WX4458;
	WX4491<= not WX4716;
	WX4492<= not WX4718;
	WX4493<= not WX4720;
	WX4494<= not WX4722;
	WX4495<= not WX4724;
	WX4496<= not WX4726;
	WX4497<= not WX4728;
	WX4498<= not WX4730;
	WX4499<= not WX4732;
	WX4500<= not WX4734;
	WX4501<= not WX4736;
	WX4502<= not WX4738;
	WX4503<= not WX4740;
	WX4504<= not WX4742;
	WX4505<= not WX4744;
	WX4506<= not WX4746;
	WX4507<= not WX4748;
	WX4508<= not WX4750;
	WX4509<= not WX4752;
	WX4510<= not WX4754;
	WX4511<= not WX4756;
	WX4512<= not WX4758;
	WX4513<= not WX4760;
	WX4514<= not WX4762;
	WX4515<= not WX4764;
	WX4516<= not WX4766;
	WX4517<= not WX4768;
	WX4518<= not WX4770;
	WX4519<= not WX4772;
	WX4520<= not WX4774;
	WX4521<= not WX4776;
	WX4522<= not WX4778;
	WX4811<= not WX4795;
	WX4812<= not WX4811;
	WX4813<= not WX4796;
	WX4814<= not WX4813;
	WX4815<= not WX4797;
	WX4816<= not WX4815;
	WX4817<= not WX4798;
	WX4818<= not WX4817;
	WX4819<= not WX4799;
	WX4820<= not WX4819;
	WX4821<= not WX4800;
	WX4822<= not WX4821;
	WX4823<= not WX4801;
	WX4824<= not WX4823;
	WX4825<= not WX4802;
	WX4826<= not WX4825;
	WX4827<= not WX4803;
	WX4828<= not WX4827;
	WX4829<= not WX4804;
	WX4830<= not WX4829;
	WX4831<= not WX4805;
	WX4832<= not WX4831;
	WX4833<= not WX4806;
	WX4834<= not WX4833;
	WX4835<= not WX4807;
	WX4836<= not WX4835;
	WX4837<= not WX4808;
	WX4838<= not WX4837;
	WX4839<= not WX4809;
	WX4840<= not WX4839;
	WX4841<= not WX4810;
	WX4842<= not WX4841;
	WX4843<= not WX4779;
	WX4844<= not WX4843;
	WX4845<= not WX4780;
	WX4846<= not WX4845;
	WX4847<= not WX4781;
	WX4848<= not WX4847;
	WX4849<= not WX4782;
	WX4850<= not WX4849;
	WX4851<= not WX4783;
	WX4852<= not WX4851;
	WX4853<= not WX4784;
	WX4854<= not WX4853;
	WX4855<= not WX4785;
	WX4856<= not WX4855;
	WX4857<= not WX4786;
	WX4858<= not WX4857;
	WX4859<= not WX4787;
	WX4860<= not WX4859;
	WX4861<= not WX4788;
	WX4862<= not WX4861;
	WX4863<= not WX4789;
	WX4864<= not WX4863;
	WX4865<= not WX4790;
	WX4866<= not WX4865;
	WX4867<= not WX4791;
	WX4868<= not WX4867;
	WX4869<= not WX4792;
	WX4870<= not WX4869;
	WX4871<= not WX4793;
	WX4872<= not WX4871;
	WX4873<= not WX4794;
	WX4874<= not WX4873;
	WX4875<= not TM0;
	WX4876<= not TM0;
	WX4877<= not TM0;
	WX4878<= not TM1;
	WX4879<= not TM1;
	WX4880<= not WX4879;
	WX4881<= not WX4877;
	WX4882<= not WX4878;
	WX4883<= not WX4876;
	WX4884<= not WX4875;
	WX4888<= not WX4884;
	WX4890<= not WX4889;
	WX4891<= not WX4890;
	WX4895<= not WX4884;
	WX4897<= not WX4896;
	WX4898<= not WX4897;
	WX4902<= not WX4884;
	WX4904<= not WX4903;
	WX4905<= not WX4904;
	WX4909<= not WX4884;
	WX4911<= not WX4910;
	WX4912<= not WX4911;
	WX4916<= not WX4884;
	WX4918<= not WX4917;
	WX4919<= not WX4918;
	WX4923<= not WX4884;
	WX4925<= not WX4924;
	WX4926<= not WX4925;
	WX4930<= not WX4884;
	WX4932<= not WX4931;
	WX4933<= not WX4932;
	WX4937<= not WX4884;
	WX4939<= not WX4938;
	WX4940<= not WX4939;
	WX4944<= not WX4884;
	WX4946<= not WX4945;
	WX4947<= not WX4946;
	WX4951<= not WX4884;
	WX4953<= not WX4952;
	WX4954<= not WX4953;
	WX4958<= not WX4884;
	WX4960<= not WX4959;
	WX4961<= not WX4960;
	WX4965<= not WX4884;
	WX4967<= not WX4966;
	WX4968<= not WX4967;
	WX4972<= not WX4884;
	WX4974<= not WX4973;
	WX4975<= not WX4974;
	WX4979<= not WX4884;
	WX4981<= not WX4980;
	WX4982<= not WX4981;
	WX4986<= not WX4884;
	WX4988<= not WX4987;
	WX4989<= not WX4988;
	WX4993<= not WX4884;
	WX4995<= not WX4994;
	WX4996<= not WX4995;
	WX5000<= not WX4884;
	WX5002<= not WX5001;
	WX5003<= not WX5002;
	WX5007<= not WX4884;
	WX5009<= not WX5008;
	WX5010<= not WX5009;
	WX5014<= not WX4884;
	WX5016<= not WX5015;
	WX5017<= not WX5016;
	WX5021<= not WX4884;
	WX5023<= not WX5022;
	WX5024<= not WX5023;
	WX5028<= not WX4884;
	WX5030<= not WX5029;
	WX5031<= not WX5030;
	WX5035<= not WX4884;
	WX5037<= not WX5036;
	WX5038<= not WX5037;
	WX5042<= not WX4884;
	WX5044<= not WX5043;
	WX5045<= not WX5044;
	WX5049<= not WX4884;
	WX5051<= not WX5050;
	WX5052<= not WX5051;
	WX5056<= not WX4884;
	WX5058<= not WX5057;
	WX5059<= not WX5058;
	WX5063<= not WX4884;
	WX5065<= not WX5064;
	WX5066<= not WX5065;
	WX5070<= not WX4884;
	WX5072<= not WX5071;
	WX5073<= not WX5072;
	WX5077<= not WX4884;
	WX5079<= not WX5078;
	WX5080<= not WX5079;
	WX5084<= not WX4884;
	WX5086<= not WX5085;
	WX5087<= not WX5086;
	WX5091<= not WX4884;
	WX5093<= not WX5092;
	WX5094<= not WX5093;
	WX5098<= not WX4884;
	WX5100<= not WX5099;
	WX5101<= not WX5100;
	WX5105<= not WX4884;
	WX5107<= not WX5106;
	WX5108<= not WX5107;
	WX5109<= not RESET;
	WX5142<= not WX5109;
	WX5209<= not WX6175;
	WX5213<= not WX6176;
	WX5217<= not WX6176;
	WX5219<= not WX5210;
	WX5220<= not WX5219;
	WX5223<= not WX6175;
	WX5227<= not WX6176;
	WX5231<= not WX6176;
	WX5233<= not WX5224;
	WX5234<= not WX5233;
	WX5237<= not WX6175;
	WX5241<= not WX6176;
	WX5245<= not WX6176;
	WX5247<= not WX5238;
	WX5248<= not WX5247;
	WX5251<= not WX6175;
	WX5255<= not WX6176;
	WX5259<= not WX6176;
	WX5261<= not WX5252;
	WX5262<= not WX5261;
	WX5265<= not WX6175;
	WX5269<= not WX6176;
	WX5273<= not WX6176;
	WX5275<= not WX5266;
	WX5276<= not WX5275;
	WX5279<= not WX6175;
	WX5283<= not WX6176;
	WX5287<= not WX6176;
	WX5289<= not WX5280;
	WX5290<= not WX5289;
	WX5293<= not WX6175;
	WX5297<= not WX6176;
	WX5301<= not WX6176;
	WX5303<= not WX5294;
	WX5304<= not WX5303;
	WX5307<= not WX6175;
	WX5311<= not WX6176;
	WX5315<= not WX6176;
	WX5317<= not WX5308;
	WX5318<= not WX5317;
	WX5321<= not WX6175;
	WX5325<= not WX6176;
	WX5329<= not WX6176;
	WX5331<= not WX5322;
	WX5332<= not WX5331;
	WX5335<= not WX6175;
	WX5339<= not WX6176;
	WX5343<= not WX6176;
	WX5345<= not WX5336;
	WX5346<= not WX5345;
	WX5349<= not WX6175;
	WX5353<= not WX6176;
	WX5357<= not WX6176;
	WX5359<= not WX5350;
	WX5360<= not WX5359;
	WX5363<= not WX6175;
	WX5367<= not WX6176;
	WX5371<= not WX6176;
	WX5373<= not WX5364;
	WX5374<= not WX5373;
	WX5377<= not WX6175;
	WX5381<= not WX6176;
	WX5385<= not WX6176;
	WX5387<= not WX5378;
	WX5388<= not WX5387;
	WX5391<= not WX6175;
	WX5395<= not WX6176;
	WX5399<= not WX6176;
	WX5401<= not WX5392;
	WX5402<= not WX5401;
	WX5405<= not WX6175;
	WX5409<= not WX6176;
	WX5413<= not WX6176;
	WX5415<= not WX5406;
	WX5416<= not WX5415;
	WX5419<= not WX6175;
	WX5423<= not WX6176;
	WX5427<= not WX6176;
	WX5429<= not WX5420;
	WX5430<= not WX5429;
	WX5433<= not WX6175;
	WX5437<= not WX6176;
	WX5441<= not WX6176;
	WX5443<= not WX5434;
	WX5444<= not WX5443;
	WX5447<= not WX6175;
	WX5451<= not WX6176;
	WX5455<= not WX6176;
	WX5457<= not WX5448;
	WX5458<= not WX5457;
	WX5461<= not WX6175;
	WX5465<= not WX6176;
	WX5469<= not WX6176;
	WX5471<= not WX5462;
	WX5472<= not WX5471;
	WX5475<= not WX6175;
	WX5479<= not WX6176;
	WX5483<= not WX6176;
	WX5485<= not WX5476;
	WX5486<= not WX5485;
	WX5489<= not WX6175;
	WX5493<= not WX6176;
	WX5497<= not WX6176;
	WX5499<= not WX5490;
	WX5500<= not WX5499;
	WX5503<= not WX6175;
	WX5507<= not WX6176;
	WX5511<= not WX6176;
	WX5513<= not WX5504;
	WX5514<= not WX5513;
	WX5517<= not WX6175;
	WX5521<= not WX6176;
	WX5525<= not WX6176;
	WX5527<= not WX5518;
	WX5528<= not WX5527;
	WX5531<= not WX6175;
	WX5535<= not WX6176;
	WX5539<= not WX6176;
	WX5541<= not WX5532;
	WX5542<= not WX5541;
	WX5545<= not WX6175;
	WX5549<= not WX6176;
	WX5553<= not WX6176;
	WX5555<= not WX5546;
	WX5556<= not WX5555;
	WX5559<= not WX6175;
	WX5563<= not WX6176;
	WX5567<= not WX6176;
	WX5569<= not WX5560;
	WX5570<= not WX5569;
	WX5573<= not WX6175;
	WX5577<= not WX6176;
	WX5581<= not WX6176;
	WX5583<= not WX5574;
	WX5584<= not WX5583;
	WX5587<= not WX6175;
	WX5591<= not WX6176;
	WX5595<= not WX6176;
	WX5597<= not WX5588;
	WX5598<= not WX5597;
	WX5601<= not WX6175;
	WX5605<= not WX6176;
	WX5609<= not WX6176;
	WX5611<= not WX5602;
	WX5612<= not WX5611;
	WX5615<= not WX6175;
	WX5619<= not WX6176;
	WX5623<= not WX6176;
	WX5625<= not WX5616;
	WX5626<= not WX5625;
	WX5629<= not WX6175;
	WX5633<= not WX6176;
	WX5637<= not WX6176;
	WX5639<= not WX5630;
	WX5640<= not WX5639;
	WX5643<= not WX6175;
	WX5647<= not WX6176;
	WX5651<= not WX6176;
	WX5653<= not WX5644;
	WX5654<= not WX5653;
	WX5655<= not WX5657;
	WX5720<= not WX6137;
	WX5721<= not WX6139;
	WX5722<= not WX6141;
	WX5723<= not WX6143;
	WX5724<= not WX6145;
	WX5725<= not WX6147;
	WX5726<= not WX6149;
	WX5727<= not WX6151;
	WX5728<= not WX6153;
	WX5729<= not WX6155;
	WX5730<= not WX6157;
	WX5731<= not WX6159;
	WX5732<= not WX6161;
	WX5733<= not WX6163;
	WX5734<= not WX6165;
	WX5735<= not WX6167;
	WX5736<= not WX6105;
	WX5737<= not WX6107;
	WX5738<= not WX6109;
	WX5739<= not WX6111;
	WX5740<= not WX6113;
	WX5741<= not WX6115;
	WX5742<= not WX6117;
	WX5743<= not WX6119;
	WX5744<= not WX6121;
	WX5745<= not WX6123;
	WX5746<= not WX6125;
	WX5747<= not WX6127;
	WX5748<= not WX6129;
	WX5749<= not WX6131;
	WX5750<= not WX6133;
	WX5751<= not WX6135;
	WX5752<= not WX5720;
	WX5753<= not WX5721;
	WX5754<= not WX5722;
	WX5755<= not WX5723;
	WX5756<= not WX5724;
	WX5757<= not WX5725;
	WX5758<= not WX5726;
	WX5759<= not WX5727;
	WX5760<= not WX5728;
	WX5761<= not WX5729;
	WX5762<= not WX5730;
	WX5763<= not WX5731;
	WX5764<= not WX5732;
	WX5765<= not WX5733;
	WX5766<= not WX5734;
	WX5767<= not WX5735;
	WX5768<= not WX5736;
	WX5769<= not WX5737;
	WX5770<= not WX5738;
	WX5771<= not WX5739;
	WX5772<= not WX5740;
	WX5773<= not WX5741;
	WX5774<= not WX5742;
	WX5775<= not WX5743;
	WX5776<= not WX5744;
	WX5777<= not WX5745;
	WX5778<= not WX5746;
	WX5779<= not WX5747;
	WX5780<= not WX5748;
	WX5781<= not WX5749;
	WX5782<= not WX5750;
	WX5783<= not WX5751;
	WX5784<= not WX6009;
	WX5785<= not WX6011;
	WX5786<= not WX6013;
	WX5787<= not WX6015;
	WX5788<= not WX6017;
	WX5789<= not WX6019;
	WX5790<= not WX6021;
	WX5791<= not WX6023;
	WX5792<= not WX6025;
	WX5793<= not WX6027;
	WX5794<= not WX6029;
	WX5795<= not WX6031;
	WX5796<= not WX6033;
	WX5797<= not WX6035;
	WX5798<= not WX6037;
	WX5799<= not WX6039;
	WX5800<= not WX6041;
	WX5801<= not WX6043;
	WX5802<= not WX6045;
	WX5803<= not WX6047;
	WX5804<= not WX6049;
	WX5805<= not WX6051;
	WX5806<= not WX6053;
	WX5807<= not WX6055;
	WX5808<= not WX6057;
	WX5809<= not WX6059;
	WX5810<= not WX6061;
	WX5811<= not WX6063;
	WX5812<= not WX6065;
	WX5813<= not WX6067;
	WX5814<= not WX6069;
	WX5815<= not WX6071;
	WX6104<= not WX6088;
	WX6105<= not WX6104;
	WX6106<= not WX6089;
	WX6107<= not WX6106;
	WX6108<= not WX6090;
	WX6109<= not WX6108;
	WX6110<= not WX6091;
	WX6111<= not WX6110;
	WX6112<= not WX6092;
	WX6113<= not WX6112;
	WX6114<= not WX6093;
	WX6115<= not WX6114;
	WX6116<= not WX6094;
	WX6117<= not WX6116;
	WX6118<= not WX6095;
	WX6119<= not WX6118;
	WX6120<= not WX6096;
	WX6121<= not WX6120;
	WX6122<= not WX6097;
	WX6123<= not WX6122;
	WX6124<= not WX6098;
	WX6125<= not WX6124;
	WX6126<= not WX6099;
	WX6127<= not WX6126;
	WX6128<= not WX6100;
	WX6129<= not WX6128;
	WX6130<= not WX6101;
	WX6131<= not WX6130;
	WX6132<= not WX6102;
	WX6133<= not WX6132;
	WX6134<= not WX6103;
	WX6135<= not WX6134;
	WX6136<= not WX6072;
	WX6137<= not WX6136;
	WX6138<= not WX6073;
	WX6139<= not WX6138;
	WX6140<= not WX6074;
	WX6141<= not WX6140;
	WX6142<= not WX6075;
	WX6143<= not WX6142;
	WX6144<= not WX6076;
	WX6145<= not WX6144;
	WX6146<= not WX6077;
	WX6147<= not WX6146;
	WX6148<= not WX6078;
	WX6149<= not WX6148;
	WX6150<= not WX6079;
	WX6151<= not WX6150;
	WX6152<= not WX6080;
	WX6153<= not WX6152;
	WX6154<= not WX6081;
	WX6155<= not WX6154;
	WX6156<= not WX6082;
	WX6157<= not WX6156;
	WX6158<= not WX6083;
	WX6159<= not WX6158;
	WX6160<= not WX6084;
	WX6161<= not WX6160;
	WX6162<= not WX6085;
	WX6163<= not WX6162;
	WX6164<= not WX6086;
	WX6165<= not WX6164;
	WX6166<= not WX6087;
	WX6167<= not WX6166;
	WX6168<= not TM0;
	WX6169<= not TM0;
	WX6170<= not TM0;
	WX6171<= not TM1;
	WX6172<= not TM1;
	WX6173<= not WX6172;
	WX6174<= not WX6170;
	WX6175<= not WX6171;
	WX6176<= not WX6169;
	WX6177<= not WX6168;
	WX6181<= not WX6177;
	WX6183<= not WX6182;
	WX6184<= not WX6183;
	WX6188<= not WX6177;
	WX6190<= not WX6189;
	WX6191<= not WX6190;
	WX6195<= not WX6177;
	WX6197<= not WX6196;
	WX6198<= not WX6197;
	WX6202<= not WX6177;
	WX6204<= not WX6203;
	WX6205<= not WX6204;
	WX6209<= not WX6177;
	WX6211<= not WX6210;
	WX6212<= not WX6211;
	WX6216<= not WX6177;
	WX6218<= not WX6217;
	WX6219<= not WX6218;
	WX6223<= not WX6177;
	WX6225<= not WX6224;
	WX6226<= not WX6225;
	WX6230<= not WX6177;
	WX6232<= not WX6231;
	WX6233<= not WX6232;
	WX6237<= not WX6177;
	WX6239<= not WX6238;
	WX6240<= not WX6239;
	WX6244<= not WX6177;
	WX6246<= not WX6245;
	WX6247<= not WX6246;
	WX6251<= not WX6177;
	WX6253<= not WX6252;
	WX6254<= not WX6253;
	WX6258<= not WX6177;
	WX6260<= not WX6259;
	WX6261<= not WX6260;
	WX6265<= not WX6177;
	WX6267<= not WX6266;
	WX6268<= not WX6267;
	WX6272<= not WX6177;
	WX6274<= not WX6273;
	WX6275<= not WX6274;
	WX6279<= not WX6177;
	WX6281<= not WX6280;
	WX6282<= not WX6281;
	WX6286<= not WX6177;
	WX6288<= not WX6287;
	WX6289<= not WX6288;
	WX6293<= not WX6177;
	WX6295<= not WX6294;
	WX6296<= not WX6295;
	WX6300<= not WX6177;
	WX6302<= not WX6301;
	WX6303<= not WX6302;
	WX6307<= not WX6177;
	WX6309<= not WX6308;
	WX6310<= not WX6309;
	WX6314<= not WX6177;
	WX6316<= not WX6315;
	WX6317<= not WX6316;
	WX6321<= not WX6177;
	WX6323<= not WX6322;
	WX6324<= not WX6323;
	WX6328<= not WX6177;
	WX6330<= not WX6329;
	WX6331<= not WX6330;
	WX6335<= not WX6177;
	WX6337<= not WX6336;
	WX6338<= not WX6337;
	WX6342<= not WX6177;
	WX6344<= not WX6343;
	WX6345<= not WX6344;
	WX6349<= not WX6177;
	WX6351<= not WX6350;
	WX6352<= not WX6351;
	WX6356<= not WX6177;
	WX6358<= not WX6357;
	WX6359<= not WX6358;
	WX6363<= not WX6177;
	WX6365<= not WX6364;
	WX6366<= not WX6365;
	WX6370<= not WX6177;
	WX6372<= not WX6371;
	WX6373<= not WX6372;
	WX6377<= not WX6177;
	WX6379<= not WX6378;
	WX6380<= not WX6379;
	WX6384<= not WX6177;
	WX6386<= not WX6385;
	WX6387<= not WX6386;
	WX6391<= not WX6177;
	WX6393<= not WX6392;
	WX6394<= not WX6393;
	WX6398<= not WX6177;
	WX6400<= not WX6399;
	WX6401<= not WX6400;
	WX6402<= not RESET;
	WX6435<= not WX6402;
	WX6502<= not WX7468;
	WX6506<= not WX7469;
	WX6510<= not WX7469;
	WX6512<= not WX6503;
	WX6513<= not WX6512;
	WX6516<= not WX7468;
	WX6520<= not WX7469;
	WX6524<= not WX7469;
	WX6526<= not WX6517;
	WX6527<= not WX6526;
	WX6530<= not WX7468;
	WX6534<= not WX7469;
	WX6538<= not WX7469;
	WX6540<= not WX6531;
	WX6541<= not WX6540;
	WX6544<= not WX7468;
	WX6548<= not WX7469;
	WX6552<= not WX7469;
	WX6554<= not WX6545;
	WX6555<= not WX6554;
	WX6558<= not WX7468;
	WX6562<= not WX7469;
	WX6566<= not WX7469;
	WX6568<= not WX6559;
	WX6569<= not WX6568;
	WX6572<= not WX7468;
	WX6576<= not WX7469;
	WX6580<= not WX7469;
	WX6582<= not WX6573;
	WX6583<= not WX6582;
	WX6586<= not WX7468;
	WX6590<= not WX7469;
	WX6594<= not WX7469;
	WX6596<= not WX6587;
	WX6597<= not WX6596;
	WX6600<= not WX7468;
	WX6604<= not WX7469;
	WX6608<= not WX7469;
	WX6610<= not WX6601;
	WX6611<= not WX6610;
	WX6614<= not WX7468;
	WX6618<= not WX7469;
	WX6622<= not WX7469;
	WX6624<= not WX6615;
	WX6625<= not WX6624;
	WX6628<= not WX7468;
	WX6632<= not WX7469;
	WX6636<= not WX7469;
	WX6638<= not WX6629;
	WX6639<= not WX6638;
	WX6642<= not WX7468;
	WX6646<= not WX7469;
	WX6650<= not WX7469;
	WX6652<= not WX6643;
	WX6653<= not WX6652;
	WX6656<= not WX7468;
	WX6660<= not WX7469;
	WX6664<= not WX7469;
	WX6666<= not WX6657;
	WX6667<= not WX6666;
	WX6670<= not WX7468;
	WX6674<= not WX7469;
	WX6678<= not WX7469;
	WX6680<= not WX6671;
	WX6681<= not WX6680;
	WX6684<= not WX7468;
	WX6688<= not WX7469;
	WX6692<= not WX7469;
	WX6694<= not WX6685;
	WX6695<= not WX6694;
	WX6698<= not WX7468;
	WX6702<= not WX7469;
	WX6706<= not WX7469;
	WX6708<= not WX6699;
	WX6709<= not WX6708;
	WX6712<= not WX7468;
	WX6716<= not WX7469;
	WX6720<= not WX7469;
	WX6722<= not WX6713;
	WX6723<= not WX6722;
	WX6726<= not WX7468;
	WX6730<= not WX7469;
	WX6734<= not WX7469;
	WX6736<= not WX6727;
	WX6737<= not WX6736;
	WX6740<= not WX7468;
	WX6744<= not WX7469;
	WX6748<= not WX7469;
	WX6750<= not WX6741;
	WX6751<= not WX6750;
	WX6754<= not WX7468;
	WX6758<= not WX7469;
	WX6762<= not WX7469;
	WX6764<= not WX6755;
	WX6765<= not WX6764;
	WX6768<= not WX7468;
	WX6772<= not WX7469;
	WX6776<= not WX7469;
	WX6778<= not WX6769;
	WX6779<= not WX6778;
	WX6782<= not WX7468;
	WX6786<= not WX7469;
	WX6790<= not WX7469;
	WX6792<= not WX6783;
	WX6793<= not WX6792;
	WX6796<= not WX7468;
	WX6800<= not WX7469;
	WX6804<= not WX7469;
	WX6806<= not WX6797;
	WX6807<= not WX6806;
	WX6810<= not WX7468;
	WX6814<= not WX7469;
	WX6818<= not WX7469;
	WX6820<= not WX6811;
	WX6821<= not WX6820;
	WX6824<= not WX7468;
	WX6828<= not WX7469;
	WX6832<= not WX7469;
	WX6834<= not WX6825;
	WX6835<= not WX6834;
	WX6838<= not WX7468;
	WX6842<= not WX7469;
	WX6846<= not WX7469;
	WX6848<= not WX6839;
	WX6849<= not WX6848;
	WX6852<= not WX7468;
	WX6856<= not WX7469;
	WX6860<= not WX7469;
	WX6862<= not WX6853;
	WX6863<= not WX6862;
	WX6866<= not WX7468;
	WX6870<= not WX7469;
	WX6874<= not WX7469;
	WX6876<= not WX6867;
	WX6877<= not WX6876;
	WX6880<= not WX7468;
	WX6884<= not WX7469;
	WX6888<= not WX7469;
	WX6890<= not WX6881;
	WX6891<= not WX6890;
	WX6894<= not WX7468;
	WX6898<= not WX7469;
	WX6902<= not WX7469;
	WX6904<= not WX6895;
	WX6905<= not WX6904;
	WX6908<= not WX7468;
	WX6912<= not WX7469;
	WX6916<= not WX7469;
	WX6918<= not WX6909;
	WX6919<= not WX6918;
	WX6922<= not WX7468;
	WX6926<= not WX7469;
	WX6930<= not WX7469;
	WX6932<= not WX6923;
	WX6933<= not WX6932;
	WX6936<= not WX7468;
	WX6940<= not WX7469;
	WX6944<= not WX7469;
	WX6946<= not WX6937;
	WX6947<= not WX6946;
	WX6948<= not WX6950;
	WX7013<= not WX7430;
	WX7014<= not WX7432;
	WX7015<= not WX7434;
	WX7016<= not WX7436;
	WX7017<= not WX7438;
	WX7018<= not WX7440;
	WX7019<= not WX7442;
	WX7020<= not WX7444;
	WX7021<= not WX7446;
	WX7022<= not WX7448;
	WX7023<= not WX7450;
	WX7024<= not WX7452;
	WX7025<= not WX7454;
	WX7026<= not WX7456;
	WX7027<= not WX7458;
	WX7028<= not WX7460;
	WX7029<= not WX7398;
	WX7030<= not WX7400;
	WX7031<= not WX7402;
	WX7032<= not WX7404;
	WX7033<= not WX7406;
	WX7034<= not WX7408;
	WX7035<= not WX7410;
	WX7036<= not WX7412;
	WX7037<= not WX7414;
	WX7038<= not WX7416;
	WX7039<= not WX7418;
	WX7040<= not WX7420;
	WX7041<= not WX7422;
	WX7042<= not WX7424;
	WX7043<= not WX7426;
	WX7044<= not WX7428;
	WX7045<= not WX7013;
	WX7046<= not WX7014;
	WX7047<= not WX7015;
	WX7048<= not WX7016;
	WX7049<= not WX7017;
	WX7050<= not WX7018;
	WX7051<= not WX7019;
	WX7052<= not WX7020;
	WX7053<= not WX7021;
	WX7054<= not WX7022;
	WX7055<= not WX7023;
	WX7056<= not WX7024;
	WX7057<= not WX7025;
	WX7058<= not WX7026;
	WX7059<= not WX7027;
	WX7060<= not WX7028;
	WX7061<= not WX7029;
	WX7062<= not WX7030;
	WX7063<= not WX7031;
	WX7064<= not WX7032;
	WX7065<= not WX7033;
	WX7066<= not WX7034;
	WX7067<= not WX7035;
	WX7068<= not WX7036;
	WX7069<= not WX7037;
	WX7070<= not WX7038;
	WX7071<= not WX7039;
	WX7072<= not WX7040;
	WX7073<= not WX7041;
	WX7074<= not WX7042;
	WX7075<= not WX7043;
	WX7076<= not WX7044;
	WX7077<= not WX7302;
	WX7078<= not WX7304;
	WX7079<= not WX7306;
	WX7080<= not WX7308;
	WX7081<= not WX7310;
	WX7082<= not WX7312;
	WX7083<= not WX7314;
	WX7084<= not WX7316;
	WX7085<= not WX7318;
	WX7086<= not WX7320;
	WX7087<= not WX7322;
	WX7088<= not WX7324;
	WX7089<= not WX7326;
	WX7090<= not WX7328;
	WX7091<= not WX7330;
	WX7092<= not WX7332;
	WX7093<= not WX7334;
	WX7094<= not WX7336;
	WX7095<= not WX7338;
	WX7096<= not WX7340;
	WX7097<= not WX7342;
	WX7098<= not WX7344;
	WX7099<= not WX7346;
	WX7100<= not WX7348;
	WX7101<= not WX7350;
	WX7102<= not WX7352;
	WX7103<= not WX7354;
	WX7104<= not WX7356;
	WX7105<= not WX7358;
	WX7106<= not WX7360;
	WX7107<= not WX7362;
	WX7108<= not WX7364;
	WX7397<= not WX7381;
	WX7398<= not WX7397;
	WX7399<= not WX7382;
	WX7400<= not WX7399;
	WX7401<= not WX7383;
	WX7402<= not WX7401;
	WX7403<= not WX7384;
	WX7404<= not WX7403;
	WX7405<= not WX7385;
	WX7406<= not WX7405;
	WX7407<= not WX7386;
	WX7408<= not WX7407;
	WX7409<= not WX7387;
	WX7410<= not WX7409;
	WX7411<= not WX7388;
	WX7412<= not WX7411;
	WX7413<= not WX7389;
	WX7414<= not WX7413;
	WX7415<= not WX7390;
	WX7416<= not WX7415;
	WX7417<= not WX7391;
	WX7418<= not WX7417;
	WX7419<= not WX7392;
	WX7420<= not WX7419;
	WX7421<= not WX7393;
	WX7422<= not WX7421;
	WX7423<= not WX7394;
	WX7424<= not WX7423;
	WX7425<= not WX7395;
	WX7426<= not WX7425;
	WX7427<= not WX7396;
	WX7428<= not WX7427;
	WX7429<= not WX7365;
	WX7430<= not WX7429;
	WX7431<= not WX7366;
	WX7432<= not WX7431;
	WX7433<= not WX7367;
	WX7434<= not WX7433;
	WX7435<= not WX7368;
	WX7436<= not WX7435;
	WX7437<= not WX7369;
	WX7438<= not WX7437;
	WX7439<= not WX7370;
	WX7440<= not WX7439;
	WX7441<= not WX7371;
	WX7442<= not WX7441;
	WX7443<= not WX7372;
	WX7444<= not WX7443;
	WX7445<= not WX7373;
	WX7446<= not WX7445;
	WX7447<= not WX7374;
	WX7448<= not WX7447;
	WX7449<= not WX7375;
	WX7450<= not WX7449;
	WX7451<= not WX7376;
	WX7452<= not WX7451;
	WX7453<= not WX7377;
	WX7454<= not WX7453;
	WX7455<= not WX7378;
	WX7456<= not WX7455;
	WX7457<= not WX7379;
	WX7458<= not WX7457;
	WX7459<= not WX7380;
	WX7460<= not WX7459;
	WX7461<= not TM0;
	WX7462<= not TM0;
	WX7463<= not TM0;
	WX7464<= not TM1;
	WX7465<= not TM1;
	WX7466<= not WX7465;
	WX7467<= not WX7463;
	WX7468<= not WX7464;
	WX7469<= not WX7462;
	WX7470<= not WX7461;
	WX7474<= not WX7470;
	WX7476<= not WX7475;
	WX7477<= not WX7476;
	WX7481<= not WX7470;
	WX7483<= not WX7482;
	WX7484<= not WX7483;
	WX7488<= not WX7470;
	WX7490<= not WX7489;
	WX7491<= not WX7490;
	WX7495<= not WX7470;
	WX7497<= not WX7496;
	WX7498<= not WX7497;
	WX7502<= not WX7470;
	WX7504<= not WX7503;
	WX7505<= not WX7504;
	WX7509<= not WX7470;
	WX7511<= not WX7510;
	WX7512<= not WX7511;
	WX7516<= not WX7470;
	WX7518<= not WX7517;
	WX7519<= not WX7518;
	WX7523<= not WX7470;
	WX7525<= not WX7524;
	WX7526<= not WX7525;
	WX7530<= not WX7470;
	WX7532<= not WX7531;
	WX7533<= not WX7532;
	WX7537<= not WX7470;
	WX7539<= not WX7538;
	WX7540<= not WX7539;
	WX7544<= not WX7470;
	WX7546<= not WX7545;
	WX7547<= not WX7546;
	WX7551<= not WX7470;
	WX7553<= not WX7552;
	WX7554<= not WX7553;
	WX7558<= not WX7470;
	WX7560<= not WX7559;
	WX7561<= not WX7560;
	WX7565<= not WX7470;
	WX7567<= not WX7566;
	WX7568<= not WX7567;
	WX7572<= not WX7470;
	WX7574<= not WX7573;
	WX7575<= not WX7574;
	WX7579<= not WX7470;
	WX7581<= not WX7580;
	WX7582<= not WX7581;
	WX7586<= not WX7470;
	WX7588<= not WX7587;
	WX7589<= not WX7588;
	WX7593<= not WX7470;
	WX7595<= not WX7594;
	WX7596<= not WX7595;
	WX7600<= not WX7470;
	WX7602<= not WX7601;
	WX7603<= not WX7602;
	WX7607<= not WX7470;
	WX7609<= not WX7608;
	WX7610<= not WX7609;
	WX7614<= not WX7470;
	WX7616<= not WX7615;
	WX7617<= not WX7616;
	WX7621<= not WX7470;
	WX7623<= not WX7622;
	WX7624<= not WX7623;
	WX7628<= not WX7470;
	WX7630<= not WX7629;
	WX7631<= not WX7630;
	WX7635<= not WX7470;
	WX7637<= not WX7636;
	WX7638<= not WX7637;
	WX7642<= not WX7470;
	WX7644<= not WX7643;
	WX7645<= not WX7644;
	WX7649<= not WX7470;
	WX7651<= not WX7650;
	WX7652<= not WX7651;
	WX7656<= not WX7470;
	WX7658<= not WX7657;
	WX7659<= not WX7658;
	WX7663<= not WX7470;
	WX7665<= not WX7664;
	WX7666<= not WX7665;
	WX7670<= not WX7470;
	WX7672<= not WX7671;
	WX7673<= not WX7672;
	WX7677<= not WX7470;
	WX7679<= not WX7678;
	WX7680<= not WX7679;
	WX7684<= not WX7470;
	WX7686<= not WX7685;
	WX7687<= not WX7686;
	WX7691<= not WX7470;
	WX7693<= not WX7692;
	WX7694<= not WX7693;
	WX7695<= not RESET;
	WX7728<= not WX7695;
	WX7795<= not WX8761;
	WX7799<= not WX8762;
	WX7803<= not WX8762;
	WX7805<= not WX7796;
	WX7806<= not WX7805;
	WX7809<= not WX8761;
	WX7813<= not WX8762;
	WX7817<= not WX8762;
	WX7819<= not WX7810;
	WX7820<= not WX7819;
	WX7823<= not WX8761;
	WX7827<= not WX8762;
	WX7831<= not WX8762;
	WX7833<= not WX7824;
	WX7834<= not WX7833;
	WX7837<= not WX8761;
	WX7841<= not WX8762;
	WX7845<= not WX8762;
	WX7847<= not WX7838;
	WX7848<= not WX7847;
	WX7851<= not WX8761;
	WX7855<= not WX8762;
	WX7859<= not WX8762;
	WX7861<= not WX7852;
	WX7862<= not WX7861;
	WX7865<= not WX8761;
	WX7869<= not WX8762;
	WX7873<= not WX8762;
	WX7875<= not WX7866;
	WX7876<= not WX7875;
	WX7879<= not WX8761;
	WX7883<= not WX8762;
	WX7887<= not WX8762;
	WX7889<= not WX7880;
	WX7890<= not WX7889;
	WX7893<= not WX8761;
	WX7897<= not WX8762;
	WX7901<= not WX8762;
	WX7903<= not WX7894;
	WX7904<= not WX7903;
	WX7907<= not WX8761;
	WX7911<= not WX8762;
	WX7915<= not WX8762;
	WX7917<= not WX7908;
	WX7918<= not WX7917;
	WX7921<= not WX8761;
	WX7925<= not WX8762;
	WX7929<= not WX8762;
	WX7931<= not WX7922;
	WX7932<= not WX7931;
	WX7935<= not WX8761;
	WX7939<= not WX8762;
	WX7943<= not WX8762;
	WX7945<= not WX7936;
	WX7946<= not WX7945;
	WX7949<= not WX8761;
	WX7953<= not WX8762;
	WX7957<= not WX8762;
	WX7959<= not WX7950;
	WX7960<= not WX7959;
	WX7963<= not WX8761;
	WX7967<= not WX8762;
	WX7971<= not WX8762;
	WX7973<= not WX7964;
	WX7974<= not WX7973;
	WX7977<= not WX8761;
	WX7981<= not WX8762;
	WX7985<= not WX8762;
	WX7987<= not WX7978;
	WX7988<= not WX7987;
	WX7991<= not WX8761;
	WX7995<= not WX8762;
	WX7999<= not WX8762;
	WX8001<= not WX7992;
	WX8002<= not WX8001;
	WX8005<= not WX8761;
	WX8009<= not WX8762;
	WX8013<= not WX8762;
	WX8015<= not WX8006;
	WX8016<= not WX8015;
	WX8019<= not WX8761;
	WX8023<= not WX8762;
	WX8027<= not WX8762;
	WX8029<= not WX8020;
	WX8030<= not WX8029;
	WX8033<= not WX8761;
	WX8037<= not WX8762;
	WX8041<= not WX8762;
	WX8043<= not WX8034;
	WX8044<= not WX8043;
	WX8047<= not WX8761;
	WX8051<= not WX8762;
	WX8055<= not WX8762;
	WX8057<= not WX8048;
	WX8058<= not WX8057;
	WX8061<= not WX8761;
	WX8065<= not WX8762;
	WX8069<= not WX8762;
	WX8071<= not WX8062;
	WX8072<= not WX8071;
	WX8075<= not WX8761;
	WX8079<= not WX8762;
	WX8083<= not WX8762;
	WX8085<= not WX8076;
	WX8086<= not WX8085;
	WX8089<= not WX8761;
	WX8093<= not WX8762;
	WX8097<= not WX8762;
	WX8099<= not WX8090;
	WX8100<= not WX8099;
	WX8103<= not WX8761;
	WX8107<= not WX8762;
	WX8111<= not WX8762;
	WX8113<= not WX8104;
	WX8114<= not WX8113;
	WX8117<= not WX8761;
	WX8121<= not WX8762;
	WX8125<= not WX8762;
	WX8127<= not WX8118;
	WX8128<= not WX8127;
	WX8131<= not WX8761;
	WX8135<= not WX8762;
	WX8139<= not WX8762;
	WX8141<= not WX8132;
	WX8142<= not WX8141;
	WX8145<= not WX8761;
	WX8149<= not WX8762;
	WX8153<= not WX8762;
	WX8155<= not WX8146;
	WX8156<= not WX8155;
	WX8159<= not WX8761;
	WX8163<= not WX8762;
	WX8167<= not WX8762;
	WX8169<= not WX8160;
	WX8170<= not WX8169;
	WX8173<= not WX8761;
	WX8177<= not WX8762;
	WX8181<= not WX8762;
	WX8183<= not WX8174;
	WX8184<= not WX8183;
	WX8187<= not WX8761;
	WX8191<= not WX8762;
	WX8195<= not WX8762;
	WX8197<= not WX8188;
	WX8198<= not WX8197;
	WX8201<= not WX8761;
	WX8205<= not WX8762;
	WX8209<= not WX8762;
	WX8211<= not WX8202;
	WX8212<= not WX8211;
	WX8215<= not WX8761;
	WX8219<= not WX8762;
	WX8223<= not WX8762;
	WX8225<= not WX8216;
	WX8226<= not WX8225;
	WX8229<= not WX8761;
	WX8233<= not WX8762;
	WX8237<= not WX8762;
	WX8239<= not WX8230;
	WX8240<= not WX8239;
	WX8241<= not WX8243;
	WX8306<= not WX8723;
	WX8307<= not WX8725;
	WX8308<= not WX8727;
	WX8309<= not WX8729;
	WX8310<= not WX8731;
	WX8311<= not WX8733;
	WX8312<= not WX8735;
	WX8313<= not WX8737;
	WX8314<= not WX8739;
	WX8315<= not WX8741;
	WX8316<= not WX8743;
	WX8317<= not WX8745;
	WX8318<= not WX8747;
	WX8319<= not WX8749;
	WX8320<= not WX8751;
	WX8321<= not WX8753;
	WX8322<= not WX8691;
	WX8323<= not WX8693;
	WX8324<= not WX8695;
	WX8325<= not WX8697;
	WX8326<= not WX8699;
	WX8327<= not WX8701;
	WX8328<= not WX8703;
	WX8329<= not WX8705;
	WX8330<= not WX8707;
	WX8331<= not WX8709;
	WX8332<= not WX8711;
	WX8333<= not WX8713;
	WX8334<= not WX8715;
	WX8335<= not WX8717;
	WX8336<= not WX8719;
	WX8337<= not WX8721;
	WX8338<= not WX8306;
	WX8339<= not WX8307;
	WX8340<= not WX8308;
	WX8341<= not WX8309;
	WX8342<= not WX8310;
	WX8343<= not WX8311;
	WX8344<= not WX8312;
	WX8345<= not WX8313;
	WX8346<= not WX8314;
	WX8347<= not WX8315;
	WX8348<= not WX8316;
	WX8349<= not WX8317;
	WX8350<= not WX8318;
	WX8351<= not WX8319;
	WX8352<= not WX8320;
	WX8353<= not WX8321;
	WX8354<= not WX8322;
	WX8355<= not WX8323;
	WX8356<= not WX8324;
	WX8357<= not WX8325;
	WX8358<= not WX8326;
	WX8359<= not WX8327;
	WX8360<= not WX8328;
	WX8361<= not WX8329;
	WX8362<= not WX8330;
	WX8363<= not WX8331;
	WX8364<= not WX8332;
	WX8365<= not WX8333;
	WX8366<= not WX8334;
	WX8367<= not WX8335;
	WX8368<= not WX8336;
	WX8369<= not WX8337;
	WX8370<= not WX8595;
	WX8371<= not WX8597;
	WX8372<= not WX8599;
	WX8373<= not WX8601;
	WX8374<= not WX8603;
	WX8375<= not WX8605;
	WX8376<= not WX8607;
	WX8377<= not WX8609;
	WX8378<= not WX8611;
	WX8379<= not WX8613;
	WX8380<= not WX8615;
	WX8381<= not WX8617;
	WX8382<= not WX8619;
	WX8383<= not WX8621;
	WX8384<= not WX8623;
	WX8385<= not WX8625;
	WX8386<= not WX8627;
	WX8387<= not WX8629;
	WX8388<= not WX8631;
	WX8389<= not WX8633;
	WX8390<= not WX8635;
	WX8391<= not WX8637;
	WX8392<= not WX8639;
	WX8393<= not WX8641;
	WX8394<= not WX8643;
	WX8395<= not WX8645;
	WX8396<= not WX8647;
	WX8397<= not WX8649;
	WX8398<= not WX8651;
	WX8399<= not WX8653;
	WX8400<= not WX8655;
	WX8401<= not WX8657;
	WX8690<= not WX8674;
	WX8691<= not WX8690;
	WX8692<= not WX8675;
	WX8693<= not WX8692;
	WX8694<= not WX8676;
	WX8695<= not WX8694;
	WX8696<= not WX8677;
	WX8697<= not WX8696;
	WX8698<= not WX8678;
	WX8699<= not WX8698;
	WX8700<= not WX8679;
	WX8701<= not WX8700;
	WX8702<= not WX8680;
	WX8703<= not WX8702;
	WX8704<= not WX8681;
	WX8705<= not WX8704;
	WX8706<= not WX8682;
	WX8707<= not WX8706;
	WX8708<= not WX8683;
	WX8709<= not WX8708;
	WX8710<= not WX8684;
	WX8711<= not WX8710;
	WX8712<= not WX8685;
	WX8713<= not WX8712;
	WX8714<= not WX8686;
	WX8715<= not WX8714;
	WX8716<= not WX8687;
	WX8717<= not WX8716;
	WX8718<= not WX8688;
	WX8719<= not WX8718;
	WX8720<= not WX8689;
	WX8721<= not WX8720;
	WX8722<= not WX8658;
	WX8723<= not WX8722;
	WX8724<= not WX8659;
	WX8725<= not WX8724;
	WX8726<= not WX8660;
	WX8727<= not WX8726;
	WX8728<= not WX8661;
	WX8729<= not WX8728;
	WX8730<= not WX8662;
	WX8731<= not WX8730;
	WX8732<= not WX8663;
	WX8733<= not WX8732;
	WX8734<= not WX8664;
	WX8735<= not WX8734;
	WX8736<= not WX8665;
	WX8737<= not WX8736;
	WX8738<= not WX8666;
	WX8739<= not WX8738;
	WX8740<= not WX8667;
	WX8741<= not WX8740;
	WX8742<= not WX8668;
	WX8743<= not WX8742;
	WX8744<= not WX8669;
	WX8745<= not WX8744;
	WX8746<= not WX8670;
	WX8747<= not WX8746;
	WX8748<= not WX8671;
	WX8749<= not WX8748;
	WX8750<= not WX8672;
	WX8751<= not WX8750;
	WX8752<= not WX8673;
	WX8753<= not WX8752;
	WX8754<= not TM0;
	WX8755<= not TM0;
	WX8756<= not TM0;
	WX8757<= not TM1;
	WX8758<= not TM1;
	WX8759<= not WX8758;
	WX8760<= not WX8756;
	WX8761<= not WX8757;
	WX8762<= not WX8755;
	WX8763<= not WX8754;
	WX8767<= not WX8763;
	WX8769<= not WX8768;
	WX8770<= not WX8769;
	WX8774<= not WX8763;
	WX8776<= not WX8775;
	WX8777<= not WX8776;
	WX8781<= not WX8763;
	WX8783<= not WX8782;
	WX8784<= not WX8783;
	WX8788<= not WX8763;
	WX8790<= not WX8789;
	WX8791<= not WX8790;
	WX8795<= not WX8763;
	WX8797<= not WX8796;
	WX8798<= not WX8797;
	WX8802<= not WX8763;
	WX8804<= not WX8803;
	WX8805<= not WX8804;
	WX8809<= not WX8763;
	WX8811<= not WX8810;
	WX8812<= not WX8811;
	WX8816<= not WX8763;
	WX8818<= not WX8817;
	WX8819<= not WX8818;
	WX8823<= not WX8763;
	WX8825<= not WX8824;
	WX8826<= not WX8825;
	WX8830<= not WX8763;
	WX8832<= not WX8831;
	WX8833<= not WX8832;
	WX8837<= not WX8763;
	WX8839<= not WX8838;
	WX8840<= not WX8839;
	WX8844<= not WX8763;
	WX8846<= not WX8845;
	WX8847<= not WX8846;
	WX8851<= not WX8763;
	WX8853<= not WX8852;
	WX8854<= not WX8853;
	WX8858<= not WX8763;
	WX8860<= not WX8859;
	WX8861<= not WX8860;
	WX8865<= not WX8763;
	WX8867<= not WX8866;
	WX8868<= not WX8867;
	WX8872<= not WX8763;
	WX8874<= not WX8873;
	WX8875<= not WX8874;
	WX8879<= not WX8763;
	WX8881<= not WX8880;
	WX8882<= not WX8881;
	WX8886<= not WX8763;
	WX8888<= not WX8887;
	WX8889<= not WX8888;
	WX8893<= not WX8763;
	WX8895<= not WX8894;
	WX8896<= not WX8895;
	WX8900<= not WX8763;
	WX8902<= not WX8901;
	WX8903<= not WX8902;
	WX8907<= not WX8763;
	WX8909<= not WX8908;
	WX8910<= not WX8909;
	WX8914<= not WX8763;
	WX8916<= not WX8915;
	WX8917<= not WX8916;
	WX8921<= not WX8763;
	WX8923<= not WX8922;
	WX8924<= not WX8923;
	WX8928<= not WX8763;
	WX8930<= not WX8929;
	WX8931<= not WX8930;
	WX8935<= not WX8763;
	WX8937<= not WX8936;
	WX8938<= not WX8937;
	WX8942<= not WX8763;
	WX8944<= not WX8943;
	WX8945<= not WX8944;
	WX8949<= not WX8763;
	WX8951<= not WX8950;
	WX8952<= not WX8951;
	WX8956<= not WX8763;
	WX8958<= not WX8957;
	WX8959<= not WX8958;
	WX8963<= not WX8763;
	WX8965<= not WX8964;
	WX8966<= not WX8965;
	WX8970<= not WX8763;
	WX8972<= not WX8971;
	WX8973<= not WX8972;
	WX8977<= not WX8763;
	WX8979<= not WX8978;
	WX8980<= not WX8979;
	WX8984<= not WX8763;
	WX8986<= not WX8985;
	WX8987<= not WX8986;
	WX8988<= not RESET;
	WX9021<= not WX8988;
	WX9088<= not WX10054;
	WX9092<= not WX10055;
	WX9096<= not WX10055;
	WX9098<= not WX9089;
	WX9099<= not WX9098;
	WX9102<= not WX10054;
	WX9106<= not WX10055;
	WX9110<= not WX10055;
	WX9112<= not WX9103;
	WX9113<= not WX9112;
	WX9116<= not WX10054;
	WX9120<= not WX10055;
	WX9124<= not WX10055;
	WX9126<= not WX9117;
	WX9127<= not WX9126;
	WX9130<= not WX10054;
	WX9134<= not WX10055;
	WX9138<= not WX10055;
	WX9140<= not WX9131;
	WX9141<= not WX9140;
	WX9144<= not WX10054;
	WX9148<= not WX10055;
	WX9152<= not WX10055;
	WX9154<= not WX9145;
	WX9155<= not WX9154;
	WX9158<= not WX10054;
	WX9162<= not WX10055;
	WX9166<= not WX10055;
	WX9168<= not WX9159;
	WX9169<= not WX9168;
	WX9172<= not WX10054;
	WX9176<= not WX10055;
	WX9180<= not WX10055;
	WX9182<= not WX9173;
	WX9183<= not WX9182;
	WX9186<= not WX10054;
	WX9190<= not WX10055;
	WX9194<= not WX10055;
	WX9196<= not WX9187;
	WX9197<= not WX9196;
	WX9200<= not WX10054;
	WX9204<= not WX10055;
	WX9208<= not WX10055;
	WX9210<= not WX9201;
	WX9211<= not WX9210;
	WX9214<= not WX10054;
	WX9218<= not WX10055;
	WX9222<= not WX10055;
	WX9224<= not WX9215;
	WX9225<= not WX9224;
	WX9228<= not WX10054;
	WX9232<= not WX10055;
	WX9236<= not WX10055;
	WX9238<= not WX9229;
	WX9239<= not WX9238;
	WX9242<= not WX10054;
	WX9246<= not WX10055;
	WX9250<= not WX10055;
	WX9252<= not WX9243;
	WX9253<= not WX9252;
	WX9256<= not WX10054;
	WX9260<= not WX10055;
	WX9264<= not WX10055;
	WX9266<= not WX9257;
	WX9267<= not WX9266;
	WX9270<= not WX10054;
	WX9274<= not WX10055;
	WX9278<= not WX10055;
	WX9280<= not WX9271;
	WX9281<= not WX9280;
	WX9284<= not WX10054;
	WX9288<= not WX10055;
	WX9292<= not WX10055;
	WX9294<= not WX9285;
	WX9295<= not WX9294;
	WX9298<= not WX10054;
	WX9302<= not WX10055;
	WX9306<= not WX10055;
	WX9308<= not WX9299;
	WX9309<= not WX9308;
	WX9312<= not WX10054;
	WX9316<= not WX10055;
	WX9320<= not WX10055;
	WX9322<= not WX9313;
	WX9323<= not WX9322;
	WX9326<= not WX10054;
	WX9330<= not WX10055;
	WX9334<= not WX10055;
	WX9336<= not WX9327;
	WX9337<= not WX9336;
	WX9340<= not WX10054;
	WX9344<= not WX10055;
	WX9348<= not WX10055;
	WX9350<= not WX9341;
	WX9351<= not WX9350;
	WX9354<= not WX10054;
	WX9358<= not WX10055;
	WX9362<= not WX10055;
	WX9364<= not WX9355;
	WX9365<= not WX9364;
	WX9368<= not WX10054;
	WX9372<= not WX10055;
	WX9376<= not WX10055;
	WX9378<= not WX9369;
	WX9379<= not WX9378;
	WX9382<= not WX10054;
	WX9386<= not WX10055;
	WX9390<= not WX10055;
	WX9392<= not WX9383;
	WX9393<= not WX9392;
	WX9396<= not WX10054;
	WX9400<= not WX10055;
	WX9404<= not WX10055;
	WX9406<= not WX9397;
	WX9407<= not WX9406;
	WX9410<= not WX10054;
	WX9414<= not WX10055;
	WX9418<= not WX10055;
	WX9420<= not WX9411;
	WX9421<= not WX9420;
	WX9424<= not WX10054;
	WX9428<= not WX10055;
	WX9432<= not WX10055;
	WX9434<= not WX9425;
	WX9435<= not WX9434;
	WX9438<= not WX10054;
	WX9442<= not WX10055;
	WX9446<= not WX10055;
	WX9448<= not WX9439;
	WX9449<= not WX9448;
	WX9452<= not WX10054;
	WX9456<= not WX10055;
	WX9460<= not WX10055;
	WX9462<= not WX9453;
	WX9463<= not WX9462;
	WX9466<= not WX10054;
	WX9470<= not WX10055;
	WX9474<= not WX10055;
	WX9476<= not WX9467;
	WX9477<= not WX9476;
	WX9480<= not WX10054;
	WX9484<= not WX10055;
	WX9488<= not WX10055;
	WX9490<= not WX9481;
	WX9491<= not WX9490;
	WX9494<= not WX10054;
	WX9498<= not WX10055;
	WX9502<= not WX10055;
	WX9504<= not WX9495;
	WX9505<= not WX9504;
	WX9508<= not WX10054;
	WX9512<= not WX10055;
	WX9516<= not WX10055;
	WX9518<= not WX9509;
	WX9519<= not WX9518;
	WX9522<= not WX10054;
	WX9526<= not WX10055;
	WX9530<= not WX10055;
	WX9532<= not WX9523;
	WX9533<= not WX9532;
	WX9534<= not WX9536;
	WX9599<= not WX10016;
	WX9600<= not WX10018;
	WX9601<= not WX10020;
	WX9602<= not WX10022;
	WX9603<= not WX10024;
	WX9604<= not WX10026;
	WX9605<= not WX10028;
	WX9606<= not WX10030;
	WX9607<= not WX10032;
	WX9608<= not WX10034;
	WX9609<= not WX10036;
	WX9610<= not WX10038;
	WX9611<= not WX10040;
	WX9612<= not WX10042;
	WX9613<= not WX10044;
	WX9614<= not WX10046;
	WX9615<= not WX9984;
	WX9616<= not WX9986;
	WX9617<= not WX9988;
	WX9618<= not WX9990;
	WX9619<= not WX9992;
	WX9620<= not WX9994;
	WX9621<= not WX9996;
	WX9622<= not WX9998;
	WX9623<= not WX10000;
	WX9624<= not WX10002;
	WX9625<= not WX10004;
	WX9626<= not WX10006;
	WX9627<= not WX10008;
	WX9628<= not WX10010;
	WX9629<= not WX10012;
	WX9630<= not WX10014;
	WX9631<= not WX9599;
	WX9632<= not WX9600;
	WX9633<= not WX9601;
	WX9634<= not WX9602;
	WX9635<= not WX9603;
	WX9636<= not WX9604;
	WX9637<= not WX9605;
	WX9638<= not WX9606;
	WX9639<= not WX9607;
	WX9640<= not WX9608;
	WX9641<= not WX9609;
	WX9642<= not WX9610;
	WX9643<= not WX9611;
	WX9644<= not WX9612;
	WX9645<= not WX9613;
	WX9646<= not WX9614;
	WX9647<= not WX9615;
	WX9648<= not WX9616;
	WX9649<= not WX9617;
	WX9650<= not WX9618;
	WX9651<= not WX9619;
	WX9652<= not WX9620;
	WX9653<= not WX9621;
	WX9654<= not WX9622;
	WX9655<= not WX9623;
	WX9656<= not WX9624;
	WX9657<= not WX9625;
	WX9658<= not WX9626;
	WX9659<= not WX9627;
	WX9660<= not WX9628;
	WX9661<= not WX9629;
	WX9662<= not WX9630;
	WX9663<= not WX9888;
	WX9664<= not WX9890;
	WX9665<= not WX9892;
	WX9666<= not WX9894;
	WX9667<= not WX9896;
	WX9668<= not WX9898;
	WX9669<= not WX9900;
	WX9670<= not WX9902;
	WX9671<= not WX9904;
	WX9672<= not WX9906;
	WX9673<= not WX9908;
	WX9674<= not WX9910;
	WX9675<= not WX9912;
	WX9676<= not WX9914;
	WX9677<= not WX9916;
	WX9678<= not WX9918;
	WX9679<= not WX9920;
	WX9680<= not WX9922;
	WX9681<= not WX9924;
	WX9682<= not WX9926;
	WX9683<= not WX9928;
	WX9684<= not WX9930;
	WX9685<= not WX9932;
	WX9686<= not WX9934;
	WX9687<= not WX9936;
	WX9688<= not WX9938;
	WX9689<= not WX9940;
	WX9690<= not WX9942;
	WX9691<= not WX9944;
	WX9692<= not WX9946;
	WX9693<= not WX9948;
	WX9694<= not WX9950;
	WX9983<= not WX9967;
	WX9984<= not WX9983;
	WX9985<= not WX9968;
	WX9986<= not WX9985;
	WX9987<= not WX9969;
	WX9988<= not WX9987;
	WX9989<= not WX9970;
	WX9990<= not WX9989;
	WX9991<= not WX9971;
	WX9992<= not WX9991;
	WX9993<= not WX9972;
	WX9994<= not WX9993;
	WX9995<= not WX9973;
	WX9996<= not WX9995;
	WX9997<= not WX9974;
	WX9998<= not WX9997;
	WX9999<= not WX9975;
	WX10000<= not WX9999;
	WX10001<= not WX9976;
	WX10002<= not WX10001;
	WX10003<= not WX9977;
	WX10004<= not WX10003;
	WX10005<= not WX9978;
	WX10006<= not WX10005;
	WX10007<= not WX9979;
	WX10008<= not WX10007;
	WX10009<= not WX9980;
	WX10010<= not WX10009;
	WX10011<= not WX9981;
	WX10012<= not WX10011;
	WX10013<= not WX9982;
	WX10014<= not WX10013;
	WX10015<= not WX9951;
	WX10016<= not WX10015;
	WX10017<= not WX9952;
	WX10018<= not WX10017;
	WX10019<= not WX9953;
	WX10020<= not WX10019;
	WX10021<= not WX9954;
	WX10022<= not WX10021;
	WX10023<= not WX9955;
	WX10024<= not WX10023;
	WX10025<= not WX9956;
	WX10026<= not WX10025;
	WX10027<= not WX9957;
	WX10028<= not WX10027;
	WX10029<= not WX9958;
	WX10030<= not WX10029;
	WX10031<= not WX9959;
	WX10032<= not WX10031;
	WX10033<= not WX9960;
	WX10034<= not WX10033;
	WX10035<= not WX9961;
	WX10036<= not WX10035;
	WX10037<= not WX9962;
	WX10038<= not WX10037;
	WX10039<= not WX9963;
	WX10040<= not WX10039;
	WX10041<= not WX9964;
	WX10042<= not WX10041;
	WX10043<= not WX9965;
	WX10044<= not WX10043;
	WX10045<= not WX9966;
	WX10046<= not WX10045;
	WX10047<= not TM0;
	WX10048<= not TM0;
	WX10049<= not TM0;
	WX10050<= not TM1;
	WX10051<= not TM1;
	WX10052<= not WX10051;
	WX10053<= not WX10049;
	WX10054<= not WX10050;
	WX10055<= not WX10048;
	WX10056<= not WX10047;
	WX10060<= not WX10056;
	WX10062<= not WX10061;
	WX10063<= not WX10062;
	WX10067<= not WX10056;
	WX10069<= not WX10068;
	WX10070<= not WX10069;
	WX10074<= not WX10056;
	WX10076<= not WX10075;
	WX10077<= not WX10076;
	WX10081<= not WX10056;
	WX10083<= not WX10082;
	WX10084<= not WX10083;
	WX10088<= not WX10056;
	WX10090<= not WX10089;
	WX10091<= not WX10090;
	WX10095<= not WX10056;
	WX10097<= not WX10096;
	WX10098<= not WX10097;
	WX10102<= not WX10056;
	WX10104<= not WX10103;
	WX10105<= not WX10104;
	WX10109<= not WX10056;
	WX10111<= not WX10110;
	WX10112<= not WX10111;
	WX10116<= not WX10056;
	WX10118<= not WX10117;
	WX10119<= not WX10118;
	WX10123<= not WX10056;
	WX10125<= not WX10124;
	WX10126<= not WX10125;
	WX10130<= not WX10056;
	WX10132<= not WX10131;
	WX10133<= not WX10132;
	WX10137<= not WX10056;
	WX10139<= not WX10138;
	WX10140<= not WX10139;
	WX10144<= not WX10056;
	WX10146<= not WX10145;
	WX10147<= not WX10146;
	WX10151<= not WX10056;
	WX10153<= not WX10152;
	WX10154<= not WX10153;
	WX10158<= not WX10056;
	WX10160<= not WX10159;
	WX10161<= not WX10160;
	WX10165<= not WX10056;
	WX10167<= not WX10166;
	WX10168<= not WX10167;
	WX10172<= not WX10056;
	WX10174<= not WX10173;
	WX10175<= not WX10174;
	WX10179<= not WX10056;
	WX10181<= not WX10180;
	WX10182<= not WX10181;
	WX10186<= not WX10056;
	WX10188<= not WX10187;
	WX10189<= not WX10188;
	WX10193<= not WX10056;
	WX10195<= not WX10194;
	WX10196<= not WX10195;
	WX10200<= not WX10056;
	WX10202<= not WX10201;
	WX10203<= not WX10202;
	WX10207<= not WX10056;
	WX10209<= not WX10208;
	WX10210<= not WX10209;
	WX10214<= not WX10056;
	WX10216<= not WX10215;
	WX10217<= not WX10216;
	WX10221<= not WX10056;
	WX10223<= not WX10222;
	WX10224<= not WX10223;
	WX10228<= not WX10056;
	WX10230<= not WX10229;
	WX10231<= not WX10230;
	WX10235<= not WX10056;
	WX10237<= not WX10236;
	WX10238<= not WX10237;
	WX10242<= not WX10056;
	WX10244<= not WX10243;
	WX10245<= not WX10244;
	WX10249<= not WX10056;
	WX10251<= not WX10250;
	WX10252<= not WX10251;
	WX10256<= not WX10056;
	WX10258<= not WX10257;
	WX10259<= not WX10258;
	WX10263<= not WX10056;
	WX10265<= not WX10264;
	WX10266<= not WX10265;
	WX10270<= not WX10056;
	WX10272<= not WX10271;
	WX10273<= not WX10272;
	WX10277<= not WX10056;
	WX10279<= not WX10278;
	WX10280<= not WX10279;
	WX10281<= not RESET;
	WX10314<= not WX10281;
	WX10381<= not WX11347;
	WX10385<= not WX11348;
	WX10389<= not WX11348;
	WX10391<= not WX10382;
	WX10392<= not WX10391;
	WX10395<= not WX11347;
	WX10399<= not WX11348;
	WX10403<= not WX11348;
	WX10405<= not WX10396;
	WX10406<= not WX10405;
	WX10409<= not WX11347;
	WX10413<= not WX11348;
	WX10417<= not WX11348;
	WX10419<= not WX10410;
	WX10420<= not WX10419;
	WX10423<= not WX11347;
	WX10427<= not WX11348;
	WX10431<= not WX11348;
	WX10433<= not WX10424;
	WX10434<= not WX10433;
	WX10437<= not WX11347;
	WX10441<= not WX11348;
	WX10445<= not WX11348;
	WX10447<= not WX10438;
	WX10448<= not WX10447;
	WX10451<= not WX11347;
	WX10455<= not WX11348;
	WX10459<= not WX11348;
	WX10461<= not WX10452;
	WX10462<= not WX10461;
	WX10465<= not WX11347;
	WX10469<= not WX11348;
	WX10473<= not WX11348;
	WX10475<= not WX10466;
	WX10476<= not WX10475;
	WX10479<= not WX11347;
	WX10483<= not WX11348;
	WX10487<= not WX11348;
	WX10489<= not WX10480;
	WX10490<= not WX10489;
	WX10493<= not WX11347;
	WX10497<= not WX11348;
	WX10501<= not WX11348;
	WX10503<= not WX10494;
	WX10504<= not WX10503;
	WX10507<= not WX11347;
	WX10511<= not WX11348;
	WX10515<= not WX11348;
	WX10517<= not WX10508;
	WX10518<= not WX10517;
	WX10521<= not WX11347;
	WX10525<= not WX11348;
	WX10529<= not WX11348;
	WX10531<= not WX10522;
	WX10532<= not WX10531;
	WX10535<= not WX11347;
	WX10539<= not WX11348;
	WX10543<= not WX11348;
	WX10545<= not WX10536;
	WX10546<= not WX10545;
	WX10549<= not WX11347;
	WX10553<= not WX11348;
	WX10557<= not WX11348;
	WX10559<= not WX10550;
	WX10560<= not WX10559;
	WX10563<= not WX11347;
	WX10567<= not WX11348;
	WX10571<= not WX11348;
	WX10573<= not WX10564;
	WX10574<= not WX10573;
	WX10577<= not WX11347;
	WX10581<= not WX11348;
	WX10585<= not WX11348;
	WX10587<= not WX10578;
	WX10588<= not WX10587;
	WX10591<= not WX11347;
	WX10595<= not WX11348;
	WX10599<= not WX11348;
	WX10601<= not WX10592;
	WX10602<= not WX10601;
	WX10605<= not WX11347;
	WX10609<= not WX11348;
	WX10613<= not WX11348;
	WX10615<= not WX10606;
	WX10616<= not WX10615;
	WX10619<= not WX11347;
	WX10623<= not WX11348;
	WX10627<= not WX11348;
	WX10629<= not WX10620;
	WX10630<= not WX10629;
	WX10633<= not WX11347;
	WX10637<= not WX11348;
	WX10641<= not WX11348;
	WX10643<= not WX10634;
	WX10644<= not WX10643;
	WX10647<= not WX11347;
	WX10651<= not WX11348;
	WX10655<= not WX11348;
	WX10657<= not WX10648;
	WX10658<= not WX10657;
	WX10661<= not WX11347;
	WX10665<= not WX11348;
	WX10669<= not WX11348;
	WX10671<= not WX10662;
	WX10672<= not WX10671;
	WX10675<= not WX11347;
	WX10679<= not WX11348;
	WX10683<= not WX11348;
	WX10685<= not WX10676;
	WX10686<= not WX10685;
	WX10689<= not WX11347;
	WX10693<= not WX11348;
	WX10697<= not WX11348;
	WX10699<= not WX10690;
	WX10700<= not WX10699;
	WX10703<= not WX11347;
	WX10707<= not WX11348;
	WX10711<= not WX11348;
	WX10713<= not WX10704;
	WX10714<= not WX10713;
	WX10717<= not WX11347;
	WX10721<= not WX11348;
	WX10725<= not WX11348;
	WX10727<= not WX10718;
	WX10728<= not WX10727;
	WX10731<= not WX11347;
	WX10735<= not WX11348;
	WX10739<= not WX11348;
	WX10741<= not WX10732;
	WX10742<= not WX10741;
	WX10745<= not WX11347;
	WX10749<= not WX11348;
	WX10753<= not WX11348;
	WX10755<= not WX10746;
	WX10756<= not WX10755;
	WX10759<= not WX11347;
	WX10763<= not WX11348;
	WX10767<= not WX11348;
	WX10769<= not WX10760;
	WX10770<= not WX10769;
	WX10773<= not WX11347;
	WX10777<= not WX11348;
	WX10781<= not WX11348;
	WX10783<= not WX10774;
	WX10784<= not WX10783;
	WX10787<= not WX11347;
	WX10791<= not WX11348;
	WX10795<= not WX11348;
	WX10797<= not WX10788;
	WX10798<= not WX10797;
	WX10801<= not WX11347;
	WX10805<= not WX11348;
	WX10809<= not WX11348;
	WX10811<= not WX10802;
	WX10812<= not WX10811;
	WX10815<= not WX11347;
	WX10819<= not WX11348;
	WX10823<= not WX11348;
	WX10825<= not WX10816;
	WX10826<= not WX10825;
	WX10827<= not WX10829;
	WX10892<= not WX11309;
	WX10893<= not WX11311;
	WX10894<= not WX11313;
	WX10895<= not WX11315;
	WX10896<= not WX11317;
	WX10897<= not WX11319;
	WX10898<= not WX11321;
	WX10899<= not WX11323;
	WX10900<= not WX11325;
	WX10901<= not WX11327;
	WX10902<= not WX11329;
	WX10903<= not WX11331;
	WX10904<= not WX11333;
	WX10905<= not WX11335;
	WX10906<= not WX11337;
	WX10907<= not WX11339;
	WX10908<= not WX11277;
	WX10909<= not WX11279;
	WX10910<= not WX11281;
	WX10911<= not WX11283;
	WX10912<= not WX11285;
	WX10913<= not WX11287;
	WX10914<= not WX11289;
	WX10915<= not WX11291;
	WX10916<= not WX11293;
	WX10917<= not WX11295;
	WX10918<= not WX11297;
	WX10919<= not WX11299;
	WX10920<= not WX11301;
	WX10921<= not WX11303;
	WX10922<= not WX11305;
	WX10923<= not WX11307;
	WX10924<= not WX10892;
	WX10925<= not WX10893;
	WX10926<= not WX10894;
	WX10927<= not WX10895;
	WX10928<= not WX10896;
	WX10929<= not WX10897;
	WX10930<= not WX10898;
	WX10931<= not WX10899;
	WX10932<= not WX10900;
	WX10933<= not WX10901;
	WX10934<= not WX10902;
	WX10935<= not WX10903;
	WX10936<= not WX10904;
	WX10937<= not WX10905;
	WX10938<= not WX10906;
	WX10939<= not WX10907;
	WX10940<= not WX10908;
	WX10941<= not WX10909;
	WX10942<= not WX10910;
	WX10943<= not WX10911;
	WX10944<= not WX10912;
	WX10945<= not WX10913;
	WX10946<= not WX10914;
	WX10947<= not WX10915;
	WX10948<= not WX10916;
	WX10949<= not WX10917;
	WX10950<= not WX10918;
	WX10951<= not WX10919;
	WX10952<= not WX10920;
	WX10953<= not WX10921;
	WX10954<= not WX10922;
	WX10955<= not WX10923;
	WX10956<= not WX11181;
	WX10957<= not WX11183;
	WX10958<= not WX11185;
	WX10959<= not WX11187;
	WX10960<= not WX11189;
	WX10961<= not WX11191;
	WX10962<= not WX11193;
	WX10963<= not WX11195;
	WX10964<= not WX11197;
	WX10965<= not WX11199;
	WX10966<= not WX11201;
	WX10967<= not WX11203;
	WX10968<= not WX11205;
	WX10969<= not WX11207;
	WX10970<= not WX11209;
	WX10971<= not WX11211;
	WX10972<= not WX11213;
	WX10973<= not WX11215;
	WX10974<= not WX11217;
	WX10975<= not WX11219;
	WX10976<= not WX11221;
	WX10977<= not WX11223;
	WX10978<= not WX11225;
	WX10979<= not WX11227;
	WX10980<= not WX11229;
	WX10981<= not WX11231;
	WX10982<= not WX11233;
	WX10983<= not WX11235;
	WX10984<= not WX11237;
	WX10985<= not WX11239;
	WX10986<= not WX11241;
	WX10987<= not WX11243;
	WX11276<= not WX11260;
	WX11277<= not WX11276;
	WX11278<= not WX11261;
	WX11279<= not WX11278;
	WX11280<= not WX11262;
	WX11281<= not WX11280;
	WX11282<= not WX11263;
	WX11283<= not WX11282;
	WX11284<= not WX11264;
	WX11285<= not WX11284;
	WX11286<= not WX11265;
	WX11287<= not WX11286;
	WX11288<= not WX11266;
	WX11289<= not WX11288;
	WX11290<= not WX11267;
	WX11291<= not WX11290;
	WX11292<= not WX11268;
	WX11293<= not WX11292;
	WX11294<= not WX11269;
	WX11295<= not WX11294;
	WX11296<= not WX11270;
	WX11297<= not WX11296;
	WX11298<= not WX11271;
	WX11299<= not WX11298;
	WX11300<= not WX11272;
	WX11301<= not WX11300;
	WX11302<= not WX11273;
	WX11303<= not WX11302;
	WX11304<= not WX11274;
	WX11305<= not WX11304;
	WX11306<= not WX11275;
	WX11307<= not WX11306;
	WX11308<= not WX11244;
	WX11309<= not WX11308;
	WX11310<= not WX11245;
	WX11311<= not WX11310;
	WX11312<= not WX11246;
	WX11313<= not WX11312;
	WX11314<= not WX11247;
	WX11315<= not WX11314;
	WX11316<= not WX11248;
	WX11317<= not WX11316;
	WX11318<= not WX11249;
	WX11319<= not WX11318;
	WX11320<= not WX11250;
	WX11321<= not WX11320;
	WX11322<= not WX11251;
	WX11323<= not WX11322;
	WX11324<= not WX11252;
	WX11325<= not WX11324;
	WX11326<= not WX11253;
	WX11327<= not WX11326;
	WX11328<= not WX11254;
	WX11329<= not WX11328;
	WX11330<= not WX11255;
	WX11331<= not WX11330;
	WX11332<= not WX11256;
	WX11333<= not WX11332;
	WX11334<= not WX11257;
	WX11335<= not WX11334;
	WX11336<= not WX11258;
	WX11337<= not WX11336;
	WX11338<= not WX11259;
	WX11339<= not WX11338;
	WX11340<= not TM0;
	WX11341<= not TM0;
	WX11342<= not TM0;
	WX11343<= not TM1;
	WX11344<= not TM1;
	WX11345<= not WX11344;
	WX11346<= not WX11342;
	WX11347<= not WX11343;
	WX11348<= not WX11341;
	WX11349<= not WX11340;
	WX11353<= not WX11349;
	WX11355<= not WX11354;
	WX11356<= not WX11355;
	WX11360<= not WX11349;
	WX11362<= not WX11361;
	WX11363<= not WX11362;
	WX11367<= not WX11349;
	WX11369<= not WX11368;
	WX11370<= not WX11369;
	WX11374<= not WX11349;
	WX11376<= not WX11375;
	WX11377<= not WX11376;
	WX11381<= not WX11349;
	WX11383<= not WX11382;
	WX11384<= not WX11383;
	WX11388<= not WX11349;
	WX11390<= not WX11389;
	WX11391<= not WX11390;
	WX11395<= not WX11349;
	WX11397<= not WX11396;
	WX11398<= not WX11397;
	WX11402<= not WX11349;
	WX11404<= not WX11403;
	WX11405<= not WX11404;
	WX11409<= not WX11349;
	WX11411<= not WX11410;
	WX11412<= not WX11411;
	WX11416<= not WX11349;
	WX11418<= not WX11417;
	WX11419<= not WX11418;
	WX11423<= not WX11349;
	WX11425<= not WX11424;
	WX11426<= not WX11425;
	WX11430<= not WX11349;
	WX11432<= not WX11431;
	WX11433<= not WX11432;
	WX11437<= not WX11349;
	WX11439<= not WX11438;
	WX11440<= not WX11439;
	WX11444<= not WX11349;
	WX11446<= not WX11445;
	WX11447<= not WX11446;
	WX11451<= not WX11349;
	WX11453<= not WX11452;
	WX11454<= not WX11453;
	WX11458<= not WX11349;
	WX11460<= not WX11459;
	WX11461<= not WX11460;
	WX11465<= not WX11349;
	WX11467<= not WX11466;
	WX11468<= not WX11467;
	WX11472<= not WX11349;
	WX11474<= not WX11473;
	WX11475<= not WX11474;
	WX11479<= not WX11349;
	WX11481<= not WX11480;
	WX11482<= not WX11481;
	WX11486<= not WX11349;
	WX11488<= not WX11487;
	WX11489<= not WX11488;
	WX11493<= not WX11349;
	WX11495<= not WX11494;
	WX11496<= not WX11495;
	WX11500<= not WX11349;
	WX11502<= not WX11501;
	WX11503<= not WX11502;
	WX11507<= not WX11349;
	WX11509<= not WX11508;
	WX11510<= not WX11509;
	WX11514<= not WX11349;
	WX11516<= not WX11515;
	WX11517<= not WX11516;
	WX11521<= not WX11349;
	WX11523<= not WX11522;
	WX11524<= not WX11523;
	WX11528<= not WX11349;
	WX11530<= not WX11529;
	WX11531<= not WX11530;
	WX11535<= not WX11349;
	WX11537<= not WX11536;
	WX11538<= not WX11537;
	WX11542<= not WX11349;
	WX11544<= not WX11543;
	WX11545<= not WX11544;
	WX11549<= not WX11349;
	WX11551<= not WX11550;
	WX11552<= not WX11551;
	WX11556<= not WX11349;
	WX11558<= not WX11557;
	WX11559<= not WX11558;
	WX11563<= not WX11349;
	WX11565<= not WX11564;
	WX11566<= not WX11565;
	WX11570<= not WX11349;
	WX11572<= not WX11571;
	WX11573<= not WX11572;
	WX11574<= not RESET;
	WX11607<= not WX11574;
	WX35<=WX46 and WX1003;
	WX36<=WX42 and WX37;
	WX39<=CRC_OUT_9_31 and WX1004;
	WX40<=WX2305 and WX41;
	WX43<=WX485 and WX1004;
	WX44<=DATA_9_31 and WX45;
	WX49<=WX60 and WX1003;
	WX50<=WX56 and WX51;
	WX53<=CRC_OUT_9_30 and WX1004;
	WX54<=WX2312 and WX55;
	WX57<=WX487 and WX1004;
	WX58<=DATA_9_30 and WX59;
	WX63<=WX74 and WX1003;
	WX64<=WX70 and WX65;
	WX67<=CRC_OUT_9_29 and WX1004;
	WX68<=WX2319 and WX69;
	WX71<=WX489 and WX1004;
	WX72<=DATA_9_29 and WX73;
	WX77<=WX88 and WX1003;
	WX78<=WX84 and WX79;
	WX81<=CRC_OUT_9_28 and WX1004;
	WX82<=WX2326 and WX83;
	WX85<=WX491 and WX1004;
	WX86<=DATA_9_28 and WX87;
	WX91<=WX102 and WX1003;
	WX92<=WX98 and WX93;
	WX95<=CRC_OUT_9_27 and WX1004;
	WX96<=WX2333 and WX97;
	WX99<=WX493 and WX1004;
	WX100<=DATA_9_27 and WX101;
	WX105<=WX116 and WX1003;
	WX106<=WX112 and WX107;
	WX109<=CRC_OUT_9_26 and WX1004;
	WX110<=WX2340 and WX111;
	WX113<=WX495 and WX1004;
	WX114<=DATA_9_26 and WX115;
	WX119<=WX130 and WX1003;
	WX120<=WX126 and WX121;
	WX123<=CRC_OUT_9_25 and WX1004;
	WX124<=WX2347 and WX125;
	WX127<=WX497 and WX1004;
	WX128<=DATA_9_25 and WX129;
	WX133<=WX144 and WX1003;
	WX134<=WX140 and WX135;
	WX137<=CRC_OUT_9_24 and WX1004;
	WX138<=WX2354 and WX139;
	WX141<=WX499 and WX1004;
	WX142<=DATA_9_24 and WX143;
	WX147<=WX158 and WX1003;
	WX148<=WX154 and WX149;
	WX151<=CRC_OUT_9_23 and WX1004;
	WX152<=WX2361 and WX153;
	WX155<=WX501 and WX1004;
	WX156<=DATA_9_23 and WX157;
	WX161<=WX172 and WX1003;
	WX162<=WX168 and WX163;
	WX165<=CRC_OUT_9_22 and WX1004;
	WX166<=WX2368 and WX167;
	WX169<=WX503 and WX1004;
	WX170<=DATA_9_22 and WX171;
	WX175<=WX186 and WX1003;
	WX176<=WX182 and WX177;
	WX179<=CRC_OUT_9_21 and WX1004;
	WX180<=WX2375 and WX181;
	WX183<=WX505 and WX1004;
	WX184<=DATA_9_21 and WX185;
	WX189<=WX200 and WX1003;
	WX190<=WX196 and WX191;
	WX193<=CRC_OUT_9_20 and WX1004;
	WX194<=WX2382 and WX195;
	WX197<=WX507 and WX1004;
	WX198<=DATA_9_20 and WX199;
	WX203<=WX214 and WX1003;
	WX204<=WX210 and WX205;
	WX207<=CRC_OUT_9_19 and WX1004;
	WX208<=WX2389 and WX209;
	WX211<=WX509 and WX1004;
	WX212<=DATA_9_19 and WX213;
	WX217<=WX228 and WX1003;
	WX218<=WX224 and WX219;
	WX221<=CRC_OUT_9_18 and WX1004;
	WX222<=WX2396 and WX223;
	WX225<=WX511 and WX1004;
	WX226<=DATA_9_18 and WX227;
	WX231<=WX242 and WX1003;
	WX232<=WX238 and WX233;
	WX235<=CRC_OUT_9_17 and WX1004;
	WX236<=WX2403 and WX237;
	WX239<=WX513 and WX1004;
	WX240<=DATA_9_17 and WX241;
	WX245<=WX256 and WX1003;
	WX246<=WX252 and WX247;
	WX249<=CRC_OUT_9_16 and WX1004;
	WX250<=WX2410 and WX251;
	WX253<=WX515 and WX1004;
	WX254<=DATA_9_16 and WX255;
	WX259<=WX270 and WX1003;
	WX260<=WX266 and WX261;
	WX263<=CRC_OUT_9_15 and WX1004;
	WX264<=WX2417 and WX265;
	WX267<=WX517 and WX1004;
	WX268<=DATA_9_15 and WX269;
	WX273<=WX284 and WX1003;
	WX274<=WX280 and WX275;
	WX277<=CRC_OUT_9_14 and WX1004;
	WX278<=WX2424 and WX279;
	WX281<=WX519 and WX1004;
	WX282<=DATA_9_14 and WX283;
	WX287<=WX298 and WX1003;
	WX288<=WX294 and WX289;
	WX291<=CRC_OUT_9_13 and WX1004;
	WX292<=WX2431 and WX293;
	WX295<=WX521 and WX1004;
	WX296<=DATA_9_13 and WX297;
	WX301<=WX312 and WX1003;
	WX302<=WX308 and WX303;
	WX305<=CRC_OUT_9_12 and WX1004;
	WX306<=WX2438 and WX307;
	WX309<=WX523 and WX1004;
	WX310<=DATA_9_12 and WX311;
	WX315<=WX326 and WX1003;
	WX316<=WX322 and WX317;
	WX319<=CRC_OUT_9_11 and WX1004;
	WX320<=WX2445 and WX321;
	WX323<=WX525 and WX1004;
	WX324<=DATA_9_11 and WX325;
	WX329<=WX340 and WX1003;
	WX330<=WX336 and WX331;
	WX333<=CRC_OUT_9_10 and WX1004;
	WX334<=WX2452 and WX335;
	WX337<=WX527 and WX1004;
	WX338<=DATA_9_10 and WX339;
	WX343<=WX354 and WX1003;
	WX344<=WX350 and WX345;
	WX347<=CRC_OUT_9_9 and WX1004;
	WX348<=WX2459 and WX349;
	WX351<=WX529 and WX1004;
	WX352<=DATA_9_9 and WX353;
	WX357<=WX368 and WX1003;
	WX358<=WX364 and WX359;
	WX361<=CRC_OUT_9_8 and WX1004;
	WX362<=WX2466 and WX363;
	WX365<=WX531 and WX1004;
	WX366<=DATA_9_8 and WX367;
	WX371<=WX382 and WX1003;
	WX372<=WX378 and WX373;
	WX375<=CRC_OUT_9_7 and WX1004;
	WX376<=WX2473 and WX377;
	WX379<=WX533 and WX1004;
	WX380<=DATA_9_7 and WX381;
	WX385<=WX396 and WX1003;
	WX386<=WX392 and WX387;
	WX389<=CRC_OUT_9_6 and WX1004;
	WX390<=WX2480 and WX391;
	WX393<=WX535 and WX1004;
	WX394<=DATA_9_6 and WX395;
	WX399<=WX410 and WX1003;
	WX400<=WX406 and WX401;
	WX403<=CRC_OUT_9_5 and WX1004;
	WX404<=WX2487 and WX405;
	WX407<=WX537 and WX1004;
	WX408<=DATA_9_5 and WX409;
	WX413<=WX424 and WX1003;
	WX414<=WX420 and WX415;
	WX417<=CRC_OUT_9_4 and WX1004;
	WX418<=WX2494 and WX419;
	WX421<=WX539 and WX1004;
	WX422<=DATA_9_4 and WX423;
	WX427<=WX438 and WX1003;
	WX428<=WX434 and WX429;
	WX431<=CRC_OUT_9_3 and WX1004;
	WX432<=WX2501 and WX433;
	WX435<=WX541 and WX1004;
	WX436<=DATA_9_3 and WX437;
	WX441<=WX452 and WX1003;
	WX442<=WX448 and WX443;
	WX445<=CRC_OUT_9_2 and WX1004;
	WX446<=WX2508 and WX447;
	WX449<=WX543 and WX1004;
	WX450<=DATA_9_2 and WX451;
	WX455<=WX466 and WX1003;
	WX456<=WX462 and WX457;
	WX459<=CRC_OUT_9_1 and WX1004;
	WX460<=WX2515 and WX461;
	WX463<=WX545 and WX1004;
	WX464<=DATA_9_1 and WX465;
	WX469<=WX480 and WX1003;
	WX470<=WX476 and WX471;
	WX473<=CRC_OUT_9_0 and WX1004;
	WX474<=WX2522 and WX475;
	WX477<=WX547 and WX1004;
	WX478<=DATA_9_0 and WX479;
	WX484<=WX487 and RESET;
	WX486<=WX489 and RESET;
	WX488<=WX491 and RESET;
	WX490<=WX493 and RESET;
	WX492<=WX495 and RESET;
	WX494<=WX497 and RESET;
	WX496<=WX499 and RESET;
	WX498<=WX501 and RESET;
	WX500<=WX503 and RESET;
	WX502<=WX505 and RESET;
	WX504<=WX507 and RESET;
	WX506<=WX509 and RESET;
	WX508<=WX511 and RESET;
	WX510<=WX513 and RESET;
	WX512<=WX515 and RESET;
	WX514<=WX517 and RESET;
	WX516<=WX519 and RESET;
	WX518<=WX521 and RESET;
	WX520<=WX523 and RESET;
	WX522<=WX525 and RESET;
	WX524<=WX527 and RESET;
	WX526<=WX529 and RESET;
	WX528<=WX531 and RESET;
	WX530<=WX533 and RESET;
	WX532<=WX535 and RESET;
	WX534<=WX537 and RESET;
	WX536<=WX539 and RESET;
	WX538<=WX541 and RESET;
	WX540<=WX543 and RESET;
	WX542<=WX545 and RESET;
	WX544<=WX547 and RESET;
	WX546<=WX483 and RESET;
	WX644<=WX48 and RESET;
	WX646<=WX62 and RESET;
	WX648<=WX76 and RESET;
	WX650<=WX90 and RESET;
	WX652<=WX104 and RESET;
	WX654<=WX118 and RESET;
	WX656<=WX132 and RESET;
	WX658<=WX146 and RESET;
	WX660<=WX160 and RESET;
	WX662<=WX174 and RESET;
	WX664<=WX188 and RESET;
	WX666<=WX202 and RESET;
	WX668<=WX216 and RESET;
	WX670<=WX230 and RESET;
	WX672<=WX244 and RESET;
	WX674<=WX258 and RESET;
	WX676<=WX272 and RESET;
	WX678<=WX286 and RESET;
	WX680<=WX300 and RESET;
	WX682<=WX314 and RESET;
	WX684<=WX328 and RESET;
	WX686<=WX342 and RESET;
	WX688<=WX356 and RESET;
	WX690<=WX370 and RESET;
	WX692<=WX384 and RESET;
	WX694<=WX398 and RESET;
	WX696<=WX412 and RESET;
	WX698<=WX426 and RESET;
	WX700<=WX440 and RESET;
	WX702<=WX454 and RESET;
	WX704<=WX468 and RESET;
	WX706<=WX482 and RESET;
	WX708<=WX645 and RESET;
	WX710<=WX647 and RESET;
	WX712<=WX649 and RESET;
	WX714<=WX651 and RESET;
	WX716<=WX653 and RESET;
	WX718<=WX655 and RESET;
	WX720<=WX657 and RESET;
	WX722<=WX659 and RESET;
	WX724<=WX661 and RESET;
	WX726<=WX663 and RESET;
	WX728<=WX665 and RESET;
	WX730<=WX667 and RESET;
	WX732<=WX669 and RESET;
	WX734<=WX671 and RESET;
	WX736<=WX673 and RESET;
	WX738<=WX675 and RESET;
	WX740<=WX677 and RESET;
	WX742<=WX679 and RESET;
	WX744<=WX681 and RESET;
	WX746<=WX683 and RESET;
	WX748<=WX685 and RESET;
	WX750<=WX687 and RESET;
	WX752<=WX689 and RESET;
	WX754<=WX691 and RESET;
	WX756<=WX693 and RESET;
	WX758<=WX695 and RESET;
	WX760<=WX697 and RESET;
	WX762<=WX699 and RESET;
	WX764<=WX701 and RESET;
	WX766<=WX703 and RESET;
	WX768<=WX705 and RESET;
	WX770<=WX707 and RESET;
	WX772<=WX709 and RESET;
	WX774<=WX711 and RESET;
	WX776<=WX713 and RESET;
	WX778<=WX715 and RESET;
	WX780<=WX717 and RESET;
	WX782<=WX719 and RESET;
	WX784<=WX721 and RESET;
	WX786<=WX723 and RESET;
	WX788<=WX725 and RESET;
	WX790<=WX727 and RESET;
	WX792<=WX729 and RESET;
	WX794<=WX731 and RESET;
	WX796<=WX733 and RESET;
	WX798<=WX735 and RESET;
	WX800<=WX737 and RESET;
	WX802<=WX739 and RESET;
	WX804<=WX741 and RESET;
	WX806<=WX743 and RESET;
	WX808<=WX745 and RESET;
	WX810<=WX747 and RESET;
	WX812<=WX749 and RESET;
	WX814<=WX751 and RESET;
	WX816<=WX753 and RESET;
	WX818<=WX755 and RESET;
	WX820<=WX757 and RESET;
	WX822<=WX759 and RESET;
	WX824<=WX761 and RESET;
	WX826<=WX763 and RESET;
	WX828<=WX765 and RESET;
	WX830<=WX767 and RESET;
	WX832<=WX769 and RESET;
	WX834<=WX771 and RESET;
	WX836<=WX773 and RESET;
	WX838<=WX775 and RESET;
	WX840<=WX777 and RESET;
	WX842<=WX779 and RESET;
	WX844<=WX781 and RESET;
	WX846<=WX783 and RESET;
	WX848<=WX785 and RESET;
	WX850<=WX787 and RESET;
	WX852<=WX789 and RESET;
	WX854<=WX791 and RESET;
	WX856<=WX793 and RESET;
	WX858<=WX795 and RESET;
	WX860<=WX797 and RESET;
	WX862<=WX799 and RESET;
	WX864<=WX801 and RESET;
	WX866<=WX803 and RESET;
	WX868<=WX805 and RESET;
	WX870<=WX807 and RESET;
	WX872<=WX809 and RESET;
	WX874<=WX811 and RESET;
	WX876<=WX813 and RESET;
	WX878<=WX815 and RESET;
	WX880<=WX817 and RESET;
	WX882<=WX819 and RESET;
	WX884<=WX821 and RESET;
	WX886<=WX823 and RESET;
	WX888<=WX825 and RESET;
	WX890<=WX827 and RESET;
	WX892<=WX829 and RESET;
	WX894<=WX831 and RESET;
	WX896<=WX833 and RESET;
	WX898<=WX835 and RESET;
	WX1007<=WX1006 and WX1005;
	WX1008<=WX580 and WX1009;
	WX1014<=WX1013 and WX1005;
	WX1015<=WX581 and WX1016;
	WX1021<=WX1020 and WX1005;
	WX1022<=WX582 and WX1023;
	WX1028<=WX1027 and WX1005;
	WX1029<=WX583 and WX1030;
	WX1035<=WX1034 and WX1005;
	WX1036<=WX584 and WX1037;
	WX1042<=WX1041 and WX1005;
	WX1043<=WX585 and WX1044;
	WX1049<=WX1048 and WX1005;
	WX1050<=WX586 and WX1051;
	WX1056<=WX1055 and WX1005;
	WX1057<=WX587 and WX1058;
	WX1063<=WX1062 and WX1005;
	WX1064<=WX588 and WX1065;
	WX1070<=WX1069 and WX1005;
	WX1071<=WX589 and WX1072;
	WX1077<=WX1076 and WX1005;
	WX1078<=WX590 and WX1079;
	WX1084<=WX1083 and WX1005;
	WX1085<=WX591 and WX1086;
	WX1091<=WX1090 and WX1005;
	WX1092<=WX592 and WX1093;
	WX1098<=WX1097 and WX1005;
	WX1099<=WX593 and WX1100;
	WX1105<=WX1104 and WX1005;
	WX1106<=WX594 and WX1107;
	WX1112<=WX1111 and WX1005;
	WX1113<=WX595 and WX1114;
	WX1119<=WX1118 and WX1005;
	WX1120<=WX596 and WX1121;
	WX1126<=WX1125 and WX1005;
	WX1127<=WX597 and WX1128;
	WX1133<=WX1132 and WX1005;
	WX1134<=WX598 and WX1135;
	WX1140<=WX1139 and WX1005;
	WX1141<=WX599 and WX1142;
	WX1147<=WX1146 and WX1005;
	WX1148<=WX600 and WX1149;
	WX1154<=WX1153 and WX1005;
	WX1155<=WX601 and WX1156;
	WX1161<=WX1160 and WX1005;
	WX1162<=WX602 and WX1163;
	WX1168<=WX1167 and WX1005;
	WX1169<=WX603 and WX1170;
	WX1175<=WX1174 and WX1005;
	WX1176<=WX604 and WX1177;
	WX1182<=WX1181 and WX1005;
	WX1183<=WX605 and WX1184;
	WX1189<=WX1188 and WX1005;
	WX1190<=WX606 and WX1191;
	WX1196<=WX1195 and WX1005;
	WX1197<=WX607 and WX1198;
	WX1203<=WX1202 and WX1005;
	WX1204<=WX608 and WX1205;
	WX1210<=WX1209 and WX1005;
	WX1211<=WX609 and WX1212;
	WX1217<=WX1216 and WX1005;
	WX1218<=WX610 and WX1219;
	WX1224<=WX1223 and WX1005;
	WX1225<=WX611 and WX1226;
	WX1264<=WX1234 and WX1263;
	WX1266<=WX1262 and WX1263;
	WX1268<=WX1261 and WX1263;
	WX1270<=WX1260 and WX1263;
	WX1272<=WX1233 and WX1263;
	WX1274<=WX1259 and WX1263;
	WX1276<=WX1258 and WX1263;
	WX1278<=WX1257 and WX1263;
	WX1280<=WX1256 and WX1263;
	WX1282<=WX1255 and WX1263;
	WX1284<=WX1254 and WX1263;
	WX1286<=WX1232 and WX1263;
	WX1288<=WX1253 and WX1263;
	WX1290<=WX1252 and WX1263;
	WX1292<=WX1251 and WX1263;
	WX1294<=WX1250 and WX1263;
	WX1296<=WX1231 and WX1263;
	WX1298<=WX1249 and WX1263;
	WX1300<=WX1248 and WX1263;
	WX1302<=WX1247 and WX1263;
	WX1304<=WX1246 and WX1263;
	WX1306<=WX1245 and WX1263;
	WX1308<=WX1244 and WX1263;
	WX1310<=WX1243 and WX1263;
	WX1312<=WX1242 and WX1263;
	WX1314<=WX1241 and WX1263;
	WX1316<=WX1240 and WX1263;
	WX1318<=WX1239 and WX1263;
	WX1320<=WX1238 and WX1263;
	WX1322<=WX1237 and WX1263;
	WX1324<=WX1236 and WX1263;
	WX1326<=WX1235 and WX1263;
	WX1328<=WX1339 and WX2296;
	WX1329<=WX1335 and WX1330;
	WX1332<=CRC_OUT_8_31 and WX2297;
	WX1333<=WX3598 and WX1334;
	WX1336<=WX1778 and WX2297;
	WX1337<=WX2305 and WX1338;
	WX1342<=WX1353 and WX2296;
	WX1343<=WX1349 and WX1344;
	WX1346<=CRC_OUT_8_30 and WX2297;
	WX1347<=WX3605 and WX1348;
	WX1350<=WX1780 and WX2297;
	WX1351<=WX2312 and WX1352;
	WX1356<=WX1367 and WX2296;
	WX1357<=WX1363 and WX1358;
	WX1360<=CRC_OUT_8_29 and WX2297;
	WX1361<=WX3612 and WX1362;
	WX1364<=WX1782 and WX2297;
	WX1365<=WX2319 and WX1366;
	WX1370<=WX1381 and WX2296;
	WX1371<=WX1377 and WX1372;
	WX1374<=CRC_OUT_8_28 and WX2297;
	WX1375<=WX3619 and WX1376;
	WX1378<=WX1784 and WX2297;
	WX1379<=WX2326 and WX1380;
	WX1384<=WX1395 and WX2296;
	WX1385<=WX1391 and WX1386;
	WX1388<=CRC_OUT_8_27 and WX2297;
	WX1389<=WX3626 and WX1390;
	WX1392<=WX1786 and WX2297;
	WX1393<=WX2333 and WX1394;
	WX1398<=WX1409 and WX2296;
	WX1399<=WX1405 and WX1400;
	WX1402<=CRC_OUT_8_26 and WX2297;
	WX1403<=WX3633 and WX1404;
	WX1406<=WX1788 and WX2297;
	WX1407<=WX2340 and WX1408;
	WX1412<=WX1423 and WX2296;
	WX1413<=WX1419 and WX1414;
	WX1416<=CRC_OUT_8_25 and WX2297;
	WX1417<=WX3640 and WX1418;
	WX1420<=WX1790 and WX2297;
	WX1421<=WX2347 and WX1422;
	WX1426<=WX1437 and WX2296;
	WX1427<=WX1433 and WX1428;
	WX1430<=CRC_OUT_8_24 and WX2297;
	WX1431<=WX3647 and WX1432;
	WX1434<=WX1792 and WX2297;
	WX1435<=WX2354 and WX1436;
	WX1440<=WX1451 and WX2296;
	WX1441<=WX1447 and WX1442;
	WX1444<=CRC_OUT_8_23 and WX2297;
	WX1445<=WX3654 and WX1446;
	WX1448<=WX1794 and WX2297;
	WX1449<=WX2361 and WX1450;
	WX1454<=WX1465 and WX2296;
	WX1455<=WX1461 and WX1456;
	WX1458<=CRC_OUT_8_22 and WX2297;
	WX1459<=WX3661 and WX1460;
	WX1462<=WX1796 and WX2297;
	WX1463<=WX2368 and WX1464;
	WX1468<=WX1479 and WX2296;
	WX1469<=WX1475 and WX1470;
	WX1472<=CRC_OUT_8_21 and WX2297;
	WX1473<=WX3668 and WX1474;
	WX1476<=WX1798 and WX2297;
	WX1477<=WX2375 and WX1478;
	WX1482<=WX1493 and WX2296;
	WX1483<=WX1489 and WX1484;
	WX1486<=CRC_OUT_8_20 and WX2297;
	WX1487<=WX3675 and WX1488;
	WX1490<=WX1800 and WX2297;
	WX1491<=WX2382 and WX1492;
	WX1496<=WX1507 and WX2296;
	WX1497<=WX1503 and WX1498;
	WX1500<=CRC_OUT_8_19 and WX2297;
	WX1501<=WX3682 and WX1502;
	WX1504<=WX1802 and WX2297;
	WX1505<=WX2389 and WX1506;
	WX1510<=WX1521 and WX2296;
	WX1511<=WX1517 and WX1512;
	WX1514<=CRC_OUT_8_18 and WX2297;
	WX1515<=WX3689 and WX1516;
	WX1518<=WX1804 and WX2297;
	WX1519<=WX2396 and WX1520;
	WX1524<=WX1535 and WX2296;
	WX1525<=WX1531 and WX1526;
	WX1528<=CRC_OUT_8_17 and WX2297;
	WX1529<=WX3696 and WX1530;
	WX1532<=WX1806 and WX2297;
	WX1533<=WX2403 and WX1534;
	WX1538<=WX1549 and WX2296;
	WX1539<=WX1545 and WX1540;
	WX1542<=CRC_OUT_8_16 and WX2297;
	WX1543<=WX3703 and WX1544;
	WX1546<=WX1808 and WX2297;
	WX1547<=WX2410 and WX1548;
	WX1552<=WX1563 and WX2296;
	WX1553<=WX1559 and WX1554;
	WX1556<=CRC_OUT_8_15 and WX2297;
	WX1557<=WX3710 and WX1558;
	WX1560<=WX1810 and WX2297;
	WX1561<=WX2417 and WX1562;
	WX1566<=WX1577 and WX2296;
	WX1567<=WX1573 and WX1568;
	WX1570<=CRC_OUT_8_14 and WX2297;
	WX1571<=WX3717 and WX1572;
	WX1574<=WX1812 and WX2297;
	WX1575<=WX2424 and WX1576;
	WX1580<=WX1591 and WX2296;
	WX1581<=WX1587 and WX1582;
	WX1584<=CRC_OUT_8_13 and WX2297;
	WX1585<=WX3724 and WX1586;
	WX1588<=WX1814 and WX2297;
	WX1589<=WX2431 and WX1590;
	WX1594<=WX1605 and WX2296;
	WX1595<=WX1601 and WX1596;
	WX1598<=CRC_OUT_8_12 and WX2297;
	WX1599<=WX3731 and WX1600;
	WX1602<=WX1816 and WX2297;
	WX1603<=WX2438 and WX1604;
	WX1608<=WX1619 and WX2296;
	WX1609<=WX1615 and WX1610;
	WX1612<=CRC_OUT_8_11 and WX2297;
	WX1613<=WX3738 and WX1614;
	WX1616<=WX1818 and WX2297;
	WX1617<=WX2445 and WX1618;
	WX1622<=WX1633 and WX2296;
	WX1623<=WX1629 and WX1624;
	WX1626<=CRC_OUT_8_10 and WX2297;
	WX1627<=WX3745 and WX1628;
	WX1630<=WX1820 and WX2297;
	WX1631<=WX2452 and WX1632;
	WX1636<=WX1647 and WX2296;
	WX1637<=WX1643 and WX1638;
	WX1640<=CRC_OUT_8_9 and WX2297;
	WX1641<=WX3752 and WX1642;
	WX1644<=WX1822 and WX2297;
	WX1645<=WX2459 and WX1646;
	WX1650<=WX1661 and WX2296;
	WX1651<=WX1657 and WX1652;
	WX1654<=CRC_OUT_8_8 and WX2297;
	WX1655<=WX3759 and WX1656;
	WX1658<=WX1824 and WX2297;
	WX1659<=WX2466 and WX1660;
	WX1664<=WX1675 and WX2296;
	WX1665<=WX1671 and WX1666;
	WX1668<=CRC_OUT_8_7 and WX2297;
	WX1669<=WX3766 and WX1670;
	WX1672<=WX1826 and WX2297;
	WX1673<=WX2473 and WX1674;
	WX1678<=WX1689 and WX2296;
	WX1679<=WX1685 and WX1680;
	WX1682<=CRC_OUT_8_6 and WX2297;
	WX1683<=WX3773 and WX1684;
	WX1686<=WX1828 and WX2297;
	WX1687<=WX2480 and WX1688;
	WX1692<=WX1703 and WX2296;
	WX1693<=WX1699 and WX1694;
	WX1696<=CRC_OUT_8_5 and WX2297;
	WX1697<=WX3780 and WX1698;
	WX1700<=WX1830 and WX2297;
	WX1701<=WX2487 and WX1702;
	WX1706<=WX1717 and WX2296;
	WX1707<=WX1713 and WX1708;
	WX1710<=CRC_OUT_8_4 and WX2297;
	WX1711<=WX3787 and WX1712;
	WX1714<=WX1832 and WX2297;
	WX1715<=WX2494 and WX1716;
	WX1720<=WX1731 and WX2296;
	WX1721<=WX1727 and WX1722;
	WX1724<=CRC_OUT_8_3 and WX2297;
	WX1725<=WX3794 and WX1726;
	WX1728<=WX1834 and WX2297;
	WX1729<=WX2501 and WX1730;
	WX1734<=WX1745 and WX2296;
	WX1735<=WX1741 and WX1736;
	WX1738<=CRC_OUT_8_2 and WX2297;
	WX1739<=WX3801 and WX1740;
	WX1742<=WX1836 and WX2297;
	WX1743<=WX2508 and WX1744;
	WX1748<=WX1759 and WX2296;
	WX1749<=WX1755 and WX1750;
	WX1752<=CRC_OUT_8_1 and WX2297;
	WX1753<=WX3808 and WX1754;
	WX1756<=WX1838 and WX2297;
	WX1757<=WX2515 and WX1758;
	WX1762<=WX1773 and WX2296;
	WX1763<=WX1769 and WX1764;
	WX1766<=CRC_OUT_8_0 and WX2297;
	WX1767<=WX3815 and WX1768;
	WX1770<=WX1840 and WX2297;
	WX1771<=WX2522 and WX1772;
	WX1777<=WX1780 and RESET;
	WX1779<=WX1782 and RESET;
	WX1781<=WX1784 and RESET;
	WX1783<=WX1786 and RESET;
	WX1785<=WX1788 and RESET;
	WX1787<=WX1790 and RESET;
	WX1789<=WX1792 and RESET;
	WX1791<=WX1794 and RESET;
	WX1793<=WX1796 and RESET;
	WX1795<=WX1798 and RESET;
	WX1797<=WX1800 and RESET;
	WX1799<=WX1802 and RESET;
	WX1801<=WX1804 and RESET;
	WX1803<=WX1806 and RESET;
	WX1805<=WX1808 and RESET;
	WX1807<=WX1810 and RESET;
	WX1809<=WX1812 and RESET;
	WX1811<=WX1814 and RESET;
	WX1813<=WX1816 and RESET;
	WX1815<=WX1818 and RESET;
	WX1817<=WX1820 and RESET;
	WX1819<=WX1822 and RESET;
	WX1821<=WX1824 and RESET;
	WX1823<=WX1826 and RESET;
	WX1825<=WX1828 and RESET;
	WX1827<=WX1830 and RESET;
	WX1829<=WX1832 and RESET;
	WX1831<=WX1834 and RESET;
	WX1833<=WX1836 and RESET;
	WX1835<=WX1838 and RESET;
	WX1837<=WX1840 and RESET;
	WX1839<=WX1776 and RESET;
	WX1937<=WX1341 and RESET;
	WX1939<=WX1355 and RESET;
	WX1941<=WX1369 and RESET;
	WX1943<=WX1383 and RESET;
	WX1945<=WX1397 and RESET;
	WX1947<=WX1411 and RESET;
	WX1949<=WX1425 and RESET;
	WX1951<=WX1439 and RESET;
	WX1953<=WX1453 and RESET;
	WX1955<=WX1467 and RESET;
	WX1957<=WX1481 and RESET;
	WX1959<=WX1495 and RESET;
	WX1961<=WX1509 and RESET;
	WX1963<=WX1523 and RESET;
	WX1965<=WX1537 and RESET;
	WX1967<=WX1551 and RESET;
	WX1969<=WX1565 and RESET;
	WX1971<=WX1579 and RESET;
	WX1973<=WX1593 and RESET;
	WX1975<=WX1607 and RESET;
	WX1977<=WX1621 and RESET;
	WX1979<=WX1635 and RESET;
	WX1981<=WX1649 and RESET;
	WX1983<=WX1663 and RESET;
	WX1985<=WX1677 and RESET;
	WX1987<=WX1691 and RESET;
	WX1989<=WX1705 and RESET;
	WX1991<=WX1719 and RESET;
	WX1993<=WX1733 and RESET;
	WX1995<=WX1747 and RESET;
	WX1997<=WX1761 and RESET;
	WX1999<=WX1775 and RESET;
	WX2001<=WX1938 and RESET;
	WX2003<=WX1940 and RESET;
	WX2005<=WX1942 and RESET;
	WX2007<=WX1944 and RESET;
	WX2009<=WX1946 and RESET;
	WX2011<=WX1948 and RESET;
	WX2013<=WX1950 and RESET;
	WX2015<=WX1952 and RESET;
	WX2017<=WX1954 and RESET;
	WX2019<=WX1956 and RESET;
	WX2021<=WX1958 and RESET;
	WX2023<=WX1960 and RESET;
	WX2025<=WX1962 and RESET;
	WX2027<=WX1964 and RESET;
	WX2029<=WX1966 and RESET;
	WX2031<=WX1968 and RESET;
	WX2033<=WX1970 and RESET;
	WX2035<=WX1972 and RESET;
	WX2037<=WX1974 and RESET;
	WX2039<=WX1976 and RESET;
	WX2041<=WX1978 and RESET;
	WX2043<=WX1980 and RESET;
	WX2045<=WX1982 and RESET;
	WX2047<=WX1984 and RESET;
	WX2049<=WX1986 and RESET;
	WX2051<=WX1988 and RESET;
	WX2053<=WX1990 and RESET;
	WX2055<=WX1992 and RESET;
	WX2057<=WX1994 and RESET;
	WX2059<=WX1996 and RESET;
	WX2061<=WX1998 and RESET;
	WX2063<=WX2000 and RESET;
	WX2065<=WX2002 and RESET;
	WX2067<=WX2004 and RESET;
	WX2069<=WX2006 and RESET;
	WX2071<=WX2008 and RESET;
	WX2073<=WX2010 and RESET;
	WX2075<=WX2012 and RESET;
	WX2077<=WX2014 and RESET;
	WX2079<=WX2016 and RESET;
	WX2081<=WX2018 and RESET;
	WX2083<=WX2020 and RESET;
	WX2085<=WX2022 and RESET;
	WX2087<=WX2024 and RESET;
	WX2089<=WX2026 and RESET;
	WX2091<=WX2028 and RESET;
	WX2093<=WX2030 and RESET;
	WX2095<=WX2032 and RESET;
	WX2097<=WX2034 and RESET;
	WX2099<=WX2036 and RESET;
	WX2101<=WX2038 and RESET;
	WX2103<=WX2040 and RESET;
	WX2105<=WX2042 and RESET;
	WX2107<=WX2044 and RESET;
	WX2109<=WX2046 and RESET;
	WX2111<=WX2048 and RESET;
	WX2113<=WX2050 and RESET;
	WX2115<=WX2052 and RESET;
	WX2117<=WX2054 and RESET;
	WX2119<=WX2056 and RESET;
	WX2121<=WX2058 and RESET;
	WX2123<=WX2060 and RESET;
	WX2125<=WX2062 and RESET;
	WX2127<=WX2064 and RESET;
	WX2129<=WX2066 and RESET;
	WX2131<=WX2068 and RESET;
	WX2133<=WX2070 and RESET;
	WX2135<=WX2072 and RESET;
	WX2137<=WX2074 and RESET;
	WX2139<=WX2076 and RESET;
	WX2141<=WX2078 and RESET;
	WX2143<=WX2080 and RESET;
	WX2145<=WX2082 and RESET;
	WX2147<=WX2084 and RESET;
	WX2149<=WX2086 and RESET;
	WX2151<=WX2088 and RESET;
	WX2153<=WX2090 and RESET;
	WX2155<=WX2092 and RESET;
	WX2157<=WX2094 and RESET;
	WX2159<=WX2096 and RESET;
	WX2161<=WX2098 and RESET;
	WX2163<=WX2100 and RESET;
	WX2165<=WX2102 and RESET;
	WX2167<=WX2104 and RESET;
	WX2169<=WX2106 and RESET;
	WX2171<=WX2108 and RESET;
	WX2173<=WX2110 and RESET;
	WX2175<=WX2112 and RESET;
	WX2177<=WX2114 and RESET;
	WX2179<=WX2116 and RESET;
	WX2181<=WX2118 and RESET;
	WX2183<=WX2120 and RESET;
	WX2185<=WX2122 and RESET;
	WX2187<=WX2124 and RESET;
	WX2189<=WX2126 and RESET;
	WX2191<=WX2128 and RESET;
	WX2300<=WX2299 and WX2298;
	WX2301<=WX1873 and WX2302;
	WX2307<=WX2306 and WX2298;
	WX2308<=WX1874 and WX2309;
	WX2314<=WX2313 and WX2298;
	WX2315<=WX1875 and WX2316;
	WX2321<=WX2320 and WX2298;
	WX2322<=WX1876 and WX2323;
	WX2328<=WX2327 and WX2298;
	WX2329<=WX1877 and WX2330;
	WX2335<=WX2334 and WX2298;
	WX2336<=WX1878 and WX2337;
	WX2342<=WX2341 and WX2298;
	WX2343<=WX1879 and WX2344;
	WX2349<=WX2348 and WX2298;
	WX2350<=WX1880 and WX2351;
	WX2356<=WX2355 and WX2298;
	WX2357<=WX1881 and WX2358;
	WX2363<=WX2362 and WX2298;
	WX2364<=WX1882 and WX2365;
	WX2370<=WX2369 and WX2298;
	WX2371<=WX1883 and WX2372;
	WX2377<=WX2376 and WX2298;
	WX2378<=WX1884 and WX2379;
	WX2384<=WX2383 and WX2298;
	WX2385<=WX1885 and WX2386;
	WX2391<=WX2390 and WX2298;
	WX2392<=WX1886 and WX2393;
	WX2398<=WX2397 and WX2298;
	WX2399<=WX1887 and WX2400;
	WX2405<=WX2404 and WX2298;
	WX2406<=WX1888 and WX2407;
	WX2412<=WX2411 and WX2298;
	WX2413<=WX1889 and WX2414;
	WX2419<=WX2418 and WX2298;
	WX2420<=WX1890 and WX2421;
	WX2426<=WX2425 and WX2298;
	WX2427<=WX1891 and WX2428;
	WX2433<=WX2432 and WX2298;
	WX2434<=WX1892 and WX2435;
	WX2440<=WX2439 and WX2298;
	WX2441<=WX1893 and WX2442;
	WX2447<=WX2446 and WX2298;
	WX2448<=WX1894 and WX2449;
	WX2454<=WX2453 and WX2298;
	WX2455<=WX1895 and WX2456;
	WX2461<=WX2460 and WX2298;
	WX2462<=WX1896 and WX2463;
	WX2468<=WX2467 and WX2298;
	WX2469<=WX1897 and WX2470;
	WX2475<=WX2474 and WX2298;
	WX2476<=WX1898 and WX2477;
	WX2482<=WX2481 and WX2298;
	WX2483<=WX1899 and WX2484;
	WX2489<=WX2488 and WX2298;
	WX2490<=WX1900 and WX2491;
	WX2496<=WX2495 and WX2298;
	WX2497<=WX1901 and WX2498;
	WX2503<=WX2502 and WX2298;
	WX2504<=WX1902 and WX2505;
	WX2510<=WX2509 and WX2298;
	WX2511<=WX1903 and WX2512;
	WX2517<=WX2516 and WX2298;
	WX2518<=WX1904 and WX2519;
	WX2557<=WX2527 and WX2556;
	WX2559<=WX2555 and WX2556;
	WX2561<=WX2554 and WX2556;
	WX2563<=WX2553 and WX2556;
	WX2565<=WX2526 and WX2556;
	WX2567<=WX2552 and WX2556;
	WX2569<=WX2551 and WX2556;
	WX2571<=WX2550 and WX2556;
	WX2573<=WX2549 and WX2556;
	WX2575<=WX2548 and WX2556;
	WX2577<=WX2547 and WX2556;
	WX2579<=WX2525 and WX2556;
	WX2581<=WX2546 and WX2556;
	WX2583<=WX2545 and WX2556;
	WX2585<=WX2544 and WX2556;
	WX2587<=WX2543 and WX2556;
	WX2589<=WX2524 and WX2556;
	WX2591<=WX2542 and WX2556;
	WX2593<=WX2541 and WX2556;
	WX2595<=WX2540 and WX2556;
	WX2597<=WX2539 and WX2556;
	WX2599<=WX2538 and WX2556;
	WX2601<=WX2537 and WX2556;
	WX2603<=WX2536 and WX2556;
	WX2605<=WX2535 and WX2556;
	WX2607<=WX2534 and WX2556;
	WX2609<=WX2533 and WX2556;
	WX2611<=WX2532 and WX2556;
	WX2613<=WX2531 and WX2556;
	WX2615<=WX2530 and WX2556;
	WX2617<=WX2529 and WX2556;
	WX2619<=WX2528 and WX2556;
	WX2621<=WX2632 and WX3589;
	WX2622<=WX2628 and WX2623;
	WX2625<=CRC_OUT_7_31 and WX3590;
	WX2626<=WX4891 and WX2627;
	WX2629<=WX3071 and WX3590;
	WX2630<=WX3598 and WX2631;
	WX2635<=WX2646 and WX3589;
	WX2636<=WX2642 and WX2637;
	WX2639<=CRC_OUT_7_30 and WX3590;
	WX2640<=WX4898 and WX2641;
	WX2643<=WX3073 and WX3590;
	WX2644<=WX3605 and WX2645;
	WX2649<=WX2660 and WX3589;
	WX2650<=WX2656 and WX2651;
	WX2653<=CRC_OUT_7_29 and WX3590;
	WX2654<=WX4905 and WX2655;
	WX2657<=WX3075 and WX3590;
	WX2658<=WX3612 and WX2659;
	WX2663<=WX2674 and WX3589;
	WX2664<=WX2670 and WX2665;
	WX2667<=CRC_OUT_7_28 and WX3590;
	WX2668<=WX4912 and WX2669;
	WX2671<=WX3077 and WX3590;
	WX2672<=WX3619 and WX2673;
	WX2677<=WX2688 and WX3589;
	WX2678<=WX2684 and WX2679;
	WX2681<=CRC_OUT_7_27 and WX3590;
	WX2682<=WX4919 and WX2683;
	WX2685<=WX3079 and WX3590;
	WX2686<=WX3626 and WX2687;
	WX2691<=WX2702 and WX3589;
	WX2692<=WX2698 and WX2693;
	WX2695<=CRC_OUT_7_26 and WX3590;
	WX2696<=WX4926 and WX2697;
	WX2699<=WX3081 and WX3590;
	WX2700<=WX3633 and WX2701;
	WX2705<=WX2716 and WX3589;
	WX2706<=WX2712 and WX2707;
	WX2709<=CRC_OUT_7_25 and WX3590;
	WX2710<=WX4933 and WX2711;
	WX2713<=WX3083 and WX3590;
	WX2714<=WX3640 and WX2715;
	WX2719<=WX2730 and WX3589;
	WX2720<=WX2726 and WX2721;
	WX2723<=CRC_OUT_7_24 and WX3590;
	WX2724<=WX4940 and WX2725;
	WX2727<=WX3085 and WX3590;
	WX2728<=WX3647 and WX2729;
	WX2733<=WX2744 and WX3589;
	WX2734<=WX2740 and WX2735;
	WX2737<=CRC_OUT_7_23 and WX3590;
	WX2738<=WX4947 and WX2739;
	WX2741<=WX3087 and WX3590;
	WX2742<=WX3654 and WX2743;
	WX2747<=WX2758 and WX3589;
	WX2748<=WX2754 and WX2749;
	WX2751<=CRC_OUT_7_22 and WX3590;
	WX2752<=WX4954 and WX2753;
	WX2755<=WX3089 and WX3590;
	WX2756<=WX3661 and WX2757;
	WX2761<=WX2772 and WX3589;
	WX2762<=WX2768 and WX2763;
	WX2765<=CRC_OUT_7_21 and WX3590;
	WX2766<=WX4961 and WX2767;
	WX2769<=WX3091 and WX3590;
	WX2770<=WX3668 and WX2771;
	WX2775<=WX2786 and WX3589;
	WX2776<=WX2782 and WX2777;
	WX2779<=CRC_OUT_7_20 and WX3590;
	WX2780<=WX4968 and WX2781;
	WX2783<=WX3093 and WX3590;
	WX2784<=WX3675 and WX2785;
	WX2789<=WX2800 and WX3589;
	WX2790<=WX2796 and WX2791;
	WX2793<=CRC_OUT_7_19 and WX3590;
	WX2794<=WX4975 and WX2795;
	WX2797<=WX3095 and WX3590;
	WX2798<=WX3682 and WX2799;
	WX2803<=WX2814 and WX3589;
	WX2804<=WX2810 and WX2805;
	WX2807<=CRC_OUT_7_18 and WX3590;
	WX2808<=WX4982 and WX2809;
	WX2811<=WX3097 and WX3590;
	WX2812<=WX3689 and WX2813;
	WX2817<=WX2828 and WX3589;
	WX2818<=WX2824 and WX2819;
	WX2821<=CRC_OUT_7_17 and WX3590;
	WX2822<=WX4989 and WX2823;
	WX2825<=WX3099 and WX3590;
	WX2826<=WX3696 and WX2827;
	WX2831<=WX2842 and WX3589;
	WX2832<=WX2838 and WX2833;
	WX2835<=CRC_OUT_7_16 and WX3590;
	WX2836<=WX4996 and WX2837;
	WX2839<=WX3101 and WX3590;
	WX2840<=WX3703 and WX2841;
	WX2845<=WX2856 and WX3589;
	WX2846<=WX2852 and WX2847;
	WX2849<=CRC_OUT_7_15 and WX3590;
	WX2850<=WX5003 and WX2851;
	WX2853<=WX3103 and WX3590;
	WX2854<=WX3710 and WX2855;
	WX2859<=WX2870 and WX3589;
	WX2860<=WX2866 and WX2861;
	WX2863<=CRC_OUT_7_14 and WX3590;
	WX2864<=WX5010 and WX2865;
	WX2867<=WX3105 and WX3590;
	WX2868<=WX3717 and WX2869;
	WX2873<=WX2884 and WX3589;
	WX2874<=WX2880 and WX2875;
	WX2877<=CRC_OUT_7_13 and WX3590;
	WX2878<=WX5017 and WX2879;
	WX2881<=WX3107 and WX3590;
	WX2882<=WX3724 and WX2883;
	WX2887<=WX2898 and WX3589;
	WX2888<=WX2894 and WX2889;
	WX2891<=CRC_OUT_7_12 and WX3590;
	WX2892<=WX5024 and WX2893;
	WX2895<=WX3109 and WX3590;
	WX2896<=WX3731 and WX2897;
	WX2901<=WX2912 and WX3589;
	WX2902<=WX2908 and WX2903;
	WX2905<=CRC_OUT_7_11 and WX3590;
	WX2906<=WX5031 and WX2907;
	WX2909<=WX3111 and WX3590;
	WX2910<=WX3738 and WX2911;
	WX2915<=WX2926 and WX3589;
	WX2916<=WX2922 and WX2917;
	WX2919<=CRC_OUT_7_10 and WX3590;
	WX2920<=WX5038 and WX2921;
	WX2923<=WX3113 and WX3590;
	WX2924<=WX3745 and WX2925;
	WX2929<=WX2940 and WX3589;
	WX2930<=WX2936 and WX2931;
	WX2933<=CRC_OUT_7_9 and WX3590;
	WX2934<=WX5045 and WX2935;
	WX2937<=WX3115 and WX3590;
	WX2938<=WX3752 and WX2939;
	WX2943<=WX2954 and WX3589;
	WX2944<=WX2950 and WX2945;
	WX2947<=CRC_OUT_7_8 and WX3590;
	WX2948<=WX5052 and WX2949;
	WX2951<=WX3117 and WX3590;
	WX2952<=WX3759 and WX2953;
	WX2957<=WX2968 and WX3589;
	WX2958<=WX2964 and WX2959;
	WX2961<=CRC_OUT_7_7 and WX3590;
	WX2962<=WX5059 and WX2963;
	WX2965<=WX3119 and WX3590;
	WX2966<=WX3766 and WX2967;
	WX2971<=WX2982 and WX3589;
	WX2972<=WX2978 and WX2973;
	WX2975<=CRC_OUT_7_6 and WX3590;
	WX2976<=WX5066 and WX2977;
	WX2979<=WX3121 and WX3590;
	WX2980<=WX3773 and WX2981;
	WX2985<=WX2996 and WX3589;
	WX2986<=WX2992 and WX2987;
	WX2989<=CRC_OUT_7_5 and WX3590;
	WX2990<=WX5073 and WX2991;
	WX2993<=WX3123 and WX3590;
	WX2994<=WX3780 and WX2995;
	WX2999<=WX3010 and WX3589;
	WX3000<=WX3006 and WX3001;
	WX3003<=CRC_OUT_7_4 and WX3590;
	WX3004<=WX5080 and WX3005;
	WX3007<=WX3125 and WX3590;
	WX3008<=WX3787 and WX3009;
	WX3013<=WX3024 and WX3589;
	WX3014<=WX3020 and WX3015;
	WX3017<=CRC_OUT_7_3 and WX3590;
	WX3018<=WX5087 and WX3019;
	WX3021<=WX3127 and WX3590;
	WX3022<=WX3794 and WX3023;
	WX3027<=WX3038 and WX3589;
	WX3028<=WX3034 and WX3029;
	WX3031<=CRC_OUT_7_2 and WX3590;
	WX3032<=WX5094 and WX3033;
	WX3035<=WX3129 and WX3590;
	WX3036<=WX3801 and WX3037;
	WX3041<=WX3052 and WX3589;
	WX3042<=WX3048 and WX3043;
	WX3045<=CRC_OUT_7_1 and WX3590;
	WX3046<=WX5101 and WX3047;
	WX3049<=WX3131 and WX3590;
	WX3050<=WX3808 and WX3051;
	WX3055<=WX3066 and WX3589;
	WX3056<=WX3062 and WX3057;
	WX3059<=CRC_OUT_7_0 and WX3590;
	WX3060<=WX5108 and WX3061;
	WX3063<=WX3133 and WX3590;
	WX3064<=WX3815 and WX3065;
	WX3070<=WX3073 and RESET;
	WX3072<=WX3075 and RESET;
	WX3074<=WX3077 and RESET;
	WX3076<=WX3079 and RESET;
	WX3078<=WX3081 and RESET;
	WX3080<=WX3083 and RESET;
	WX3082<=WX3085 and RESET;
	WX3084<=WX3087 and RESET;
	WX3086<=WX3089 and RESET;
	WX3088<=WX3091 and RESET;
	WX3090<=WX3093 and RESET;
	WX3092<=WX3095 and RESET;
	WX3094<=WX3097 and RESET;
	WX3096<=WX3099 and RESET;
	WX3098<=WX3101 and RESET;
	WX3100<=WX3103 and RESET;
	WX3102<=WX3105 and RESET;
	WX3104<=WX3107 and RESET;
	WX3106<=WX3109 and RESET;
	WX3108<=WX3111 and RESET;
	WX3110<=WX3113 and RESET;
	WX3112<=WX3115 and RESET;
	WX3114<=WX3117 and RESET;
	WX3116<=WX3119 and RESET;
	WX3118<=WX3121 and RESET;
	WX3120<=WX3123 and RESET;
	WX3122<=WX3125 and RESET;
	WX3124<=WX3127 and RESET;
	WX3126<=WX3129 and RESET;
	WX3128<=WX3131 and RESET;
	WX3130<=WX3133 and RESET;
	WX3132<=WX3069 and RESET;
	WX3230<=WX2634 and RESET;
	WX3232<=WX2648 and RESET;
	WX3234<=WX2662 and RESET;
	WX3236<=WX2676 and RESET;
	WX3238<=WX2690 and RESET;
	WX3240<=WX2704 and RESET;
	WX3242<=WX2718 and RESET;
	WX3244<=WX2732 and RESET;
	WX3246<=WX2746 and RESET;
	WX3248<=WX2760 and RESET;
	WX3250<=WX2774 and RESET;
	WX3252<=WX2788 and RESET;
	WX3254<=WX2802 and RESET;
	WX3256<=WX2816 and RESET;
	WX3258<=WX2830 and RESET;
	WX3260<=WX2844 and RESET;
	WX3262<=WX2858 and RESET;
	WX3264<=WX2872 and RESET;
	WX3266<=WX2886 and RESET;
	WX3268<=WX2900 and RESET;
	WX3270<=WX2914 and RESET;
	WX3272<=WX2928 and RESET;
	WX3274<=WX2942 and RESET;
	WX3276<=WX2956 and RESET;
	WX3278<=WX2970 and RESET;
	WX3280<=WX2984 and RESET;
	WX3282<=WX2998 and RESET;
	WX3284<=WX3012 and RESET;
	WX3286<=WX3026 and RESET;
	WX3288<=WX3040 and RESET;
	WX3290<=WX3054 and RESET;
	WX3292<=WX3068 and RESET;
	WX3294<=WX3231 and RESET;
	WX3296<=WX3233 and RESET;
	WX3298<=WX3235 and RESET;
	WX3300<=WX3237 and RESET;
	WX3302<=WX3239 and RESET;
	WX3304<=WX3241 and RESET;
	WX3306<=WX3243 and RESET;
	WX3308<=WX3245 and RESET;
	WX3310<=WX3247 and RESET;
	WX3312<=WX3249 and RESET;
	WX3314<=WX3251 and RESET;
	WX3316<=WX3253 and RESET;
	WX3318<=WX3255 and RESET;
	WX3320<=WX3257 and RESET;
	WX3322<=WX3259 and RESET;
	WX3324<=WX3261 and RESET;
	WX3326<=WX3263 and RESET;
	WX3328<=WX3265 and RESET;
	WX3330<=WX3267 and RESET;
	WX3332<=WX3269 and RESET;
	WX3334<=WX3271 and RESET;
	WX3336<=WX3273 and RESET;
	WX3338<=WX3275 and RESET;
	WX3340<=WX3277 and RESET;
	WX3342<=WX3279 and RESET;
	WX3344<=WX3281 and RESET;
	WX3346<=WX3283 and RESET;
	WX3348<=WX3285 and RESET;
	WX3350<=WX3287 and RESET;
	WX3352<=WX3289 and RESET;
	WX3354<=WX3291 and RESET;
	WX3356<=WX3293 and RESET;
	WX3358<=WX3295 and RESET;
	WX3360<=WX3297 and RESET;
	WX3362<=WX3299 and RESET;
	WX3364<=WX3301 and RESET;
	WX3366<=WX3303 and RESET;
	WX3368<=WX3305 and RESET;
	WX3370<=WX3307 and RESET;
	WX3372<=WX3309 and RESET;
	WX3374<=WX3311 and RESET;
	WX3376<=WX3313 and RESET;
	WX3378<=WX3315 and RESET;
	WX3380<=WX3317 and RESET;
	WX3382<=WX3319 and RESET;
	WX3384<=WX3321 and RESET;
	WX3386<=WX3323 and RESET;
	WX3388<=WX3325 and RESET;
	WX3390<=WX3327 and RESET;
	WX3392<=WX3329 and RESET;
	WX3394<=WX3331 and RESET;
	WX3396<=WX3333 and RESET;
	WX3398<=WX3335 and RESET;
	WX3400<=WX3337 and RESET;
	WX3402<=WX3339 and RESET;
	WX3404<=WX3341 and RESET;
	WX3406<=WX3343 and RESET;
	WX3408<=WX3345 and RESET;
	WX3410<=WX3347 and RESET;
	WX3412<=WX3349 and RESET;
	WX3414<=WX3351 and RESET;
	WX3416<=WX3353 and RESET;
	WX3418<=WX3355 and RESET;
	WX3420<=WX3357 and RESET;
	WX3422<=WX3359 and RESET;
	WX3424<=WX3361 and RESET;
	WX3426<=WX3363 and RESET;
	WX3428<=WX3365 and RESET;
	WX3430<=WX3367 and RESET;
	WX3432<=WX3369 and RESET;
	WX3434<=WX3371 and RESET;
	WX3436<=WX3373 and RESET;
	WX3438<=WX3375 and RESET;
	WX3440<=WX3377 and RESET;
	WX3442<=WX3379 and RESET;
	WX3444<=WX3381 and RESET;
	WX3446<=WX3383 and RESET;
	WX3448<=WX3385 and RESET;
	WX3450<=WX3387 and RESET;
	WX3452<=WX3389 and RESET;
	WX3454<=WX3391 and RESET;
	WX3456<=WX3393 and RESET;
	WX3458<=WX3395 and RESET;
	WX3460<=WX3397 and RESET;
	WX3462<=WX3399 and RESET;
	WX3464<=WX3401 and RESET;
	WX3466<=WX3403 and RESET;
	WX3468<=WX3405 and RESET;
	WX3470<=WX3407 and RESET;
	WX3472<=WX3409 and RESET;
	WX3474<=WX3411 and RESET;
	WX3476<=WX3413 and RESET;
	WX3478<=WX3415 and RESET;
	WX3480<=WX3417 and RESET;
	WX3482<=WX3419 and RESET;
	WX3484<=WX3421 and RESET;
	WX3593<=WX3592 and WX3591;
	WX3594<=WX3166 and WX3595;
	WX3600<=WX3599 and WX3591;
	WX3601<=WX3167 and WX3602;
	WX3607<=WX3606 and WX3591;
	WX3608<=WX3168 and WX3609;
	WX3614<=WX3613 and WX3591;
	WX3615<=WX3169 and WX3616;
	WX3621<=WX3620 and WX3591;
	WX3622<=WX3170 and WX3623;
	WX3628<=WX3627 and WX3591;
	WX3629<=WX3171 and WX3630;
	WX3635<=WX3634 and WX3591;
	WX3636<=WX3172 and WX3637;
	WX3642<=WX3641 and WX3591;
	WX3643<=WX3173 and WX3644;
	WX3649<=WX3648 and WX3591;
	WX3650<=WX3174 and WX3651;
	WX3656<=WX3655 and WX3591;
	WX3657<=WX3175 and WX3658;
	WX3663<=WX3662 and WX3591;
	WX3664<=WX3176 and WX3665;
	WX3670<=WX3669 and WX3591;
	WX3671<=WX3177 and WX3672;
	WX3677<=WX3676 and WX3591;
	WX3678<=WX3178 and WX3679;
	WX3684<=WX3683 and WX3591;
	WX3685<=WX3179 and WX3686;
	WX3691<=WX3690 and WX3591;
	WX3692<=WX3180 and WX3693;
	WX3698<=WX3697 and WX3591;
	WX3699<=WX3181 and WX3700;
	WX3705<=WX3704 and WX3591;
	WX3706<=WX3182 and WX3707;
	WX3712<=WX3711 and WX3591;
	WX3713<=WX3183 and WX3714;
	WX3719<=WX3718 and WX3591;
	WX3720<=WX3184 and WX3721;
	WX3726<=WX3725 and WX3591;
	WX3727<=WX3185 and WX3728;
	WX3733<=WX3732 and WX3591;
	WX3734<=WX3186 and WX3735;
	WX3740<=WX3739 and WX3591;
	WX3741<=WX3187 and WX3742;
	WX3747<=WX3746 and WX3591;
	WX3748<=WX3188 and WX3749;
	WX3754<=WX3753 and WX3591;
	WX3755<=WX3189 and WX3756;
	WX3761<=WX3760 and WX3591;
	WX3762<=WX3190 and WX3763;
	WX3768<=WX3767 and WX3591;
	WX3769<=WX3191 and WX3770;
	WX3775<=WX3774 and WX3591;
	WX3776<=WX3192 and WX3777;
	WX3782<=WX3781 and WX3591;
	WX3783<=WX3193 and WX3784;
	WX3789<=WX3788 and WX3591;
	WX3790<=WX3194 and WX3791;
	WX3796<=WX3795 and WX3591;
	WX3797<=WX3195 and WX3798;
	WX3803<=WX3802 and WX3591;
	WX3804<=WX3196 and WX3805;
	WX3810<=WX3809 and WX3591;
	WX3811<=WX3197 and WX3812;
	WX3850<=WX3820 and WX3849;
	WX3852<=WX3848 and WX3849;
	WX3854<=WX3847 and WX3849;
	WX3856<=WX3846 and WX3849;
	WX3858<=WX3819 and WX3849;
	WX3860<=WX3845 and WX3849;
	WX3862<=WX3844 and WX3849;
	WX3864<=WX3843 and WX3849;
	WX3866<=WX3842 and WX3849;
	WX3868<=WX3841 and WX3849;
	WX3870<=WX3840 and WX3849;
	WX3872<=WX3818 and WX3849;
	WX3874<=WX3839 and WX3849;
	WX3876<=WX3838 and WX3849;
	WX3878<=WX3837 and WX3849;
	WX3880<=WX3836 and WX3849;
	WX3882<=WX3817 and WX3849;
	WX3884<=WX3835 and WX3849;
	WX3886<=WX3834 and WX3849;
	WX3888<=WX3833 and WX3849;
	WX3890<=WX3832 and WX3849;
	WX3892<=WX3831 and WX3849;
	WX3894<=WX3830 and WX3849;
	WX3896<=WX3829 and WX3849;
	WX3898<=WX3828 and WX3849;
	WX3900<=WX3827 and WX3849;
	WX3902<=WX3826 and WX3849;
	WX3904<=WX3825 and WX3849;
	WX3906<=WX3824 and WX3849;
	WX3908<=WX3823 and WX3849;
	WX3910<=WX3822 and WX3849;
	WX3912<=WX3821 and WX3849;
	WX3914<=WX3925 and WX4882;
	WX3915<=WX3921 and WX3916;
	WX3918<=CRC_OUT_6_31 and WX4883;
	WX3919<=WX6184 and WX3920;
	WX3922<=WX4364 and WX4883;
	WX3923<=WX4891 and WX3924;
	WX3928<=WX3939 and WX4882;
	WX3929<=WX3935 and WX3930;
	WX3932<=CRC_OUT_6_30 and WX4883;
	WX3933<=WX6191 and WX3934;
	WX3936<=WX4366 and WX4883;
	WX3937<=WX4898 and WX3938;
	WX3942<=WX3953 and WX4882;
	WX3943<=WX3949 and WX3944;
	WX3946<=CRC_OUT_6_29 and WX4883;
	WX3947<=WX6198 and WX3948;
	WX3950<=WX4368 and WX4883;
	WX3951<=WX4905 and WX3952;
	WX3956<=WX3967 and WX4882;
	WX3957<=WX3963 and WX3958;
	WX3960<=CRC_OUT_6_28 and WX4883;
	WX3961<=WX6205 and WX3962;
	WX3964<=WX4370 and WX4883;
	WX3965<=WX4912 and WX3966;
	WX3970<=WX3981 and WX4882;
	WX3971<=WX3977 and WX3972;
	WX3974<=CRC_OUT_6_27 and WX4883;
	WX3975<=WX6212 and WX3976;
	WX3978<=WX4372 and WX4883;
	WX3979<=WX4919 and WX3980;
	WX3984<=WX3995 and WX4882;
	WX3985<=WX3991 and WX3986;
	WX3988<=CRC_OUT_6_26 and WX4883;
	WX3989<=WX6219 and WX3990;
	WX3992<=WX4374 and WX4883;
	WX3993<=WX4926 and WX3994;
	WX3998<=WX4009 and WX4882;
	WX3999<=WX4005 and WX4000;
	WX4002<=CRC_OUT_6_25 and WX4883;
	WX4003<=WX6226 and WX4004;
	WX4006<=WX4376 and WX4883;
	WX4007<=WX4933 and WX4008;
	WX4012<=WX4023 and WX4882;
	WX4013<=WX4019 and WX4014;
	WX4016<=CRC_OUT_6_24 and WX4883;
	WX4017<=WX6233 and WX4018;
	WX4020<=WX4378 and WX4883;
	WX4021<=WX4940 and WX4022;
	WX4026<=WX4037 and WX4882;
	WX4027<=WX4033 and WX4028;
	WX4030<=CRC_OUT_6_23 and WX4883;
	WX4031<=WX6240 and WX4032;
	WX4034<=WX4380 and WX4883;
	WX4035<=WX4947 and WX4036;
	WX4040<=WX4051 and WX4882;
	WX4041<=WX4047 and WX4042;
	WX4044<=CRC_OUT_6_22 and WX4883;
	WX4045<=WX6247 and WX4046;
	WX4048<=WX4382 and WX4883;
	WX4049<=WX4954 and WX4050;
	WX4054<=WX4065 and WX4882;
	WX4055<=WX4061 and WX4056;
	WX4058<=CRC_OUT_6_21 and WX4883;
	WX4059<=WX6254 and WX4060;
	WX4062<=WX4384 and WX4883;
	WX4063<=WX4961 and WX4064;
	WX4068<=WX4079 and WX4882;
	WX4069<=WX4075 and WX4070;
	WX4072<=CRC_OUT_6_20 and WX4883;
	WX4073<=WX6261 and WX4074;
	WX4076<=WX4386 and WX4883;
	WX4077<=WX4968 and WX4078;
	WX4082<=WX4093 and WX4882;
	WX4083<=WX4089 and WX4084;
	WX4086<=CRC_OUT_6_19 and WX4883;
	WX4087<=WX6268 and WX4088;
	WX4090<=WX4388 and WX4883;
	WX4091<=WX4975 and WX4092;
	WX4096<=WX4107 and WX4882;
	WX4097<=WX4103 and WX4098;
	WX4100<=CRC_OUT_6_18 and WX4883;
	WX4101<=WX6275 and WX4102;
	WX4104<=WX4390 and WX4883;
	WX4105<=WX4982 and WX4106;
	WX4110<=WX4121 and WX4882;
	WX4111<=WX4117 and WX4112;
	WX4114<=CRC_OUT_6_17 and WX4883;
	WX4115<=WX6282 and WX4116;
	WX4118<=WX4392 and WX4883;
	WX4119<=WX4989 and WX4120;
	WX4124<=WX4135 and WX4882;
	WX4125<=WX4131 and WX4126;
	WX4128<=CRC_OUT_6_16 and WX4883;
	WX4129<=WX6289 and WX4130;
	WX4132<=WX4394 and WX4883;
	WX4133<=WX4996 and WX4134;
	WX4138<=WX4149 and WX4882;
	WX4139<=WX4145 and WX4140;
	WX4142<=CRC_OUT_6_15 and WX4883;
	WX4143<=WX6296 and WX4144;
	WX4146<=WX4396 and WX4883;
	WX4147<=WX5003 and WX4148;
	WX4152<=WX4163 and WX4882;
	WX4153<=WX4159 and WX4154;
	WX4156<=CRC_OUT_6_14 and WX4883;
	WX4157<=WX6303 and WX4158;
	WX4160<=WX4398 and WX4883;
	WX4161<=WX5010 and WX4162;
	WX4166<=WX4177 and WX4882;
	WX4167<=WX4173 and WX4168;
	WX4170<=CRC_OUT_6_13 and WX4883;
	WX4171<=WX6310 and WX4172;
	WX4174<=WX4400 and WX4883;
	WX4175<=WX5017 and WX4176;
	WX4180<=WX4191 and WX4882;
	WX4181<=WX4187 and WX4182;
	WX4184<=CRC_OUT_6_12 and WX4883;
	WX4185<=WX6317 and WX4186;
	WX4188<=WX4402 and WX4883;
	WX4189<=WX5024 and WX4190;
	WX4194<=WX4205 and WX4882;
	WX4195<=WX4201 and WX4196;
	WX4198<=CRC_OUT_6_11 and WX4883;
	WX4199<=WX6324 and WX4200;
	WX4202<=WX4404 and WX4883;
	WX4203<=WX5031 and WX4204;
	WX4208<=WX4219 and WX4882;
	WX4209<=WX4215 and WX4210;
	WX4212<=CRC_OUT_6_10 and WX4883;
	WX4213<=WX6331 and WX4214;
	WX4216<=WX4406 and WX4883;
	WX4217<=WX5038 and WX4218;
	WX4222<=WX4233 and WX4882;
	WX4223<=WX4229 and WX4224;
	WX4226<=CRC_OUT_6_9 and WX4883;
	WX4227<=WX6338 and WX4228;
	WX4230<=WX4408 and WX4883;
	WX4231<=WX5045 and WX4232;
	WX4236<=WX4247 and WX4882;
	WX4237<=WX4243 and WX4238;
	WX4240<=CRC_OUT_6_8 and WX4883;
	WX4241<=WX6345 and WX4242;
	WX4244<=WX4410 and WX4883;
	WX4245<=WX5052 and WX4246;
	WX4250<=WX4261 and WX4882;
	WX4251<=WX4257 and WX4252;
	WX4254<=CRC_OUT_6_7 and WX4883;
	WX4255<=WX6352 and WX4256;
	WX4258<=WX4412 and WX4883;
	WX4259<=WX5059 and WX4260;
	WX4264<=WX4275 and WX4882;
	WX4265<=WX4271 and WX4266;
	WX4268<=CRC_OUT_6_6 and WX4883;
	WX4269<=WX6359 and WX4270;
	WX4272<=WX4414 and WX4883;
	WX4273<=WX5066 and WX4274;
	WX4278<=WX4289 and WX4882;
	WX4279<=WX4285 and WX4280;
	WX4282<=CRC_OUT_6_5 and WX4883;
	WX4283<=WX6366 and WX4284;
	WX4286<=WX4416 and WX4883;
	WX4287<=WX5073 and WX4288;
	WX4292<=WX4303 and WX4882;
	WX4293<=WX4299 and WX4294;
	WX4296<=CRC_OUT_6_4 and WX4883;
	WX4297<=WX6373 and WX4298;
	WX4300<=WX4418 and WX4883;
	WX4301<=WX5080 and WX4302;
	WX4306<=WX4317 and WX4882;
	WX4307<=WX4313 and WX4308;
	WX4310<=CRC_OUT_6_3 and WX4883;
	WX4311<=WX6380 and WX4312;
	WX4314<=WX4420 and WX4883;
	WX4315<=WX5087 and WX4316;
	WX4320<=WX4331 and WX4882;
	WX4321<=WX4327 and WX4322;
	WX4324<=CRC_OUT_6_2 and WX4883;
	WX4325<=WX6387 and WX4326;
	WX4328<=WX4422 and WX4883;
	WX4329<=WX5094 and WX4330;
	WX4334<=WX4345 and WX4882;
	WX4335<=WX4341 and WX4336;
	WX4338<=CRC_OUT_6_1 and WX4883;
	WX4339<=WX6394 and WX4340;
	WX4342<=WX4424 and WX4883;
	WX4343<=WX5101 and WX4344;
	WX4348<=WX4359 and WX4882;
	WX4349<=WX4355 and WX4350;
	WX4352<=CRC_OUT_6_0 and WX4883;
	WX4353<=WX6401 and WX4354;
	WX4356<=WX4426 and WX4883;
	WX4357<=WX5108 and WX4358;
	WX4363<=WX4366 and RESET;
	WX4365<=WX4368 and RESET;
	WX4367<=WX4370 and RESET;
	WX4369<=WX4372 and RESET;
	WX4371<=WX4374 and RESET;
	WX4373<=WX4376 and RESET;
	WX4375<=WX4378 and RESET;
	WX4377<=WX4380 and RESET;
	WX4379<=WX4382 and RESET;
	WX4381<=WX4384 and RESET;
	WX4383<=WX4386 and RESET;
	WX4385<=WX4388 and RESET;
	WX4387<=WX4390 and RESET;
	WX4389<=WX4392 and RESET;
	WX4391<=WX4394 and RESET;
	WX4393<=WX4396 and RESET;
	WX4395<=WX4398 and RESET;
	WX4397<=WX4400 and RESET;
	WX4399<=WX4402 and RESET;
	WX4401<=WX4404 and RESET;
	WX4403<=WX4406 and RESET;
	WX4405<=WX4408 and RESET;
	WX4407<=WX4410 and RESET;
	WX4409<=WX4412 and RESET;
	WX4411<=WX4414 and RESET;
	WX4413<=WX4416 and RESET;
	WX4415<=WX4418 and RESET;
	WX4417<=WX4420 and RESET;
	WX4419<=WX4422 and RESET;
	WX4421<=WX4424 and RESET;
	WX4423<=WX4426 and RESET;
	WX4425<=WX4362 and RESET;
	WX4523<=WX3927 and RESET;
	WX4525<=WX3941 and RESET;
	WX4527<=WX3955 and RESET;
	WX4529<=WX3969 and RESET;
	WX4531<=WX3983 and RESET;
	WX4533<=WX3997 and RESET;
	WX4535<=WX4011 and RESET;
	WX4537<=WX4025 and RESET;
	WX4539<=WX4039 and RESET;
	WX4541<=WX4053 and RESET;
	WX4543<=WX4067 and RESET;
	WX4545<=WX4081 and RESET;
	WX4547<=WX4095 and RESET;
	WX4549<=WX4109 and RESET;
	WX4551<=WX4123 and RESET;
	WX4553<=WX4137 and RESET;
	WX4555<=WX4151 and RESET;
	WX4557<=WX4165 and RESET;
	WX4559<=WX4179 and RESET;
	WX4561<=WX4193 and RESET;
	WX4563<=WX4207 and RESET;
	WX4565<=WX4221 and RESET;
	WX4567<=WX4235 and RESET;
	WX4569<=WX4249 and RESET;
	WX4571<=WX4263 and RESET;
	WX4573<=WX4277 and RESET;
	WX4575<=WX4291 and RESET;
	WX4577<=WX4305 and RESET;
	WX4579<=WX4319 and RESET;
	WX4581<=WX4333 and RESET;
	WX4583<=WX4347 and RESET;
	WX4585<=WX4361 and RESET;
	WX4587<=WX4524 and RESET;
	WX4589<=WX4526 and RESET;
	WX4591<=WX4528 and RESET;
	WX4593<=WX4530 and RESET;
	WX4595<=WX4532 and RESET;
	WX4597<=WX4534 and RESET;
	WX4599<=WX4536 and RESET;
	WX4601<=WX4538 and RESET;
	WX4603<=WX4540 and RESET;
	WX4605<=WX4542 and RESET;
	WX4607<=WX4544 and RESET;
	WX4609<=WX4546 and RESET;
	WX4611<=WX4548 and RESET;
	WX4613<=WX4550 and RESET;
	WX4615<=WX4552 and RESET;
	WX4617<=WX4554 and RESET;
	WX4619<=WX4556 and RESET;
	WX4621<=WX4558 and RESET;
	WX4623<=WX4560 and RESET;
	WX4625<=WX4562 and RESET;
	WX4627<=WX4564 and RESET;
	WX4629<=WX4566 and RESET;
	WX4631<=WX4568 and RESET;
	WX4633<=WX4570 and RESET;
	WX4635<=WX4572 and RESET;
	WX4637<=WX4574 and RESET;
	WX4639<=WX4576 and RESET;
	WX4641<=WX4578 and RESET;
	WX4643<=WX4580 and RESET;
	WX4645<=WX4582 and RESET;
	WX4647<=WX4584 and RESET;
	WX4649<=WX4586 and RESET;
	WX4651<=WX4588 and RESET;
	WX4653<=WX4590 and RESET;
	WX4655<=WX4592 and RESET;
	WX4657<=WX4594 and RESET;
	WX4659<=WX4596 and RESET;
	WX4661<=WX4598 and RESET;
	WX4663<=WX4600 and RESET;
	WX4665<=WX4602 and RESET;
	WX4667<=WX4604 and RESET;
	WX4669<=WX4606 and RESET;
	WX4671<=WX4608 and RESET;
	WX4673<=WX4610 and RESET;
	WX4675<=WX4612 and RESET;
	WX4677<=WX4614 and RESET;
	WX4679<=WX4616 and RESET;
	WX4681<=WX4618 and RESET;
	WX4683<=WX4620 and RESET;
	WX4685<=WX4622 and RESET;
	WX4687<=WX4624 and RESET;
	WX4689<=WX4626 and RESET;
	WX4691<=WX4628 and RESET;
	WX4693<=WX4630 and RESET;
	WX4695<=WX4632 and RESET;
	WX4697<=WX4634 and RESET;
	WX4699<=WX4636 and RESET;
	WX4701<=WX4638 and RESET;
	WX4703<=WX4640 and RESET;
	WX4705<=WX4642 and RESET;
	WX4707<=WX4644 and RESET;
	WX4709<=WX4646 and RESET;
	WX4711<=WX4648 and RESET;
	WX4713<=WX4650 and RESET;
	WX4715<=WX4652 and RESET;
	WX4717<=WX4654 and RESET;
	WX4719<=WX4656 and RESET;
	WX4721<=WX4658 and RESET;
	WX4723<=WX4660 and RESET;
	WX4725<=WX4662 and RESET;
	WX4727<=WX4664 and RESET;
	WX4729<=WX4666 and RESET;
	WX4731<=WX4668 and RESET;
	WX4733<=WX4670 and RESET;
	WX4735<=WX4672 and RESET;
	WX4737<=WX4674 and RESET;
	WX4739<=WX4676 and RESET;
	WX4741<=WX4678 and RESET;
	WX4743<=WX4680 and RESET;
	WX4745<=WX4682 and RESET;
	WX4747<=WX4684 and RESET;
	WX4749<=WX4686 and RESET;
	WX4751<=WX4688 and RESET;
	WX4753<=WX4690 and RESET;
	WX4755<=WX4692 and RESET;
	WX4757<=WX4694 and RESET;
	WX4759<=WX4696 and RESET;
	WX4761<=WX4698 and RESET;
	WX4763<=WX4700 and RESET;
	WX4765<=WX4702 and RESET;
	WX4767<=WX4704 and RESET;
	WX4769<=WX4706 and RESET;
	WX4771<=WX4708 and RESET;
	WX4773<=WX4710 and RESET;
	WX4775<=WX4712 and RESET;
	WX4777<=WX4714 and RESET;
	WX4886<=WX4885 and WX4884;
	WX4887<=WX4459 and WX4888;
	WX4893<=WX4892 and WX4884;
	WX4894<=WX4460 and WX4895;
	WX4900<=WX4899 and WX4884;
	WX4901<=WX4461 and WX4902;
	WX4907<=WX4906 and WX4884;
	WX4908<=WX4462 and WX4909;
	WX4914<=WX4913 and WX4884;
	WX4915<=WX4463 and WX4916;
	WX4921<=WX4920 and WX4884;
	WX4922<=WX4464 and WX4923;
	WX4928<=WX4927 and WX4884;
	WX4929<=WX4465 and WX4930;
	WX4935<=WX4934 and WX4884;
	WX4936<=WX4466 and WX4937;
	WX4942<=WX4941 and WX4884;
	WX4943<=WX4467 and WX4944;
	WX4949<=WX4948 and WX4884;
	WX4950<=WX4468 and WX4951;
	WX4956<=WX4955 and WX4884;
	WX4957<=WX4469 and WX4958;
	WX4963<=WX4962 and WX4884;
	WX4964<=WX4470 and WX4965;
	WX4970<=WX4969 and WX4884;
	WX4971<=WX4471 and WX4972;
	WX4977<=WX4976 and WX4884;
	WX4978<=WX4472 and WX4979;
	WX4984<=WX4983 and WX4884;
	WX4985<=WX4473 and WX4986;
	WX4991<=WX4990 and WX4884;
	WX4992<=WX4474 and WX4993;
	WX4998<=WX4997 and WX4884;
	WX4999<=WX4475 and WX5000;
	WX5005<=WX5004 and WX4884;
	WX5006<=WX4476 and WX5007;
	WX5012<=WX5011 and WX4884;
	WX5013<=WX4477 and WX5014;
	WX5019<=WX5018 and WX4884;
	WX5020<=WX4478 and WX5021;
	WX5026<=WX5025 and WX4884;
	WX5027<=WX4479 and WX5028;
	WX5033<=WX5032 and WX4884;
	WX5034<=WX4480 and WX5035;
	WX5040<=WX5039 and WX4884;
	WX5041<=WX4481 and WX5042;
	WX5047<=WX5046 and WX4884;
	WX5048<=WX4482 and WX5049;
	WX5054<=WX5053 and WX4884;
	WX5055<=WX4483 and WX5056;
	WX5061<=WX5060 and WX4884;
	WX5062<=WX4484 and WX5063;
	WX5068<=WX5067 and WX4884;
	WX5069<=WX4485 and WX5070;
	WX5075<=WX5074 and WX4884;
	WX5076<=WX4486 and WX5077;
	WX5082<=WX5081 and WX4884;
	WX5083<=WX4487 and WX5084;
	WX5089<=WX5088 and WX4884;
	WX5090<=WX4488 and WX5091;
	WX5096<=WX5095 and WX4884;
	WX5097<=WX4489 and WX5098;
	WX5103<=WX5102 and WX4884;
	WX5104<=WX4490 and WX5105;
	WX5143<=WX5113 and WX5142;
	WX5145<=WX5141 and WX5142;
	WX5147<=WX5140 and WX5142;
	WX5149<=WX5139 and WX5142;
	WX5151<=WX5112 and WX5142;
	WX5153<=WX5138 and WX5142;
	WX5155<=WX5137 and WX5142;
	WX5157<=WX5136 and WX5142;
	WX5159<=WX5135 and WX5142;
	WX5161<=WX5134 and WX5142;
	WX5163<=WX5133 and WX5142;
	WX5165<=WX5111 and WX5142;
	WX5167<=WX5132 and WX5142;
	WX5169<=WX5131 and WX5142;
	WX5171<=WX5130 and WX5142;
	WX5173<=WX5129 and WX5142;
	WX5175<=WX5110 and WX5142;
	WX5177<=WX5128 and WX5142;
	WX5179<=WX5127 and WX5142;
	WX5181<=WX5126 and WX5142;
	WX5183<=WX5125 and WX5142;
	WX5185<=WX5124 and WX5142;
	WX5187<=WX5123 and WX5142;
	WX5189<=WX5122 and WX5142;
	WX5191<=WX5121 and WX5142;
	WX5193<=WX5120 and WX5142;
	WX5195<=WX5119 and WX5142;
	WX5197<=WX5118 and WX5142;
	WX5199<=WX5117 and WX5142;
	WX5201<=WX5116 and WX5142;
	WX5203<=WX5115 and WX5142;
	WX5205<=WX5114 and WX5142;
	WX5207<=WX5218 and WX6175;
	WX5208<=WX5214 and WX5209;
	WX5211<=CRC_OUT_5_31 and WX6176;
	WX5212<=WX7477 and WX5213;
	WX5215<=WX5657 and WX6176;
	WX5216<=WX6184 and WX5217;
	WX5221<=WX5232 and WX6175;
	WX5222<=WX5228 and WX5223;
	WX5225<=CRC_OUT_5_30 and WX6176;
	WX5226<=WX7484 and WX5227;
	WX5229<=WX5659 and WX6176;
	WX5230<=WX6191 and WX5231;
	WX5235<=WX5246 and WX6175;
	WX5236<=WX5242 and WX5237;
	WX5239<=CRC_OUT_5_29 and WX6176;
	WX5240<=WX7491 and WX5241;
	WX5243<=WX5661 and WX6176;
	WX5244<=WX6198 and WX5245;
	WX5249<=WX5260 and WX6175;
	WX5250<=WX5256 and WX5251;
	WX5253<=CRC_OUT_5_28 and WX6176;
	WX5254<=WX7498 and WX5255;
	WX5257<=WX5663 and WX6176;
	WX5258<=WX6205 and WX5259;
	WX5263<=WX5274 and WX6175;
	WX5264<=WX5270 and WX5265;
	WX5267<=CRC_OUT_5_27 and WX6176;
	WX5268<=WX7505 and WX5269;
	WX5271<=WX5665 and WX6176;
	WX5272<=WX6212 and WX5273;
	WX5277<=WX5288 and WX6175;
	WX5278<=WX5284 and WX5279;
	WX5281<=CRC_OUT_5_26 and WX6176;
	WX5282<=WX7512 and WX5283;
	WX5285<=WX5667 and WX6176;
	WX5286<=WX6219 and WX5287;
	WX5291<=WX5302 and WX6175;
	WX5292<=WX5298 and WX5293;
	WX5295<=CRC_OUT_5_25 and WX6176;
	WX5296<=WX7519 and WX5297;
	WX5299<=WX5669 and WX6176;
	WX5300<=WX6226 and WX5301;
	WX5305<=WX5316 and WX6175;
	WX5306<=WX5312 and WX5307;
	WX5309<=CRC_OUT_5_24 and WX6176;
	WX5310<=WX7526 and WX5311;
	WX5313<=WX5671 and WX6176;
	WX5314<=WX6233 and WX5315;
	WX5319<=WX5330 and WX6175;
	WX5320<=WX5326 and WX5321;
	WX5323<=CRC_OUT_5_23 and WX6176;
	WX5324<=WX7533 and WX5325;
	WX5327<=WX5673 and WX6176;
	WX5328<=WX6240 and WX5329;
	WX5333<=WX5344 and WX6175;
	WX5334<=WX5340 and WX5335;
	WX5337<=CRC_OUT_5_22 and WX6176;
	WX5338<=WX7540 and WX5339;
	WX5341<=WX5675 and WX6176;
	WX5342<=WX6247 and WX5343;
	WX5347<=WX5358 and WX6175;
	WX5348<=WX5354 and WX5349;
	WX5351<=CRC_OUT_5_21 and WX6176;
	WX5352<=WX7547 and WX5353;
	WX5355<=WX5677 and WX6176;
	WX5356<=WX6254 and WX5357;
	WX5361<=WX5372 and WX6175;
	WX5362<=WX5368 and WX5363;
	WX5365<=CRC_OUT_5_20 and WX6176;
	WX5366<=WX7554 and WX5367;
	WX5369<=WX5679 and WX6176;
	WX5370<=WX6261 and WX5371;
	WX5375<=WX5386 and WX6175;
	WX5376<=WX5382 and WX5377;
	WX5379<=CRC_OUT_5_19 and WX6176;
	WX5380<=WX7561 and WX5381;
	WX5383<=WX5681 and WX6176;
	WX5384<=WX6268 and WX5385;
	WX5389<=WX5400 and WX6175;
	WX5390<=WX5396 and WX5391;
	WX5393<=CRC_OUT_5_18 and WX6176;
	WX5394<=WX7568 and WX5395;
	WX5397<=WX5683 and WX6176;
	WX5398<=WX6275 and WX5399;
	WX5403<=WX5414 and WX6175;
	WX5404<=WX5410 and WX5405;
	WX5407<=CRC_OUT_5_17 and WX6176;
	WX5408<=WX7575 and WX5409;
	WX5411<=WX5685 and WX6176;
	WX5412<=WX6282 and WX5413;
	WX5417<=WX5428 and WX6175;
	WX5418<=WX5424 and WX5419;
	WX5421<=CRC_OUT_5_16 and WX6176;
	WX5422<=WX7582 and WX5423;
	WX5425<=WX5687 and WX6176;
	WX5426<=WX6289 and WX5427;
	WX5431<=WX5442 and WX6175;
	WX5432<=WX5438 and WX5433;
	WX5435<=CRC_OUT_5_15 and WX6176;
	WX5436<=WX7589 and WX5437;
	WX5439<=WX5689 and WX6176;
	WX5440<=WX6296 and WX5441;
	WX5445<=WX5456 and WX6175;
	WX5446<=WX5452 and WX5447;
	WX5449<=CRC_OUT_5_14 and WX6176;
	WX5450<=WX7596 and WX5451;
	WX5453<=WX5691 and WX6176;
	WX5454<=WX6303 and WX5455;
	WX5459<=WX5470 and WX6175;
	WX5460<=WX5466 and WX5461;
	WX5463<=CRC_OUT_5_13 and WX6176;
	WX5464<=WX7603 and WX5465;
	WX5467<=WX5693 and WX6176;
	WX5468<=WX6310 and WX5469;
	WX5473<=WX5484 and WX6175;
	WX5474<=WX5480 and WX5475;
	WX5477<=CRC_OUT_5_12 and WX6176;
	WX5478<=WX7610 and WX5479;
	WX5481<=WX5695 and WX6176;
	WX5482<=WX6317 and WX5483;
	WX5487<=WX5498 and WX6175;
	WX5488<=WX5494 and WX5489;
	WX5491<=CRC_OUT_5_11 and WX6176;
	WX5492<=WX7617 and WX5493;
	WX5495<=WX5697 and WX6176;
	WX5496<=WX6324 and WX5497;
	WX5501<=WX5512 and WX6175;
	WX5502<=WX5508 and WX5503;
	WX5505<=CRC_OUT_5_10 and WX6176;
	WX5506<=WX7624 and WX5507;
	WX5509<=WX5699 and WX6176;
	WX5510<=WX6331 and WX5511;
	WX5515<=WX5526 and WX6175;
	WX5516<=WX5522 and WX5517;
	WX5519<=CRC_OUT_5_9 and WX6176;
	WX5520<=WX7631 and WX5521;
	WX5523<=WX5701 and WX6176;
	WX5524<=WX6338 and WX5525;
	WX5529<=WX5540 and WX6175;
	WX5530<=WX5536 and WX5531;
	WX5533<=CRC_OUT_5_8 and WX6176;
	WX5534<=WX7638 and WX5535;
	WX5537<=WX5703 and WX6176;
	WX5538<=WX6345 and WX5539;
	WX5543<=WX5554 and WX6175;
	WX5544<=WX5550 and WX5545;
	WX5547<=CRC_OUT_5_7 and WX6176;
	WX5548<=WX7645 and WX5549;
	WX5551<=WX5705 and WX6176;
	WX5552<=WX6352 and WX5553;
	WX5557<=WX5568 and WX6175;
	WX5558<=WX5564 and WX5559;
	WX5561<=CRC_OUT_5_6 and WX6176;
	WX5562<=WX7652 and WX5563;
	WX5565<=WX5707 and WX6176;
	WX5566<=WX6359 and WX5567;
	WX5571<=WX5582 and WX6175;
	WX5572<=WX5578 and WX5573;
	WX5575<=CRC_OUT_5_5 and WX6176;
	WX5576<=WX7659 and WX5577;
	WX5579<=WX5709 and WX6176;
	WX5580<=WX6366 and WX5581;
	WX5585<=WX5596 and WX6175;
	WX5586<=WX5592 and WX5587;
	WX5589<=CRC_OUT_5_4 and WX6176;
	WX5590<=WX7666 and WX5591;
	WX5593<=WX5711 and WX6176;
	WX5594<=WX6373 and WX5595;
	WX5599<=WX5610 and WX6175;
	WX5600<=WX5606 and WX5601;
	WX5603<=CRC_OUT_5_3 and WX6176;
	WX5604<=WX7673 and WX5605;
	WX5607<=WX5713 and WX6176;
	WX5608<=WX6380 and WX5609;
	WX5613<=WX5624 and WX6175;
	WX5614<=WX5620 and WX5615;
	WX5617<=CRC_OUT_5_2 and WX6176;
	WX5618<=WX7680 and WX5619;
	WX5621<=WX5715 and WX6176;
	WX5622<=WX6387 and WX5623;
	WX5627<=WX5638 and WX6175;
	WX5628<=WX5634 and WX5629;
	WX5631<=CRC_OUT_5_1 and WX6176;
	WX5632<=WX7687 and WX5633;
	WX5635<=WX5717 and WX6176;
	WX5636<=WX6394 and WX5637;
	WX5641<=WX5652 and WX6175;
	WX5642<=WX5648 and WX5643;
	WX5645<=CRC_OUT_5_0 and WX6176;
	WX5646<=WX7694 and WX5647;
	WX5649<=WX5719 and WX6176;
	WX5650<=WX6401 and WX5651;
	WX5656<=WX5659 and RESET;
	WX5658<=WX5661 and RESET;
	WX5660<=WX5663 and RESET;
	WX5662<=WX5665 and RESET;
	WX5664<=WX5667 and RESET;
	WX5666<=WX5669 and RESET;
	WX5668<=WX5671 and RESET;
	WX5670<=WX5673 and RESET;
	WX5672<=WX5675 and RESET;
	WX5674<=WX5677 and RESET;
	WX5676<=WX5679 and RESET;
	WX5678<=WX5681 and RESET;
	WX5680<=WX5683 and RESET;
	WX5682<=WX5685 and RESET;
	WX5684<=WX5687 and RESET;
	WX5686<=WX5689 and RESET;
	WX5688<=WX5691 and RESET;
	WX5690<=WX5693 and RESET;
	WX5692<=WX5695 and RESET;
	WX5694<=WX5697 and RESET;
	WX5696<=WX5699 and RESET;
	WX5698<=WX5701 and RESET;
	WX5700<=WX5703 and RESET;
	WX5702<=WX5705 and RESET;
	WX5704<=WX5707 and RESET;
	WX5706<=WX5709 and RESET;
	WX5708<=WX5711 and RESET;
	WX5710<=WX5713 and RESET;
	WX5712<=WX5715 and RESET;
	WX5714<=WX5717 and RESET;
	WX5716<=WX5719 and RESET;
	WX5718<=WX5655 and RESET;
	WX5816<=WX5220 and RESET;
	WX5818<=WX5234 and RESET;
	WX5820<=WX5248 and RESET;
	WX5822<=WX5262 and RESET;
	WX5824<=WX5276 and RESET;
	WX5826<=WX5290 and RESET;
	WX5828<=WX5304 and RESET;
	WX5830<=WX5318 and RESET;
	WX5832<=WX5332 and RESET;
	WX5834<=WX5346 and RESET;
	WX5836<=WX5360 and RESET;
	WX5838<=WX5374 and RESET;
	WX5840<=WX5388 and RESET;
	WX5842<=WX5402 and RESET;
	WX5844<=WX5416 and RESET;
	WX5846<=WX5430 and RESET;
	WX5848<=WX5444 and RESET;
	WX5850<=WX5458 and RESET;
	WX5852<=WX5472 and RESET;
	WX5854<=WX5486 and RESET;
	WX5856<=WX5500 and RESET;
	WX5858<=WX5514 and RESET;
	WX5860<=WX5528 and RESET;
	WX5862<=WX5542 and RESET;
	WX5864<=WX5556 and RESET;
	WX5866<=WX5570 and RESET;
	WX5868<=WX5584 and RESET;
	WX5870<=WX5598 and RESET;
	WX5872<=WX5612 and RESET;
	WX5874<=WX5626 and RESET;
	WX5876<=WX5640 and RESET;
	WX5878<=WX5654 and RESET;
	WX5880<=WX5817 and RESET;
	WX5882<=WX5819 and RESET;
	WX5884<=WX5821 and RESET;
	WX5886<=WX5823 and RESET;
	WX5888<=WX5825 and RESET;
	WX5890<=WX5827 and RESET;
	WX5892<=WX5829 and RESET;
	WX5894<=WX5831 and RESET;
	WX5896<=WX5833 and RESET;
	WX5898<=WX5835 and RESET;
	WX5900<=WX5837 and RESET;
	WX5902<=WX5839 and RESET;
	WX5904<=WX5841 and RESET;
	WX5906<=WX5843 and RESET;
	WX5908<=WX5845 and RESET;
	WX5910<=WX5847 and RESET;
	WX5912<=WX5849 and RESET;
	WX5914<=WX5851 and RESET;
	WX5916<=WX5853 and RESET;
	WX5918<=WX5855 and RESET;
	WX5920<=WX5857 and RESET;
	WX5922<=WX5859 and RESET;
	WX5924<=WX5861 and RESET;
	WX5926<=WX5863 and RESET;
	WX5928<=WX5865 and RESET;
	WX5930<=WX5867 and RESET;
	WX5932<=WX5869 and RESET;
	WX5934<=WX5871 and RESET;
	WX5936<=WX5873 and RESET;
	WX5938<=WX5875 and RESET;
	WX5940<=WX5877 and RESET;
	WX5942<=WX5879 and RESET;
	WX5944<=WX5881 and RESET;
	WX5946<=WX5883 and RESET;
	WX5948<=WX5885 and RESET;
	WX5950<=WX5887 and RESET;
	WX5952<=WX5889 and RESET;
	WX5954<=WX5891 and RESET;
	WX5956<=WX5893 and RESET;
	WX5958<=WX5895 and RESET;
	WX5960<=WX5897 and RESET;
	WX5962<=WX5899 and RESET;
	WX5964<=WX5901 and RESET;
	WX5966<=WX5903 and RESET;
	WX5968<=WX5905 and RESET;
	WX5970<=WX5907 and RESET;
	WX5972<=WX5909 and RESET;
	WX5974<=WX5911 and RESET;
	WX5976<=WX5913 and RESET;
	WX5978<=WX5915 and RESET;
	WX5980<=WX5917 and RESET;
	WX5982<=WX5919 and RESET;
	WX5984<=WX5921 and RESET;
	WX5986<=WX5923 and RESET;
	WX5988<=WX5925 and RESET;
	WX5990<=WX5927 and RESET;
	WX5992<=WX5929 and RESET;
	WX5994<=WX5931 and RESET;
	WX5996<=WX5933 and RESET;
	WX5998<=WX5935 and RESET;
	WX6000<=WX5937 and RESET;
	WX6002<=WX5939 and RESET;
	WX6004<=WX5941 and RESET;
	WX6006<=WX5943 and RESET;
	WX6008<=WX5945 and RESET;
	WX6010<=WX5947 and RESET;
	WX6012<=WX5949 and RESET;
	WX6014<=WX5951 and RESET;
	WX6016<=WX5953 and RESET;
	WX6018<=WX5955 and RESET;
	WX6020<=WX5957 and RESET;
	WX6022<=WX5959 and RESET;
	WX6024<=WX5961 and RESET;
	WX6026<=WX5963 and RESET;
	WX6028<=WX5965 and RESET;
	WX6030<=WX5967 and RESET;
	WX6032<=WX5969 and RESET;
	WX6034<=WX5971 and RESET;
	WX6036<=WX5973 and RESET;
	WX6038<=WX5975 and RESET;
	WX6040<=WX5977 and RESET;
	WX6042<=WX5979 and RESET;
	WX6044<=WX5981 and RESET;
	WX6046<=WX5983 and RESET;
	WX6048<=WX5985 and RESET;
	WX6050<=WX5987 and RESET;
	WX6052<=WX5989 and RESET;
	WX6054<=WX5991 and RESET;
	WX6056<=WX5993 and RESET;
	WX6058<=WX5995 and RESET;
	WX6060<=WX5997 and RESET;
	WX6062<=WX5999 and RESET;
	WX6064<=WX6001 and RESET;
	WX6066<=WX6003 and RESET;
	WX6068<=WX6005 and RESET;
	WX6070<=WX6007 and RESET;
	WX6179<=WX6178 and WX6177;
	WX6180<=WX5752 and WX6181;
	WX6186<=WX6185 and WX6177;
	WX6187<=WX5753 and WX6188;
	WX6193<=WX6192 and WX6177;
	WX6194<=WX5754 and WX6195;
	WX6200<=WX6199 and WX6177;
	WX6201<=WX5755 and WX6202;
	WX6207<=WX6206 and WX6177;
	WX6208<=WX5756 and WX6209;
	WX6214<=WX6213 and WX6177;
	WX6215<=WX5757 and WX6216;
	WX6221<=WX6220 and WX6177;
	WX6222<=WX5758 and WX6223;
	WX6228<=WX6227 and WX6177;
	WX6229<=WX5759 and WX6230;
	WX6235<=WX6234 and WX6177;
	WX6236<=WX5760 and WX6237;
	WX6242<=WX6241 and WX6177;
	WX6243<=WX5761 and WX6244;
	WX6249<=WX6248 and WX6177;
	WX6250<=WX5762 and WX6251;
	WX6256<=WX6255 and WX6177;
	WX6257<=WX5763 and WX6258;
	WX6263<=WX6262 and WX6177;
	WX6264<=WX5764 and WX6265;
	WX6270<=WX6269 and WX6177;
	WX6271<=WX5765 and WX6272;
	WX6277<=WX6276 and WX6177;
	WX6278<=WX5766 and WX6279;
	WX6284<=WX6283 and WX6177;
	WX6285<=WX5767 and WX6286;
	WX6291<=WX6290 and WX6177;
	WX6292<=WX5768 and WX6293;
	WX6298<=WX6297 and WX6177;
	WX6299<=WX5769 and WX6300;
	WX6305<=WX6304 and WX6177;
	WX6306<=WX5770 and WX6307;
	WX6312<=WX6311 and WX6177;
	WX6313<=WX5771 and WX6314;
	WX6319<=WX6318 and WX6177;
	WX6320<=WX5772 and WX6321;
	WX6326<=WX6325 and WX6177;
	WX6327<=WX5773 and WX6328;
	WX6333<=WX6332 and WX6177;
	WX6334<=WX5774 and WX6335;
	WX6340<=WX6339 and WX6177;
	WX6341<=WX5775 and WX6342;
	WX6347<=WX6346 and WX6177;
	WX6348<=WX5776 and WX6349;
	WX6354<=WX6353 and WX6177;
	WX6355<=WX5777 and WX6356;
	WX6361<=WX6360 and WX6177;
	WX6362<=WX5778 and WX6363;
	WX6368<=WX6367 and WX6177;
	WX6369<=WX5779 and WX6370;
	WX6375<=WX6374 and WX6177;
	WX6376<=WX5780 and WX6377;
	WX6382<=WX6381 and WX6177;
	WX6383<=WX5781 and WX6384;
	WX6389<=WX6388 and WX6177;
	WX6390<=WX5782 and WX6391;
	WX6396<=WX6395 and WX6177;
	WX6397<=WX5783 and WX6398;
	WX6436<=WX6406 and WX6435;
	WX6438<=WX6434 and WX6435;
	WX6440<=WX6433 and WX6435;
	WX6442<=WX6432 and WX6435;
	WX6444<=WX6405 and WX6435;
	WX6446<=WX6431 and WX6435;
	WX6448<=WX6430 and WX6435;
	WX6450<=WX6429 and WX6435;
	WX6452<=WX6428 and WX6435;
	WX6454<=WX6427 and WX6435;
	WX6456<=WX6426 and WX6435;
	WX6458<=WX6404 and WX6435;
	WX6460<=WX6425 and WX6435;
	WX6462<=WX6424 and WX6435;
	WX6464<=WX6423 and WX6435;
	WX6466<=WX6422 and WX6435;
	WX6468<=WX6403 and WX6435;
	WX6470<=WX6421 and WX6435;
	WX6472<=WX6420 and WX6435;
	WX6474<=WX6419 and WX6435;
	WX6476<=WX6418 and WX6435;
	WX6478<=WX6417 and WX6435;
	WX6480<=WX6416 and WX6435;
	WX6482<=WX6415 and WX6435;
	WX6484<=WX6414 and WX6435;
	WX6486<=WX6413 and WX6435;
	WX6488<=WX6412 and WX6435;
	WX6490<=WX6411 and WX6435;
	WX6492<=WX6410 and WX6435;
	WX6494<=WX6409 and WX6435;
	WX6496<=WX6408 and WX6435;
	WX6498<=WX6407 and WX6435;
	WX6500<=WX6511 and WX7468;
	WX6501<=WX6507 and WX6502;
	WX6504<=CRC_OUT_4_31 and WX7469;
	WX6505<=WX8770 and WX6506;
	WX6508<=WX6950 and WX7469;
	WX6509<=WX7477 and WX6510;
	WX6514<=WX6525 and WX7468;
	WX6515<=WX6521 and WX6516;
	WX6518<=CRC_OUT_4_30 and WX7469;
	WX6519<=WX8777 and WX6520;
	WX6522<=WX6952 and WX7469;
	WX6523<=WX7484 and WX6524;
	WX6528<=WX6539 and WX7468;
	WX6529<=WX6535 and WX6530;
	WX6532<=CRC_OUT_4_29 and WX7469;
	WX6533<=WX8784 and WX6534;
	WX6536<=WX6954 and WX7469;
	WX6537<=WX7491 and WX6538;
	WX6542<=WX6553 and WX7468;
	WX6543<=WX6549 and WX6544;
	WX6546<=CRC_OUT_4_28 and WX7469;
	WX6547<=WX8791 and WX6548;
	WX6550<=WX6956 and WX7469;
	WX6551<=WX7498 and WX6552;
	WX6556<=WX6567 and WX7468;
	WX6557<=WX6563 and WX6558;
	WX6560<=CRC_OUT_4_27 and WX7469;
	WX6561<=WX8798 and WX6562;
	WX6564<=WX6958 and WX7469;
	WX6565<=WX7505 and WX6566;
	WX6570<=WX6581 and WX7468;
	WX6571<=WX6577 and WX6572;
	WX6574<=CRC_OUT_4_26 and WX7469;
	WX6575<=WX8805 and WX6576;
	WX6578<=WX6960 and WX7469;
	WX6579<=WX7512 and WX6580;
	WX6584<=WX6595 and WX7468;
	WX6585<=WX6591 and WX6586;
	WX6588<=CRC_OUT_4_25 and WX7469;
	WX6589<=WX8812 and WX6590;
	WX6592<=WX6962 and WX7469;
	WX6593<=WX7519 and WX6594;
	WX6598<=WX6609 and WX7468;
	WX6599<=WX6605 and WX6600;
	WX6602<=CRC_OUT_4_24 and WX7469;
	WX6603<=WX8819 and WX6604;
	WX6606<=WX6964 and WX7469;
	WX6607<=WX7526 and WX6608;
	WX6612<=WX6623 and WX7468;
	WX6613<=WX6619 and WX6614;
	WX6616<=CRC_OUT_4_23 and WX7469;
	WX6617<=WX8826 and WX6618;
	WX6620<=WX6966 and WX7469;
	WX6621<=WX7533 and WX6622;
	WX6626<=WX6637 and WX7468;
	WX6627<=WX6633 and WX6628;
	WX6630<=CRC_OUT_4_22 and WX7469;
	WX6631<=WX8833 and WX6632;
	WX6634<=WX6968 and WX7469;
	WX6635<=WX7540 and WX6636;
	WX6640<=WX6651 and WX7468;
	WX6641<=WX6647 and WX6642;
	WX6644<=CRC_OUT_4_21 and WX7469;
	WX6645<=WX8840 and WX6646;
	WX6648<=WX6970 and WX7469;
	WX6649<=WX7547 and WX6650;
	WX6654<=WX6665 and WX7468;
	WX6655<=WX6661 and WX6656;
	WX6658<=CRC_OUT_4_20 and WX7469;
	WX6659<=WX8847 and WX6660;
	WX6662<=WX6972 and WX7469;
	WX6663<=WX7554 and WX6664;
	WX6668<=WX6679 and WX7468;
	WX6669<=WX6675 and WX6670;
	WX6672<=CRC_OUT_4_19 and WX7469;
	WX6673<=WX8854 and WX6674;
	WX6676<=WX6974 and WX7469;
	WX6677<=WX7561 and WX6678;
	WX6682<=WX6693 and WX7468;
	WX6683<=WX6689 and WX6684;
	WX6686<=CRC_OUT_4_18 and WX7469;
	WX6687<=WX8861 and WX6688;
	WX6690<=WX6976 and WX7469;
	WX6691<=WX7568 and WX6692;
	WX6696<=WX6707 and WX7468;
	WX6697<=WX6703 and WX6698;
	WX6700<=CRC_OUT_4_17 and WX7469;
	WX6701<=WX8868 and WX6702;
	WX6704<=WX6978 and WX7469;
	WX6705<=WX7575 and WX6706;
	WX6710<=WX6721 and WX7468;
	WX6711<=WX6717 and WX6712;
	WX6714<=CRC_OUT_4_16 and WX7469;
	WX6715<=WX8875 and WX6716;
	WX6718<=WX6980 and WX7469;
	WX6719<=WX7582 and WX6720;
	WX6724<=WX6735 and WX7468;
	WX6725<=WX6731 and WX6726;
	WX6728<=CRC_OUT_4_15 and WX7469;
	WX6729<=WX8882 and WX6730;
	WX6732<=WX6982 and WX7469;
	WX6733<=WX7589 and WX6734;
	WX6738<=WX6749 and WX7468;
	WX6739<=WX6745 and WX6740;
	WX6742<=CRC_OUT_4_14 and WX7469;
	WX6743<=WX8889 and WX6744;
	WX6746<=WX6984 and WX7469;
	WX6747<=WX7596 and WX6748;
	WX6752<=WX6763 and WX7468;
	WX6753<=WX6759 and WX6754;
	WX6756<=CRC_OUT_4_13 and WX7469;
	WX6757<=WX8896 and WX6758;
	WX6760<=WX6986 and WX7469;
	WX6761<=WX7603 and WX6762;
	WX6766<=WX6777 and WX7468;
	WX6767<=WX6773 and WX6768;
	WX6770<=CRC_OUT_4_12 and WX7469;
	WX6771<=WX8903 and WX6772;
	WX6774<=WX6988 and WX7469;
	WX6775<=WX7610 and WX6776;
	WX6780<=WX6791 and WX7468;
	WX6781<=WX6787 and WX6782;
	WX6784<=CRC_OUT_4_11 and WX7469;
	WX6785<=WX8910 and WX6786;
	WX6788<=WX6990 and WX7469;
	WX6789<=WX7617 and WX6790;
	WX6794<=WX6805 and WX7468;
	WX6795<=WX6801 and WX6796;
	WX6798<=CRC_OUT_4_10 and WX7469;
	WX6799<=WX8917 and WX6800;
	WX6802<=WX6992 and WX7469;
	WX6803<=WX7624 and WX6804;
	WX6808<=WX6819 and WX7468;
	WX6809<=WX6815 and WX6810;
	WX6812<=CRC_OUT_4_9 and WX7469;
	WX6813<=WX8924 and WX6814;
	WX6816<=WX6994 and WX7469;
	WX6817<=WX7631 and WX6818;
	WX6822<=WX6833 and WX7468;
	WX6823<=WX6829 and WX6824;
	WX6826<=CRC_OUT_4_8 and WX7469;
	WX6827<=WX8931 and WX6828;
	WX6830<=WX6996 and WX7469;
	WX6831<=WX7638 and WX6832;
	WX6836<=WX6847 and WX7468;
	WX6837<=WX6843 and WX6838;
	WX6840<=CRC_OUT_4_7 and WX7469;
	WX6841<=WX8938 and WX6842;
	WX6844<=WX6998 and WX7469;
	WX6845<=WX7645 and WX6846;
	WX6850<=WX6861 and WX7468;
	WX6851<=WX6857 and WX6852;
	WX6854<=CRC_OUT_4_6 and WX7469;
	WX6855<=WX8945 and WX6856;
	WX6858<=WX7000 and WX7469;
	WX6859<=WX7652 and WX6860;
	WX6864<=WX6875 and WX7468;
	WX6865<=WX6871 and WX6866;
	WX6868<=CRC_OUT_4_5 and WX7469;
	WX6869<=WX8952 and WX6870;
	WX6872<=WX7002 and WX7469;
	WX6873<=WX7659 and WX6874;
	WX6878<=WX6889 and WX7468;
	WX6879<=WX6885 and WX6880;
	WX6882<=CRC_OUT_4_4 and WX7469;
	WX6883<=WX8959 and WX6884;
	WX6886<=WX7004 and WX7469;
	WX6887<=WX7666 and WX6888;
	WX6892<=WX6903 and WX7468;
	WX6893<=WX6899 and WX6894;
	WX6896<=CRC_OUT_4_3 and WX7469;
	WX6897<=WX8966 and WX6898;
	WX6900<=WX7006 and WX7469;
	WX6901<=WX7673 and WX6902;
	WX6906<=WX6917 and WX7468;
	WX6907<=WX6913 and WX6908;
	WX6910<=CRC_OUT_4_2 and WX7469;
	WX6911<=WX8973 and WX6912;
	WX6914<=WX7008 and WX7469;
	WX6915<=WX7680 and WX6916;
	WX6920<=WX6931 and WX7468;
	WX6921<=WX6927 and WX6922;
	WX6924<=CRC_OUT_4_1 and WX7469;
	WX6925<=WX8980 and WX6926;
	WX6928<=WX7010 and WX7469;
	WX6929<=WX7687 and WX6930;
	WX6934<=WX6945 and WX7468;
	WX6935<=WX6941 and WX6936;
	WX6938<=CRC_OUT_4_0 and WX7469;
	WX6939<=WX8987 and WX6940;
	WX6942<=WX7012 and WX7469;
	WX6943<=WX7694 and WX6944;
	WX6949<=WX6952 and RESET;
	WX6951<=WX6954 and RESET;
	WX6953<=WX6956 and RESET;
	WX6955<=WX6958 and RESET;
	WX6957<=WX6960 and RESET;
	WX6959<=WX6962 and RESET;
	WX6961<=WX6964 and RESET;
	WX6963<=WX6966 and RESET;
	WX6965<=WX6968 and RESET;
	WX6967<=WX6970 and RESET;
	WX6969<=WX6972 and RESET;
	WX6971<=WX6974 and RESET;
	WX6973<=WX6976 and RESET;
	WX6975<=WX6978 and RESET;
	WX6977<=WX6980 and RESET;
	WX6979<=WX6982 and RESET;
	WX6981<=WX6984 and RESET;
	WX6983<=WX6986 and RESET;
	WX6985<=WX6988 and RESET;
	WX6987<=WX6990 and RESET;
	WX6989<=WX6992 and RESET;
	WX6991<=WX6994 and RESET;
	WX6993<=WX6996 and RESET;
	WX6995<=WX6998 and RESET;
	WX6997<=WX7000 and RESET;
	WX6999<=WX7002 and RESET;
	WX7001<=WX7004 and RESET;
	WX7003<=WX7006 and RESET;
	WX7005<=WX7008 and RESET;
	WX7007<=WX7010 and RESET;
	WX7009<=WX7012 and RESET;
	WX7011<=WX6948 and RESET;
	WX7109<=WX6513 and RESET;
	WX7111<=WX6527 and RESET;
	WX7113<=WX6541 and RESET;
	WX7115<=WX6555 and RESET;
	WX7117<=WX6569 and RESET;
	WX7119<=WX6583 and RESET;
	WX7121<=WX6597 and RESET;
	WX7123<=WX6611 and RESET;
	WX7125<=WX6625 and RESET;
	WX7127<=WX6639 and RESET;
	WX7129<=WX6653 and RESET;
	WX7131<=WX6667 and RESET;
	WX7133<=WX6681 and RESET;
	WX7135<=WX6695 and RESET;
	WX7137<=WX6709 and RESET;
	WX7139<=WX6723 and RESET;
	WX7141<=WX6737 and RESET;
	WX7143<=WX6751 and RESET;
	WX7145<=WX6765 and RESET;
	WX7147<=WX6779 and RESET;
	WX7149<=WX6793 and RESET;
	WX7151<=WX6807 and RESET;
	WX7153<=WX6821 and RESET;
	WX7155<=WX6835 and RESET;
	WX7157<=WX6849 and RESET;
	WX7159<=WX6863 and RESET;
	WX7161<=WX6877 and RESET;
	WX7163<=WX6891 and RESET;
	WX7165<=WX6905 and RESET;
	WX7167<=WX6919 and RESET;
	WX7169<=WX6933 and RESET;
	WX7171<=WX6947 and RESET;
	WX7173<=WX7110 and RESET;
	WX7175<=WX7112 and RESET;
	WX7177<=WX7114 and RESET;
	WX7179<=WX7116 and RESET;
	WX7181<=WX7118 and RESET;
	WX7183<=WX7120 and RESET;
	WX7185<=WX7122 and RESET;
	WX7187<=WX7124 and RESET;
	WX7189<=WX7126 and RESET;
	WX7191<=WX7128 and RESET;
	WX7193<=WX7130 and RESET;
	WX7195<=WX7132 and RESET;
	WX7197<=WX7134 and RESET;
	WX7199<=WX7136 and RESET;
	WX7201<=WX7138 and RESET;
	WX7203<=WX7140 and RESET;
	WX7205<=WX7142 and RESET;
	WX7207<=WX7144 and RESET;
	WX7209<=WX7146 and RESET;
	WX7211<=WX7148 and RESET;
	WX7213<=WX7150 and RESET;
	WX7215<=WX7152 and RESET;
	WX7217<=WX7154 and RESET;
	WX7219<=WX7156 and RESET;
	WX7221<=WX7158 and RESET;
	WX7223<=WX7160 and RESET;
	WX7225<=WX7162 and RESET;
	WX7227<=WX7164 and RESET;
	WX7229<=WX7166 and RESET;
	WX7231<=WX7168 and RESET;
	WX7233<=WX7170 and RESET;
	WX7235<=WX7172 and RESET;
	WX7237<=WX7174 and RESET;
	WX7239<=WX7176 and RESET;
	WX7241<=WX7178 and RESET;
	WX7243<=WX7180 and RESET;
	WX7245<=WX7182 and RESET;
	WX7247<=WX7184 and RESET;
	WX7249<=WX7186 and RESET;
	WX7251<=WX7188 and RESET;
	WX7253<=WX7190 and RESET;
	WX7255<=WX7192 and RESET;
	WX7257<=WX7194 and RESET;
	WX7259<=WX7196 and RESET;
	WX7261<=WX7198 and RESET;
	WX7263<=WX7200 and RESET;
	WX7265<=WX7202 and RESET;
	WX7267<=WX7204 and RESET;
	WX7269<=WX7206 and RESET;
	WX7271<=WX7208 and RESET;
	WX7273<=WX7210 and RESET;
	WX7275<=WX7212 and RESET;
	WX7277<=WX7214 and RESET;
	WX7279<=WX7216 and RESET;
	WX7281<=WX7218 and RESET;
	WX7283<=WX7220 and RESET;
	WX7285<=WX7222 and RESET;
	WX7287<=WX7224 and RESET;
	WX7289<=WX7226 and RESET;
	WX7291<=WX7228 and RESET;
	WX7293<=WX7230 and RESET;
	WX7295<=WX7232 and RESET;
	WX7297<=WX7234 and RESET;
	WX7299<=WX7236 and RESET;
	WX7301<=WX7238 and RESET;
	WX7303<=WX7240 and RESET;
	WX7305<=WX7242 and RESET;
	WX7307<=WX7244 and RESET;
	WX7309<=WX7246 and RESET;
	WX7311<=WX7248 and RESET;
	WX7313<=WX7250 and RESET;
	WX7315<=WX7252 and RESET;
	WX7317<=WX7254 and RESET;
	WX7319<=WX7256 and RESET;
	WX7321<=WX7258 and RESET;
	WX7323<=WX7260 and RESET;
	WX7325<=WX7262 and RESET;
	WX7327<=WX7264 and RESET;
	WX7329<=WX7266 and RESET;
	WX7331<=WX7268 and RESET;
	WX7333<=WX7270 and RESET;
	WX7335<=WX7272 and RESET;
	WX7337<=WX7274 and RESET;
	WX7339<=WX7276 and RESET;
	WX7341<=WX7278 and RESET;
	WX7343<=WX7280 and RESET;
	WX7345<=WX7282 and RESET;
	WX7347<=WX7284 and RESET;
	WX7349<=WX7286 and RESET;
	WX7351<=WX7288 and RESET;
	WX7353<=WX7290 and RESET;
	WX7355<=WX7292 and RESET;
	WX7357<=WX7294 and RESET;
	WX7359<=WX7296 and RESET;
	WX7361<=WX7298 and RESET;
	WX7363<=WX7300 and RESET;
	WX7472<=WX7471 and WX7470;
	WX7473<=WX7045 and WX7474;
	WX7479<=WX7478 and WX7470;
	WX7480<=WX7046 and WX7481;
	WX7486<=WX7485 and WX7470;
	WX7487<=WX7047 and WX7488;
	WX7493<=WX7492 and WX7470;
	WX7494<=WX7048 and WX7495;
	WX7500<=WX7499 and WX7470;
	WX7501<=WX7049 and WX7502;
	WX7507<=WX7506 and WX7470;
	WX7508<=WX7050 and WX7509;
	WX7514<=WX7513 and WX7470;
	WX7515<=WX7051 and WX7516;
	WX7521<=WX7520 and WX7470;
	WX7522<=WX7052 and WX7523;
	WX7528<=WX7527 and WX7470;
	WX7529<=WX7053 and WX7530;
	WX7535<=WX7534 and WX7470;
	WX7536<=WX7054 and WX7537;
	WX7542<=WX7541 and WX7470;
	WX7543<=WX7055 and WX7544;
	WX7549<=WX7548 and WX7470;
	WX7550<=WX7056 and WX7551;
	WX7556<=WX7555 and WX7470;
	WX7557<=WX7057 and WX7558;
	WX7563<=WX7562 and WX7470;
	WX7564<=WX7058 and WX7565;
	WX7570<=WX7569 and WX7470;
	WX7571<=WX7059 and WX7572;
	WX7577<=WX7576 and WX7470;
	WX7578<=WX7060 and WX7579;
	WX7584<=WX7583 and WX7470;
	WX7585<=WX7061 and WX7586;
	WX7591<=WX7590 and WX7470;
	WX7592<=WX7062 and WX7593;
	WX7598<=WX7597 and WX7470;
	WX7599<=WX7063 and WX7600;
	WX7605<=WX7604 and WX7470;
	WX7606<=WX7064 and WX7607;
	WX7612<=WX7611 and WX7470;
	WX7613<=WX7065 and WX7614;
	WX7619<=WX7618 and WX7470;
	WX7620<=WX7066 and WX7621;
	WX7626<=WX7625 and WX7470;
	WX7627<=WX7067 and WX7628;
	WX7633<=WX7632 and WX7470;
	WX7634<=WX7068 and WX7635;
	WX7640<=WX7639 and WX7470;
	WX7641<=WX7069 and WX7642;
	WX7647<=WX7646 and WX7470;
	WX7648<=WX7070 and WX7649;
	WX7654<=WX7653 and WX7470;
	WX7655<=WX7071 and WX7656;
	WX7661<=WX7660 and WX7470;
	WX7662<=WX7072 and WX7663;
	WX7668<=WX7667 and WX7470;
	WX7669<=WX7073 and WX7670;
	WX7675<=WX7674 and WX7470;
	WX7676<=WX7074 and WX7677;
	WX7682<=WX7681 and WX7470;
	WX7683<=WX7075 and WX7684;
	WX7689<=WX7688 and WX7470;
	WX7690<=WX7076 and WX7691;
	WX7729<=WX7699 and WX7728;
	WX7731<=WX7727 and WX7728;
	WX7733<=WX7726 and WX7728;
	WX7735<=WX7725 and WX7728;
	WX7737<=WX7698 and WX7728;
	WX7739<=WX7724 and WX7728;
	WX7741<=WX7723 and WX7728;
	WX7743<=WX7722 and WX7728;
	WX7745<=WX7721 and WX7728;
	WX7747<=WX7720 and WX7728;
	WX7749<=WX7719 and WX7728;
	WX7751<=WX7697 and WX7728;
	WX7753<=WX7718 and WX7728;
	WX7755<=WX7717 and WX7728;
	WX7757<=WX7716 and WX7728;
	WX7759<=WX7715 and WX7728;
	WX7761<=WX7696 and WX7728;
	WX7763<=WX7714 and WX7728;
	WX7765<=WX7713 and WX7728;
	WX7767<=WX7712 and WX7728;
	WX7769<=WX7711 and WX7728;
	WX7771<=WX7710 and WX7728;
	WX7773<=WX7709 and WX7728;
	WX7775<=WX7708 and WX7728;
	WX7777<=WX7707 and WX7728;
	WX7779<=WX7706 and WX7728;
	WX7781<=WX7705 and WX7728;
	WX7783<=WX7704 and WX7728;
	WX7785<=WX7703 and WX7728;
	WX7787<=WX7702 and WX7728;
	WX7789<=WX7701 and WX7728;
	WX7791<=WX7700 and WX7728;
	WX7793<=WX7804 and WX8761;
	WX7794<=WX7800 and WX7795;
	WX7797<=CRC_OUT_3_31 and WX8762;
	WX7798<=WX10063 and WX7799;
	WX7801<=WX8243 and WX8762;
	WX7802<=WX8770 and WX7803;
	WX7807<=WX7818 and WX8761;
	WX7808<=WX7814 and WX7809;
	WX7811<=CRC_OUT_3_30 and WX8762;
	WX7812<=WX10070 and WX7813;
	WX7815<=WX8245 and WX8762;
	WX7816<=WX8777 and WX7817;
	WX7821<=WX7832 and WX8761;
	WX7822<=WX7828 and WX7823;
	WX7825<=CRC_OUT_3_29 and WX8762;
	WX7826<=WX10077 and WX7827;
	WX7829<=WX8247 and WX8762;
	WX7830<=WX8784 and WX7831;
	WX7835<=WX7846 and WX8761;
	WX7836<=WX7842 and WX7837;
	WX7839<=CRC_OUT_3_28 and WX8762;
	WX7840<=WX10084 and WX7841;
	WX7843<=WX8249 and WX8762;
	WX7844<=WX8791 and WX7845;
	WX7849<=WX7860 and WX8761;
	WX7850<=WX7856 and WX7851;
	WX7853<=CRC_OUT_3_27 and WX8762;
	WX7854<=WX10091 and WX7855;
	WX7857<=WX8251 and WX8762;
	WX7858<=WX8798 and WX7859;
	WX7863<=WX7874 and WX8761;
	WX7864<=WX7870 and WX7865;
	WX7867<=CRC_OUT_3_26 and WX8762;
	WX7868<=WX10098 and WX7869;
	WX7871<=WX8253 and WX8762;
	WX7872<=WX8805 and WX7873;
	WX7877<=WX7888 and WX8761;
	WX7878<=WX7884 and WX7879;
	WX7881<=CRC_OUT_3_25 and WX8762;
	WX7882<=WX10105 and WX7883;
	WX7885<=WX8255 and WX8762;
	WX7886<=WX8812 and WX7887;
	WX7891<=WX7902 and WX8761;
	WX7892<=WX7898 and WX7893;
	WX7895<=CRC_OUT_3_24 and WX8762;
	WX7896<=WX10112 and WX7897;
	WX7899<=WX8257 and WX8762;
	WX7900<=WX8819 and WX7901;
	WX7905<=WX7916 and WX8761;
	WX7906<=WX7912 and WX7907;
	WX7909<=CRC_OUT_3_23 and WX8762;
	WX7910<=WX10119 and WX7911;
	WX7913<=WX8259 and WX8762;
	WX7914<=WX8826 and WX7915;
	WX7919<=WX7930 and WX8761;
	WX7920<=WX7926 and WX7921;
	WX7923<=CRC_OUT_3_22 and WX8762;
	WX7924<=WX10126 and WX7925;
	WX7927<=WX8261 and WX8762;
	WX7928<=WX8833 and WX7929;
	WX7933<=WX7944 and WX8761;
	WX7934<=WX7940 and WX7935;
	WX7937<=CRC_OUT_3_21 and WX8762;
	WX7938<=WX10133 and WX7939;
	WX7941<=WX8263 and WX8762;
	WX7942<=WX8840 and WX7943;
	WX7947<=WX7958 and WX8761;
	WX7948<=WX7954 and WX7949;
	WX7951<=CRC_OUT_3_20 and WX8762;
	WX7952<=WX10140 and WX7953;
	WX7955<=WX8265 and WX8762;
	WX7956<=WX8847 and WX7957;
	WX7961<=WX7972 and WX8761;
	WX7962<=WX7968 and WX7963;
	WX7965<=CRC_OUT_3_19 and WX8762;
	WX7966<=WX10147 and WX7967;
	WX7969<=WX8267 and WX8762;
	WX7970<=WX8854 and WX7971;
	WX7975<=WX7986 and WX8761;
	WX7976<=WX7982 and WX7977;
	WX7979<=CRC_OUT_3_18 and WX8762;
	WX7980<=WX10154 and WX7981;
	WX7983<=WX8269 and WX8762;
	WX7984<=WX8861 and WX7985;
	WX7989<=WX8000 and WX8761;
	WX7990<=WX7996 and WX7991;
	WX7993<=CRC_OUT_3_17 and WX8762;
	WX7994<=WX10161 and WX7995;
	WX7997<=WX8271 and WX8762;
	WX7998<=WX8868 and WX7999;
	WX8003<=WX8014 and WX8761;
	WX8004<=WX8010 and WX8005;
	WX8007<=CRC_OUT_3_16 and WX8762;
	WX8008<=WX10168 and WX8009;
	WX8011<=WX8273 and WX8762;
	WX8012<=WX8875 and WX8013;
	WX8017<=WX8028 and WX8761;
	WX8018<=WX8024 and WX8019;
	WX8021<=CRC_OUT_3_15 and WX8762;
	WX8022<=WX10175 and WX8023;
	WX8025<=WX8275 and WX8762;
	WX8026<=WX8882 and WX8027;
	WX8031<=WX8042 and WX8761;
	WX8032<=WX8038 and WX8033;
	WX8035<=CRC_OUT_3_14 and WX8762;
	WX8036<=WX10182 and WX8037;
	WX8039<=WX8277 and WX8762;
	WX8040<=WX8889 and WX8041;
	WX8045<=WX8056 and WX8761;
	WX8046<=WX8052 and WX8047;
	WX8049<=CRC_OUT_3_13 and WX8762;
	WX8050<=WX10189 and WX8051;
	WX8053<=WX8279 and WX8762;
	WX8054<=WX8896 and WX8055;
	WX8059<=WX8070 and WX8761;
	WX8060<=WX8066 and WX8061;
	WX8063<=CRC_OUT_3_12 and WX8762;
	WX8064<=WX10196 and WX8065;
	WX8067<=WX8281 and WX8762;
	WX8068<=WX8903 and WX8069;
	WX8073<=WX8084 and WX8761;
	WX8074<=WX8080 and WX8075;
	WX8077<=CRC_OUT_3_11 and WX8762;
	WX8078<=WX10203 and WX8079;
	WX8081<=WX8283 and WX8762;
	WX8082<=WX8910 and WX8083;
	WX8087<=WX8098 and WX8761;
	WX8088<=WX8094 and WX8089;
	WX8091<=CRC_OUT_3_10 and WX8762;
	WX8092<=WX10210 and WX8093;
	WX8095<=WX8285 and WX8762;
	WX8096<=WX8917 and WX8097;
	WX8101<=WX8112 and WX8761;
	WX8102<=WX8108 and WX8103;
	WX8105<=CRC_OUT_3_9 and WX8762;
	WX8106<=WX10217 and WX8107;
	WX8109<=WX8287 and WX8762;
	WX8110<=WX8924 and WX8111;
	WX8115<=WX8126 and WX8761;
	WX8116<=WX8122 and WX8117;
	WX8119<=CRC_OUT_3_8 and WX8762;
	WX8120<=WX10224 and WX8121;
	WX8123<=WX8289 and WX8762;
	WX8124<=WX8931 and WX8125;
	WX8129<=WX8140 and WX8761;
	WX8130<=WX8136 and WX8131;
	WX8133<=CRC_OUT_3_7 and WX8762;
	WX8134<=WX10231 and WX8135;
	WX8137<=WX8291 and WX8762;
	WX8138<=WX8938 and WX8139;
	WX8143<=WX8154 and WX8761;
	WX8144<=WX8150 and WX8145;
	WX8147<=CRC_OUT_3_6 and WX8762;
	WX8148<=WX10238 and WX8149;
	WX8151<=WX8293 and WX8762;
	WX8152<=WX8945 and WX8153;
	WX8157<=WX8168 and WX8761;
	WX8158<=WX8164 and WX8159;
	WX8161<=CRC_OUT_3_5 and WX8762;
	WX8162<=WX10245 and WX8163;
	WX8165<=WX8295 and WX8762;
	WX8166<=WX8952 and WX8167;
	WX8171<=WX8182 and WX8761;
	WX8172<=WX8178 and WX8173;
	WX8175<=CRC_OUT_3_4 and WX8762;
	WX8176<=WX10252 and WX8177;
	WX8179<=WX8297 and WX8762;
	WX8180<=WX8959 and WX8181;
	WX8185<=WX8196 and WX8761;
	WX8186<=WX8192 and WX8187;
	WX8189<=CRC_OUT_3_3 and WX8762;
	WX8190<=WX10259 and WX8191;
	WX8193<=WX8299 and WX8762;
	WX8194<=WX8966 and WX8195;
	WX8199<=WX8210 and WX8761;
	WX8200<=WX8206 and WX8201;
	WX8203<=CRC_OUT_3_2 and WX8762;
	WX8204<=WX10266 and WX8205;
	WX8207<=WX8301 and WX8762;
	WX8208<=WX8973 and WX8209;
	WX8213<=WX8224 and WX8761;
	WX8214<=WX8220 and WX8215;
	WX8217<=CRC_OUT_3_1 and WX8762;
	WX8218<=WX10273 and WX8219;
	WX8221<=WX8303 and WX8762;
	WX8222<=WX8980 and WX8223;
	WX8227<=WX8238 and WX8761;
	WX8228<=WX8234 and WX8229;
	WX8231<=CRC_OUT_3_0 and WX8762;
	WX8232<=WX10280 and WX8233;
	WX8235<=WX8305 and WX8762;
	WX8236<=WX8987 and WX8237;
	WX8242<=WX8245 and RESET;
	WX8244<=WX8247 and RESET;
	WX8246<=WX8249 and RESET;
	WX8248<=WX8251 and RESET;
	WX8250<=WX8253 and RESET;
	WX8252<=WX8255 and RESET;
	WX8254<=WX8257 and RESET;
	WX8256<=WX8259 and RESET;
	WX8258<=WX8261 and RESET;
	WX8260<=WX8263 and RESET;
	WX8262<=WX8265 and RESET;
	WX8264<=WX8267 and RESET;
	WX8266<=WX8269 and RESET;
	WX8268<=WX8271 and RESET;
	WX8270<=WX8273 and RESET;
	WX8272<=WX8275 and RESET;
	WX8274<=WX8277 and RESET;
	WX8276<=WX8279 and RESET;
	WX8278<=WX8281 and RESET;
	WX8280<=WX8283 and RESET;
	WX8282<=WX8285 and RESET;
	WX8284<=WX8287 and RESET;
	WX8286<=WX8289 and RESET;
	WX8288<=WX8291 and RESET;
	WX8290<=WX8293 and RESET;
	WX8292<=WX8295 and RESET;
	WX8294<=WX8297 and RESET;
	WX8296<=WX8299 and RESET;
	WX8298<=WX8301 and RESET;
	WX8300<=WX8303 and RESET;
	WX8302<=WX8305 and RESET;
	WX8304<=WX8241 and RESET;
	WX8402<=WX7806 and RESET;
	WX8404<=WX7820 and RESET;
	WX8406<=WX7834 and RESET;
	WX8408<=WX7848 and RESET;
	WX8410<=WX7862 and RESET;
	WX8412<=WX7876 and RESET;
	WX8414<=WX7890 and RESET;
	WX8416<=WX7904 and RESET;
	WX8418<=WX7918 and RESET;
	WX8420<=WX7932 and RESET;
	WX8422<=WX7946 and RESET;
	WX8424<=WX7960 and RESET;
	WX8426<=WX7974 and RESET;
	WX8428<=WX7988 and RESET;
	WX8430<=WX8002 and RESET;
	WX8432<=WX8016 and RESET;
	WX8434<=WX8030 and RESET;
	WX8436<=WX8044 and RESET;
	WX8438<=WX8058 and RESET;
	WX8440<=WX8072 and RESET;
	WX8442<=WX8086 and RESET;
	WX8444<=WX8100 and RESET;
	WX8446<=WX8114 and RESET;
	WX8448<=WX8128 and RESET;
	WX8450<=WX8142 and RESET;
	WX8452<=WX8156 and RESET;
	WX8454<=WX8170 and RESET;
	WX8456<=WX8184 and RESET;
	WX8458<=WX8198 and RESET;
	WX8460<=WX8212 and RESET;
	WX8462<=WX8226 and RESET;
	WX8464<=WX8240 and RESET;
	WX8466<=WX8403 and RESET;
	WX8468<=WX8405 and RESET;
	WX8470<=WX8407 and RESET;
	WX8472<=WX8409 and RESET;
	WX8474<=WX8411 and RESET;
	WX8476<=WX8413 and RESET;
	WX8478<=WX8415 and RESET;
	WX8480<=WX8417 and RESET;
	WX8482<=WX8419 and RESET;
	WX8484<=WX8421 and RESET;
	WX8486<=WX8423 and RESET;
	WX8488<=WX8425 and RESET;
	WX8490<=WX8427 and RESET;
	WX8492<=WX8429 and RESET;
	WX8494<=WX8431 and RESET;
	WX8496<=WX8433 and RESET;
	WX8498<=WX8435 and RESET;
	WX8500<=WX8437 and RESET;
	WX8502<=WX8439 and RESET;
	WX8504<=WX8441 and RESET;
	WX8506<=WX8443 and RESET;
	WX8508<=WX8445 and RESET;
	WX8510<=WX8447 and RESET;
	WX8512<=WX8449 and RESET;
	WX8514<=WX8451 and RESET;
	WX8516<=WX8453 and RESET;
	WX8518<=WX8455 and RESET;
	WX8520<=WX8457 and RESET;
	WX8522<=WX8459 and RESET;
	WX8524<=WX8461 and RESET;
	WX8526<=WX8463 and RESET;
	WX8528<=WX8465 and RESET;
	WX8530<=WX8467 and RESET;
	WX8532<=WX8469 and RESET;
	WX8534<=WX8471 and RESET;
	WX8536<=WX8473 and RESET;
	WX8538<=WX8475 and RESET;
	WX8540<=WX8477 and RESET;
	WX8542<=WX8479 and RESET;
	WX8544<=WX8481 and RESET;
	WX8546<=WX8483 and RESET;
	WX8548<=WX8485 and RESET;
	WX8550<=WX8487 and RESET;
	WX8552<=WX8489 and RESET;
	WX8554<=WX8491 and RESET;
	WX8556<=WX8493 and RESET;
	WX8558<=WX8495 and RESET;
	WX8560<=WX8497 and RESET;
	WX8562<=WX8499 and RESET;
	WX8564<=WX8501 and RESET;
	WX8566<=WX8503 and RESET;
	WX8568<=WX8505 and RESET;
	WX8570<=WX8507 and RESET;
	WX8572<=WX8509 and RESET;
	WX8574<=WX8511 and RESET;
	WX8576<=WX8513 and RESET;
	WX8578<=WX8515 and RESET;
	WX8580<=WX8517 and RESET;
	WX8582<=WX8519 and RESET;
	WX8584<=WX8521 and RESET;
	WX8586<=WX8523 and RESET;
	WX8588<=WX8525 and RESET;
	WX8590<=WX8527 and RESET;
	WX8592<=WX8529 and RESET;
	WX8594<=WX8531 and RESET;
	WX8596<=WX8533 and RESET;
	WX8598<=WX8535 and RESET;
	WX8600<=WX8537 and RESET;
	WX8602<=WX8539 and RESET;
	WX8604<=WX8541 and RESET;
	WX8606<=WX8543 and RESET;
	WX8608<=WX8545 and RESET;
	WX8610<=WX8547 and RESET;
	WX8612<=WX8549 and RESET;
	WX8614<=WX8551 and RESET;
	WX8616<=WX8553 and RESET;
	WX8618<=WX8555 and RESET;
	WX8620<=WX8557 and RESET;
	WX8622<=WX8559 and RESET;
	WX8624<=WX8561 and RESET;
	WX8626<=WX8563 and RESET;
	WX8628<=WX8565 and RESET;
	WX8630<=WX8567 and RESET;
	WX8632<=WX8569 and RESET;
	WX8634<=WX8571 and RESET;
	WX8636<=WX8573 and RESET;
	WX8638<=WX8575 and RESET;
	WX8640<=WX8577 and RESET;
	WX8642<=WX8579 and RESET;
	WX8644<=WX8581 and RESET;
	WX8646<=WX8583 and RESET;
	WX8648<=WX8585 and RESET;
	WX8650<=WX8587 and RESET;
	WX8652<=WX8589 and RESET;
	WX8654<=WX8591 and RESET;
	WX8656<=WX8593 and RESET;
	WX8765<=WX8764 and WX8763;
	WX8766<=WX8338 and WX8767;
	WX8772<=WX8771 and WX8763;
	WX8773<=WX8339 and WX8774;
	WX8779<=WX8778 and WX8763;
	WX8780<=WX8340 and WX8781;
	WX8786<=WX8785 and WX8763;
	WX8787<=WX8341 and WX8788;
	WX8793<=WX8792 and WX8763;
	WX8794<=WX8342 and WX8795;
	WX8800<=WX8799 and WX8763;
	WX8801<=WX8343 and WX8802;
	WX8807<=WX8806 and WX8763;
	WX8808<=WX8344 and WX8809;
	WX8814<=WX8813 and WX8763;
	WX8815<=WX8345 and WX8816;
	WX8821<=WX8820 and WX8763;
	WX8822<=WX8346 and WX8823;
	WX8828<=WX8827 and WX8763;
	WX8829<=WX8347 and WX8830;
	WX8835<=WX8834 and WX8763;
	WX8836<=WX8348 and WX8837;
	WX8842<=WX8841 and WX8763;
	WX8843<=WX8349 and WX8844;
	WX8849<=WX8848 and WX8763;
	WX8850<=WX8350 and WX8851;
	WX8856<=WX8855 and WX8763;
	WX8857<=WX8351 and WX8858;
	WX8863<=WX8862 and WX8763;
	WX8864<=WX8352 and WX8865;
	WX8870<=WX8869 and WX8763;
	WX8871<=WX8353 and WX8872;
	WX8877<=WX8876 and WX8763;
	WX8878<=WX8354 and WX8879;
	WX8884<=WX8883 and WX8763;
	WX8885<=WX8355 and WX8886;
	WX8891<=WX8890 and WX8763;
	WX8892<=WX8356 and WX8893;
	WX8898<=WX8897 and WX8763;
	WX8899<=WX8357 and WX8900;
	WX8905<=WX8904 and WX8763;
	WX8906<=WX8358 and WX8907;
	WX8912<=WX8911 and WX8763;
	WX8913<=WX8359 and WX8914;
	WX8919<=WX8918 and WX8763;
	WX8920<=WX8360 and WX8921;
	WX8926<=WX8925 and WX8763;
	WX8927<=WX8361 and WX8928;
	WX8933<=WX8932 and WX8763;
	WX8934<=WX8362 and WX8935;
	WX8940<=WX8939 and WX8763;
	WX8941<=WX8363 and WX8942;
	WX8947<=WX8946 and WX8763;
	WX8948<=WX8364 and WX8949;
	WX8954<=WX8953 and WX8763;
	WX8955<=WX8365 and WX8956;
	WX8961<=WX8960 and WX8763;
	WX8962<=WX8366 and WX8963;
	WX8968<=WX8967 and WX8763;
	WX8969<=WX8367 and WX8970;
	WX8975<=WX8974 and WX8763;
	WX8976<=WX8368 and WX8977;
	WX8982<=WX8981 and WX8763;
	WX8983<=WX8369 and WX8984;
	WX9022<=WX8992 and WX9021;
	WX9024<=WX9020 and WX9021;
	WX9026<=WX9019 and WX9021;
	WX9028<=WX9018 and WX9021;
	WX9030<=WX8991 and WX9021;
	WX9032<=WX9017 and WX9021;
	WX9034<=WX9016 and WX9021;
	WX9036<=WX9015 and WX9021;
	WX9038<=WX9014 and WX9021;
	WX9040<=WX9013 and WX9021;
	WX9042<=WX9012 and WX9021;
	WX9044<=WX8990 and WX9021;
	WX9046<=WX9011 and WX9021;
	WX9048<=WX9010 and WX9021;
	WX9050<=WX9009 and WX9021;
	WX9052<=WX9008 and WX9021;
	WX9054<=WX8989 and WX9021;
	WX9056<=WX9007 and WX9021;
	WX9058<=WX9006 and WX9021;
	WX9060<=WX9005 and WX9021;
	WX9062<=WX9004 and WX9021;
	WX9064<=WX9003 and WX9021;
	WX9066<=WX9002 and WX9021;
	WX9068<=WX9001 and WX9021;
	WX9070<=WX9000 and WX9021;
	WX9072<=WX8999 and WX9021;
	WX9074<=WX8998 and WX9021;
	WX9076<=WX8997 and WX9021;
	WX9078<=WX8996 and WX9021;
	WX9080<=WX8995 and WX9021;
	WX9082<=WX8994 and WX9021;
	WX9084<=WX8993 and WX9021;
	WX9086<=WX9097 and WX10054;
	WX9087<=WX9093 and WX9088;
	WX9090<=CRC_OUT_2_31 and WX10055;
	WX9091<=WX11356 and WX9092;
	WX9094<=WX9536 and WX10055;
	WX9095<=WX10063 and WX9096;
	WX9100<=WX9111 and WX10054;
	WX9101<=WX9107 and WX9102;
	WX9104<=CRC_OUT_2_30 and WX10055;
	WX9105<=WX11363 and WX9106;
	WX9108<=WX9538 and WX10055;
	WX9109<=WX10070 and WX9110;
	WX9114<=WX9125 and WX10054;
	WX9115<=WX9121 and WX9116;
	WX9118<=CRC_OUT_2_29 and WX10055;
	WX9119<=WX11370 and WX9120;
	WX9122<=WX9540 and WX10055;
	WX9123<=WX10077 and WX9124;
	WX9128<=WX9139 and WX10054;
	WX9129<=WX9135 and WX9130;
	WX9132<=CRC_OUT_2_28 and WX10055;
	WX9133<=WX11377 and WX9134;
	WX9136<=WX9542 and WX10055;
	WX9137<=WX10084 and WX9138;
	WX9142<=WX9153 and WX10054;
	WX9143<=WX9149 and WX9144;
	WX9146<=CRC_OUT_2_27 and WX10055;
	WX9147<=WX11384 and WX9148;
	WX9150<=WX9544 and WX10055;
	WX9151<=WX10091 and WX9152;
	WX9156<=WX9167 and WX10054;
	WX9157<=WX9163 and WX9158;
	WX9160<=CRC_OUT_2_26 and WX10055;
	WX9161<=WX11391 and WX9162;
	WX9164<=WX9546 and WX10055;
	WX9165<=WX10098 and WX9166;
	WX9170<=WX9181 and WX10054;
	WX9171<=WX9177 and WX9172;
	WX9174<=CRC_OUT_2_25 and WX10055;
	WX9175<=WX11398 and WX9176;
	WX9178<=WX9548 and WX10055;
	WX9179<=WX10105 and WX9180;
	WX9184<=WX9195 and WX10054;
	WX9185<=WX9191 and WX9186;
	WX9188<=CRC_OUT_2_24 and WX10055;
	WX9189<=WX11405 and WX9190;
	WX9192<=WX9550 and WX10055;
	WX9193<=WX10112 and WX9194;
	WX9198<=WX9209 and WX10054;
	WX9199<=WX9205 and WX9200;
	WX9202<=CRC_OUT_2_23 and WX10055;
	WX9203<=WX11412 and WX9204;
	WX9206<=WX9552 and WX10055;
	WX9207<=WX10119 and WX9208;
	WX9212<=WX9223 and WX10054;
	WX9213<=WX9219 and WX9214;
	WX9216<=CRC_OUT_2_22 and WX10055;
	WX9217<=WX11419 and WX9218;
	WX9220<=WX9554 and WX10055;
	WX9221<=WX10126 and WX9222;
	WX9226<=WX9237 and WX10054;
	WX9227<=WX9233 and WX9228;
	WX9230<=CRC_OUT_2_21 and WX10055;
	WX9231<=WX11426 and WX9232;
	WX9234<=WX9556 and WX10055;
	WX9235<=WX10133 and WX9236;
	WX9240<=WX9251 and WX10054;
	WX9241<=WX9247 and WX9242;
	WX9244<=CRC_OUT_2_20 and WX10055;
	WX9245<=WX11433 and WX9246;
	WX9248<=WX9558 and WX10055;
	WX9249<=WX10140 and WX9250;
	WX9254<=WX9265 and WX10054;
	WX9255<=WX9261 and WX9256;
	WX9258<=CRC_OUT_2_19 and WX10055;
	WX9259<=WX11440 and WX9260;
	WX9262<=WX9560 and WX10055;
	WX9263<=WX10147 and WX9264;
	WX9268<=WX9279 and WX10054;
	WX9269<=WX9275 and WX9270;
	WX9272<=CRC_OUT_2_18 and WX10055;
	WX9273<=WX11447 and WX9274;
	WX9276<=WX9562 and WX10055;
	WX9277<=WX10154 and WX9278;
	WX9282<=WX9293 and WX10054;
	WX9283<=WX9289 and WX9284;
	WX9286<=CRC_OUT_2_17 and WX10055;
	WX9287<=WX11454 and WX9288;
	WX9290<=WX9564 and WX10055;
	WX9291<=WX10161 and WX9292;
	WX9296<=WX9307 and WX10054;
	WX9297<=WX9303 and WX9298;
	WX9300<=CRC_OUT_2_16 and WX10055;
	WX9301<=WX11461 and WX9302;
	WX9304<=WX9566 and WX10055;
	WX9305<=WX10168 and WX9306;
	WX9310<=WX9321 and WX10054;
	WX9311<=WX9317 and WX9312;
	WX9314<=CRC_OUT_2_15 and WX10055;
	WX9315<=WX11468 and WX9316;
	WX9318<=WX9568 and WX10055;
	WX9319<=WX10175 and WX9320;
	WX9324<=WX9335 and WX10054;
	WX9325<=WX9331 and WX9326;
	WX9328<=CRC_OUT_2_14 and WX10055;
	WX9329<=WX11475 and WX9330;
	WX9332<=WX9570 and WX10055;
	WX9333<=WX10182 and WX9334;
	WX9338<=WX9349 and WX10054;
	WX9339<=WX9345 and WX9340;
	WX9342<=CRC_OUT_2_13 and WX10055;
	WX9343<=WX11482 and WX9344;
	WX9346<=WX9572 and WX10055;
	WX9347<=WX10189 and WX9348;
	WX9352<=WX9363 and WX10054;
	WX9353<=WX9359 and WX9354;
	WX9356<=CRC_OUT_2_12 and WX10055;
	WX9357<=WX11489 and WX9358;
	WX9360<=WX9574 and WX10055;
	WX9361<=WX10196 and WX9362;
	WX9366<=WX9377 and WX10054;
	WX9367<=WX9373 and WX9368;
	WX9370<=CRC_OUT_2_11 and WX10055;
	WX9371<=WX11496 and WX9372;
	WX9374<=WX9576 and WX10055;
	WX9375<=WX10203 and WX9376;
	WX9380<=WX9391 and WX10054;
	WX9381<=WX9387 and WX9382;
	WX9384<=CRC_OUT_2_10 and WX10055;
	WX9385<=WX11503 and WX9386;
	WX9388<=WX9578 and WX10055;
	WX9389<=WX10210 and WX9390;
	WX9394<=WX9405 and WX10054;
	WX9395<=WX9401 and WX9396;
	WX9398<=CRC_OUT_2_9 and WX10055;
	WX9399<=WX11510 and WX9400;
	WX9402<=WX9580 and WX10055;
	WX9403<=WX10217 and WX9404;
	WX9408<=WX9419 and WX10054;
	WX9409<=WX9415 and WX9410;
	WX9412<=CRC_OUT_2_8 and WX10055;
	WX9413<=WX11517 and WX9414;
	WX9416<=WX9582 and WX10055;
	WX9417<=WX10224 and WX9418;
	WX9422<=WX9433 and WX10054;
	WX9423<=WX9429 and WX9424;
	WX9426<=CRC_OUT_2_7 and WX10055;
	WX9427<=WX11524 and WX9428;
	WX9430<=WX9584 and WX10055;
	WX9431<=WX10231 and WX9432;
	WX9436<=WX9447 and WX10054;
	WX9437<=WX9443 and WX9438;
	WX9440<=CRC_OUT_2_6 and WX10055;
	WX9441<=WX11531 and WX9442;
	WX9444<=WX9586 and WX10055;
	WX9445<=WX10238 and WX9446;
	WX9450<=WX9461 and WX10054;
	WX9451<=WX9457 and WX9452;
	WX9454<=CRC_OUT_2_5 and WX10055;
	WX9455<=WX11538 and WX9456;
	WX9458<=WX9588 and WX10055;
	WX9459<=WX10245 and WX9460;
	WX9464<=WX9475 and WX10054;
	WX9465<=WX9471 and WX9466;
	WX9468<=CRC_OUT_2_4 and WX10055;
	WX9469<=WX11545 and WX9470;
	WX9472<=WX9590 and WX10055;
	WX9473<=WX10252 and WX9474;
	WX9478<=WX9489 and WX10054;
	WX9479<=WX9485 and WX9480;
	WX9482<=CRC_OUT_2_3 and WX10055;
	WX9483<=WX11552 and WX9484;
	WX9486<=WX9592 and WX10055;
	WX9487<=WX10259 and WX9488;
	WX9492<=WX9503 and WX10054;
	WX9493<=WX9499 and WX9494;
	WX9496<=CRC_OUT_2_2 and WX10055;
	WX9497<=WX11559 and WX9498;
	WX9500<=WX9594 and WX10055;
	WX9501<=WX10266 and WX9502;
	WX9506<=WX9517 and WX10054;
	WX9507<=WX9513 and WX9508;
	WX9510<=CRC_OUT_2_1 and WX10055;
	WX9511<=WX11566 and WX9512;
	WX9514<=WX9596 and WX10055;
	WX9515<=WX10273 and WX9516;
	WX9520<=WX9531 and WX10054;
	WX9521<=WX9527 and WX9522;
	WX9524<=CRC_OUT_2_0 and WX10055;
	WX9525<=WX11573 and WX9526;
	WX9528<=WX9598 and WX10055;
	WX9529<=WX10280 and WX9530;
	WX9535<=WX9538 and RESET;
	WX9537<=WX9540 and RESET;
	WX9539<=WX9542 and RESET;
	WX9541<=WX9544 and RESET;
	WX9543<=WX9546 and RESET;
	WX9545<=WX9548 and RESET;
	WX9547<=WX9550 and RESET;
	WX9549<=WX9552 and RESET;
	WX9551<=WX9554 and RESET;
	WX9553<=WX9556 and RESET;
	WX9555<=WX9558 and RESET;
	WX9557<=WX9560 and RESET;
	WX9559<=WX9562 and RESET;
	WX9561<=WX9564 and RESET;
	WX9563<=WX9566 and RESET;
	WX9565<=WX9568 and RESET;
	WX9567<=WX9570 and RESET;
	WX9569<=WX9572 and RESET;
	WX9571<=WX9574 and RESET;
	WX9573<=WX9576 and RESET;
	WX9575<=WX9578 and RESET;
	WX9577<=WX9580 and RESET;
	WX9579<=WX9582 and RESET;
	WX9581<=WX9584 and RESET;
	WX9583<=WX9586 and RESET;
	WX9585<=WX9588 and RESET;
	WX9587<=WX9590 and RESET;
	WX9589<=WX9592 and RESET;
	WX9591<=WX9594 and RESET;
	WX9593<=WX9596 and RESET;
	WX9595<=WX9598 and RESET;
	WX9597<=WX9534 and RESET;
	WX9695<=WX9099 and RESET;
	WX9697<=WX9113 and RESET;
	WX9699<=WX9127 and RESET;
	WX9701<=WX9141 and RESET;
	WX9703<=WX9155 and RESET;
	WX9705<=WX9169 and RESET;
	WX9707<=WX9183 and RESET;
	WX9709<=WX9197 and RESET;
	WX9711<=WX9211 and RESET;
	WX9713<=WX9225 and RESET;
	WX9715<=WX9239 and RESET;
	WX9717<=WX9253 and RESET;
	WX9719<=WX9267 and RESET;
	WX9721<=WX9281 and RESET;
	WX9723<=WX9295 and RESET;
	WX9725<=WX9309 and RESET;
	WX9727<=WX9323 and RESET;
	WX9729<=WX9337 and RESET;
	WX9731<=WX9351 and RESET;
	WX9733<=WX9365 and RESET;
	WX9735<=WX9379 and RESET;
	WX9737<=WX9393 and RESET;
	WX9739<=WX9407 and RESET;
	WX9741<=WX9421 and RESET;
	WX9743<=WX9435 and RESET;
	WX9745<=WX9449 and RESET;
	WX9747<=WX9463 and RESET;
	WX9749<=WX9477 and RESET;
	WX9751<=WX9491 and RESET;
	WX9753<=WX9505 and RESET;
	WX9755<=WX9519 and RESET;
	WX9757<=WX9533 and RESET;
	WX9759<=WX9696 and RESET;
	WX9761<=WX9698 and RESET;
	WX9763<=WX9700 and RESET;
	WX9765<=WX9702 and RESET;
	WX9767<=WX9704 and RESET;
	WX9769<=WX9706 and RESET;
	WX9771<=WX9708 and RESET;
	WX9773<=WX9710 and RESET;
	WX9775<=WX9712 and RESET;
	WX9777<=WX9714 and RESET;
	WX9779<=WX9716 and RESET;
	WX9781<=WX9718 and RESET;
	WX9783<=WX9720 and RESET;
	WX9785<=WX9722 and RESET;
	WX9787<=WX9724 and RESET;
	WX9789<=WX9726 and RESET;
	WX9791<=WX9728 and RESET;
	WX9793<=WX9730 and RESET;
	WX9795<=WX9732 and RESET;
	WX9797<=WX9734 and RESET;
	WX9799<=WX9736 and RESET;
	WX9801<=WX9738 and RESET;
	WX9803<=WX9740 and RESET;
	WX9805<=WX9742 and RESET;
	WX9807<=WX9744 and RESET;
	WX9809<=WX9746 and RESET;
	WX9811<=WX9748 and RESET;
	WX9813<=WX9750 and RESET;
	WX9815<=WX9752 and RESET;
	WX9817<=WX9754 and RESET;
	WX9819<=WX9756 and RESET;
	WX9821<=WX9758 and RESET;
	WX9823<=WX9760 and RESET;
	WX9825<=WX9762 and RESET;
	WX9827<=WX9764 and RESET;
	WX9829<=WX9766 and RESET;
	WX9831<=WX9768 and RESET;
	WX9833<=WX9770 and RESET;
	WX9835<=WX9772 and RESET;
	WX9837<=WX9774 and RESET;
	WX9839<=WX9776 and RESET;
	WX9841<=WX9778 and RESET;
	WX9843<=WX9780 and RESET;
	WX9845<=WX9782 and RESET;
	WX9847<=WX9784 and RESET;
	WX9849<=WX9786 and RESET;
	WX9851<=WX9788 and RESET;
	WX9853<=WX9790 and RESET;
	WX9855<=WX9792 and RESET;
	WX9857<=WX9794 and RESET;
	WX9859<=WX9796 and RESET;
	WX9861<=WX9798 and RESET;
	WX9863<=WX9800 and RESET;
	WX9865<=WX9802 and RESET;
	WX9867<=WX9804 and RESET;
	WX9869<=WX9806 and RESET;
	WX9871<=WX9808 and RESET;
	WX9873<=WX9810 and RESET;
	WX9875<=WX9812 and RESET;
	WX9877<=WX9814 and RESET;
	WX9879<=WX9816 and RESET;
	WX9881<=WX9818 and RESET;
	WX9883<=WX9820 and RESET;
	WX9885<=WX9822 and RESET;
	WX9887<=WX9824 and RESET;
	WX9889<=WX9826 and RESET;
	WX9891<=WX9828 and RESET;
	WX9893<=WX9830 and RESET;
	WX9895<=WX9832 and RESET;
	WX9897<=WX9834 and RESET;
	WX9899<=WX9836 and RESET;
	WX9901<=WX9838 and RESET;
	WX9903<=WX9840 and RESET;
	WX9905<=WX9842 and RESET;
	WX9907<=WX9844 and RESET;
	WX9909<=WX9846 and RESET;
	WX9911<=WX9848 and RESET;
	WX9913<=WX9850 and RESET;
	WX9915<=WX9852 and RESET;
	WX9917<=WX9854 and RESET;
	WX9919<=WX9856 and RESET;
	WX9921<=WX9858 and RESET;
	WX9923<=WX9860 and RESET;
	WX9925<=WX9862 and RESET;
	WX9927<=WX9864 and RESET;
	WX9929<=WX9866 and RESET;
	WX9931<=WX9868 and RESET;
	WX9933<=WX9870 and RESET;
	WX9935<=WX9872 and RESET;
	WX9937<=WX9874 and RESET;
	WX9939<=WX9876 and RESET;
	WX9941<=WX9878 and RESET;
	WX9943<=WX9880 and RESET;
	WX9945<=WX9882 and RESET;
	WX9947<=WX9884 and RESET;
	WX9949<=WX9886 and RESET;
	WX10058<=WX10057 and WX10056;
	WX10059<=WX9631 and WX10060;
	WX10065<=WX10064 and WX10056;
	WX10066<=WX9632 and WX10067;
	WX10072<=WX10071 and WX10056;
	WX10073<=WX9633 and WX10074;
	WX10079<=WX10078 and WX10056;
	WX10080<=WX9634 and WX10081;
	WX10086<=WX10085 and WX10056;
	WX10087<=WX9635 and WX10088;
	WX10093<=WX10092 and WX10056;
	WX10094<=WX9636 and WX10095;
	WX10100<=WX10099 and WX10056;
	WX10101<=WX9637 and WX10102;
	WX10107<=WX10106 and WX10056;
	WX10108<=WX9638 and WX10109;
	WX10114<=WX10113 and WX10056;
	WX10115<=WX9639 and WX10116;
	WX10121<=WX10120 and WX10056;
	WX10122<=WX9640 and WX10123;
	WX10128<=WX10127 and WX10056;
	WX10129<=WX9641 and WX10130;
	WX10135<=WX10134 and WX10056;
	WX10136<=WX9642 and WX10137;
	WX10142<=WX10141 and WX10056;
	WX10143<=WX9643 and WX10144;
	WX10149<=WX10148 and WX10056;
	WX10150<=WX9644 and WX10151;
	WX10156<=WX10155 and WX10056;
	WX10157<=WX9645 and WX10158;
	WX10163<=WX10162 and WX10056;
	WX10164<=WX9646 and WX10165;
	WX10170<=WX10169 and WX10056;
	WX10171<=WX9647 and WX10172;
	WX10177<=WX10176 and WX10056;
	WX10178<=WX9648 and WX10179;
	WX10184<=WX10183 and WX10056;
	WX10185<=WX9649 and WX10186;
	WX10191<=WX10190 and WX10056;
	WX10192<=WX9650 and WX10193;
	WX10198<=WX10197 and WX10056;
	WX10199<=WX9651 and WX10200;
	WX10205<=WX10204 and WX10056;
	WX10206<=WX9652 and WX10207;
	WX10212<=WX10211 and WX10056;
	WX10213<=WX9653 and WX10214;
	WX10219<=WX10218 and WX10056;
	WX10220<=WX9654 and WX10221;
	WX10226<=WX10225 and WX10056;
	WX10227<=WX9655 and WX10228;
	WX10233<=WX10232 and WX10056;
	WX10234<=WX9656 and WX10235;
	WX10240<=WX10239 and WX10056;
	WX10241<=WX9657 and WX10242;
	WX10247<=WX10246 and WX10056;
	WX10248<=WX9658 and WX10249;
	WX10254<=WX10253 and WX10056;
	WX10255<=WX9659 and WX10256;
	WX10261<=WX10260 and WX10056;
	WX10262<=WX9660 and WX10263;
	WX10268<=WX10267 and WX10056;
	WX10269<=WX9661 and WX10270;
	WX10275<=WX10274 and WX10056;
	WX10276<=WX9662 and WX10277;
	WX10315<=WX10285 and WX10314;
	WX10317<=WX10313 and WX10314;
	WX10319<=WX10312 and WX10314;
	WX10321<=WX10311 and WX10314;
	WX10323<=WX10284 and WX10314;
	WX10325<=WX10310 and WX10314;
	WX10327<=WX10309 and WX10314;
	WX10329<=WX10308 and WX10314;
	WX10331<=WX10307 and WX10314;
	WX10333<=WX10306 and WX10314;
	WX10335<=WX10305 and WX10314;
	WX10337<=WX10283 and WX10314;
	WX10339<=WX10304 and WX10314;
	WX10341<=WX10303 and WX10314;
	WX10343<=WX10302 and WX10314;
	WX10345<=WX10301 and WX10314;
	WX10347<=WX10282 and WX10314;
	WX10349<=WX10300 and WX10314;
	WX10351<=WX10299 and WX10314;
	WX10353<=WX10298 and WX10314;
	WX10355<=WX10297 and WX10314;
	WX10357<=WX10296 and WX10314;
	WX10359<=WX10295 and WX10314;
	WX10361<=WX10294 and WX10314;
	WX10363<=WX10293 and WX10314;
	WX10365<=WX10292 and WX10314;
	WX10367<=WX10291 and WX10314;
	WX10369<=WX10290 and WX10314;
	WX10371<=WX10289 and WX10314;
	WX10373<=WX10288 and WX10314;
	WX10375<=WX10287 and WX10314;
	WX10377<=WX10286 and WX10314;
	WX10379<=WX10390 and WX11347;
	WX10380<=WX10386 and WX10381;
	WX10383<=CRC_OUT_1_31 and WX11348;
	WX10384<=DATA_0_31 and WX10385;
	WX10387<=WX10829 and WX11348;
	WX10388<=WX11356 and WX10389;
	WX10393<=WX10404 and WX11347;
	WX10394<=WX10400 and WX10395;
	WX10397<=CRC_OUT_1_30 and WX11348;
	WX10398<=DATA_0_30 and WX10399;
	WX10401<=WX10831 and WX11348;
	WX10402<=WX11363 and WX10403;
	WX10407<=WX10418 and WX11347;
	WX10408<=WX10414 and WX10409;
	WX10411<=CRC_OUT_1_29 and WX11348;
	WX10412<=DATA_0_29 and WX10413;
	WX10415<=WX10833 and WX11348;
	WX10416<=WX11370 and WX10417;
	WX10421<=WX10432 and WX11347;
	WX10422<=WX10428 and WX10423;
	WX10425<=CRC_OUT_1_28 and WX11348;
	WX10426<=DATA_0_28 and WX10427;
	WX10429<=WX10835 and WX11348;
	WX10430<=WX11377 and WX10431;
	WX10435<=WX10446 and WX11347;
	WX10436<=WX10442 and WX10437;
	WX10439<=CRC_OUT_1_27 and WX11348;
	WX10440<=DATA_0_27 and WX10441;
	WX10443<=WX10837 and WX11348;
	WX10444<=WX11384 and WX10445;
	WX10449<=WX10460 and WX11347;
	WX10450<=WX10456 and WX10451;
	WX10453<=CRC_OUT_1_26 and WX11348;
	WX10454<=DATA_0_26 and WX10455;
	WX10457<=WX10839 and WX11348;
	WX10458<=WX11391 and WX10459;
	WX10463<=WX10474 and WX11347;
	WX10464<=WX10470 and WX10465;
	WX10467<=CRC_OUT_1_25 and WX11348;
	WX10468<=DATA_0_25 and WX10469;
	WX10471<=WX10841 and WX11348;
	WX10472<=WX11398 and WX10473;
	WX10477<=WX10488 and WX11347;
	WX10478<=WX10484 and WX10479;
	WX10481<=CRC_OUT_1_24 and WX11348;
	WX10482<=DATA_0_24 and WX10483;
	WX10485<=WX10843 and WX11348;
	WX10486<=WX11405 and WX10487;
	WX10491<=WX10502 and WX11347;
	WX10492<=WX10498 and WX10493;
	WX10495<=CRC_OUT_1_23 and WX11348;
	WX10496<=DATA_0_23 and WX10497;
	WX10499<=WX10845 and WX11348;
	WX10500<=WX11412 and WX10501;
	WX10505<=WX10516 and WX11347;
	WX10506<=WX10512 and WX10507;
	WX10509<=CRC_OUT_1_22 and WX11348;
	WX10510<=DATA_0_22 and WX10511;
	WX10513<=WX10847 and WX11348;
	WX10514<=WX11419 and WX10515;
	WX10519<=WX10530 and WX11347;
	WX10520<=WX10526 and WX10521;
	WX10523<=CRC_OUT_1_21 and WX11348;
	WX10524<=DATA_0_21 and WX10525;
	WX10527<=WX10849 and WX11348;
	WX10528<=WX11426 and WX10529;
	WX10533<=WX10544 and WX11347;
	WX10534<=WX10540 and WX10535;
	WX10537<=CRC_OUT_1_20 and WX11348;
	WX10538<=DATA_0_20 and WX10539;
	WX10541<=WX10851 and WX11348;
	WX10542<=WX11433 and WX10543;
	WX10547<=WX10558 and WX11347;
	WX10548<=WX10554 and WX10549;
	WX10551<=CRC_OUT_1_19 and WX11348;
	WX10552<=DATA_0_19 and WX10553;
	WX10555<=WX10853 and WX11348;
	WX10556<=WX11440 and WX10557;
	WX10561<=WX10572 and WX11347;
	WX10562<=WX10568 and WX10563;
	WX10565<=CRC_OUT_1_18 and WX11348;
	WX10566<=DATA_0_18 and WX10567;
	WX10569<=WX10855 and WX11348;
	WX10570<=WX11447 and WX10571;
	WX10575<=WX10586 and WX11347;
	WX10576<=WX10582 and WX10577;
	WX10579<=CRC_OUT_1_17 and WX11348;
	WX10580<=DATA_0_17 and WX10581;
	WX10583<=WX10857 and WX11348;
	WX10584<=WX11454 and WX10585;
	WX10589<=WX10600 and WX11347;
	WX10590<=WX10596 and WX10591;
	WX10593<=CRC_OUT_1_16 and WX11348;
	WX10594<=DATA_0_16 and WX10595;
	WX10597<=WX10859 and WX11348;
	WX10598<=WX11461 and WX10599;
	WX10603<=WX10614 and WX11347;
	WX10604<=WX10610 and WX10605;
	WX10607<=CRC_OUT_1_15 and WX11348;
	WX10608<=DATA_0_15 and WX10609;
	WX10611<=WX10861 and WX11348;
	WX10612<=WX11468 and WX10613;
	WX10617<=WX10628 and WX11347;
	WX10618<=WX10624 and WX10619;
	WX10621<=CRC_OUT_1_14 and WX11348;
	WX10622<=DATA_0_14 and WX10623;
	WX10625<=WX10863 and WX11348;
	WX10626<=WX11475 and WX10627;
	WX10631<=WX10642 and WX11347;
	WX10632<=WX10638 and WX10633;
	WX10635<=CRC_OUT_1_13 and WX11348;
	WX10636<=DATA_0_13 and WX10637;
	WX10639<=WX10865 and WX11348;
	WX10640<=WX11482 and WX10641;
	WX10645<=WX10656 and WX11347;
	WX10646<=WX10652 and WX10647;
	WX10649<=CRC_OUT_1_12 and WX11348;
	WX10650<=DATA_0_12 and WX10651;
	WX10653<=WX10867 and WX11348;
	WX10654<=WX11489 and WX10655;
	WX10659<=WX10670 and WX11347;
	WX10660<=WX10666 and WX10661;
	WX10663<=CRC_OUT_1_11 and WX11348;
	WX10664<=DATA_0_11 and WX10665;
	WX10667<=WX10869 and WX11348;
	WX10668<=WX11496 and WX10669;
	WX10673<=WX10684 and WX11347;
	WX10674<=WX10680 and WX10675;
	WX10677<=CRC_OUT_1_10 and WX11348;
	WX10678<=DATA_0_10 and WX10679;
	WX10681<=WX10871 and WX11348;
	WX10682<=WX11503 and WX10683;
	WX10687<=WX10698 and WX11347;
	WX10688<=WX10694 and WX10689;
	WX10691<=CRC_OUT_1_9 and WX11348;
	WX10692<=DATA_0_9 and WX10693;
	WX10695<=WX10873 and WX11348;
	WX10696<=WX11510 and WX10697;
	WX10701<=WX10712 and WX11347;
	WX10702<=WX10708 and WX10703;
	WX10705<=CRC_OUT_1_8 and WX11348;
	WX10706<=DATA_0_8 and WX10707;
	WX10709<=WX10875 and WX11348;
	WX10710<=WX11517 and WX10711;
	WX10715<=WX10726 and WX11347;
	WX10716<=WX10722 and WX10717;
	WX10719<=CRC_OUT_1_7 and WX11348;
	WX10720<=DATA_0_7 and WX10721;
	WX10723<=WX10877 and WX11348;
	WX10724<=WX11524 and WX10725;
	WX10729<=WX10740 and WX11347;
	WX10730<=WX10736 and WX10731;
	WX10733<=CRC_OUT_1_6 and WX11348;
	WX10734<=DATA_0_6 and WX10735;
	WX10737<=WX10879 and WX11348;
	WX10738<=WX11531 and WX10739;
	WX10743<=WX10754 and WX11347;
	WX10744<=WX10750 and WX10745;
	WX10747<=CRC_OUT_1_5 and WX11348;
	WX10748<=DATA_0_5 and WX10749;
	WX10751<=WX10881 and WX11348;
	WX10752<=WX11538 and WX10753;
	WX10757<=WX10768 and WX11347;
	WX10758<=WX10764 and WX10759;
	WX10761<=CRC_OUT_1_4 and WX11348;
	WX10762<=DATA_0_4 and WX10763;
	WX10765<=WX10883 and WX11348;
	WX10766<=WX11545 and WX10767;
	WX10771<=WX10782 and WX11347;
	WX10772<=WX10778 and WX10773;
	WX10775<=CRC_OUT_1_3 and WX11348;
	WX10776<=DATA_0_3 and WX10777;
	WX10779<=WX10885 and WX11348;
	WX10780<=WX11552 and WX10781;
	WX10785<=WX10796 and WX11347;
	WX10786<=WX10792 and WX10787;
	WX10789<=CRC_OUT_1_2 and WX11348;
	WX10790<=DATA_0_2 and WX10791;
	WX10793<=WX10887 and WX11348;
	WX10794<=WX11559 and WX10795;
	WX10799<=WX10810 and WX11347;
	WX10800<=WX10806 and WX10801;
	WX10803<=CRC_OUT_1_1 and WX11348;
	WX10804<=DATA_0_1 and WX10805;
	WX10807<=WX10889 and WX11348;
	WX10808<=WX11566 and WX10809;
	WX10813<=WX10824 and WX11347;
	WX10814<=WX10820 and WX10815;
	WX10817<=CRC_OUT_1_0 and WX11348;
	WX10818<=DATA_0_0 and WX10819;
	WX10821<=WX10891 and WX11348;
	WX10822<=WX11573 and WX10823;
	WX10828<=WX10831 and RESET;
	WX10830<=WX10833 and RESET;
	WX10832<=WX10835 and RESET;
	WX10834<=WX10837 and RESET;
	WX10836<=WX10839 and RESET;
	WX10838<=WX10841 and RESET;
	WX10840<=WX10843 and RESET;
	WX10842<=WX10845 and RESET;
	WX10844<=WX10847 and RESET;
	WX10846<=WX10849 and RESET;
	WX10848<=WX10851 and RESET;
	WX10850<=WX10853 and RESET;
	WX10852<=WX10855 and RESET;
	WX10854<=WX10857 and RESET;
	WX10856<=WX10859 and RESET;
	WX10858<=WX10861 and RESET;
	WX10860<=WX10863 and RESET;
	WX10862<=WX10865 and RESET;
	WX10864<=WX10867 and RESET;
	WX10866<=WX10869 and RESET;
	WX10868<=WX10871 and RESET;
	WX10870<=WX10873 and RESET;
	WX10872<=WX10875 and RESET;
	WX10874<=WX10877 and RESET;
	WX10876<=WX10879 and RESET;
	WX10878<=WX10881 and RESET;
	WX10880<=WX10883 and RESET;
	WX10882<=WX10885 and RESET;
	WX10884<=WX10887 and RESET;
	WX10886<=WX10889 and RESET;
	WX10888<=WX10891 and RESET;
	WX10890<=WX10827 and RESET;
	WX10988<=WX10392 and RESET;
	WX10990<=WX10406 and RESET;
	WX10992<=WX10420 and RESET;
	WX10994<=WX10434 and RESET;
	WX10996<=WX10448 and RESET;
	WX10998<=WX10462 and RESET;
	WX11000<=WX10476 and RESET;
	WX11002<=WX10490 and RESET;
	WX11004<=WX10504 and RESET;
	WX11006<=WX10518 and RESET;
	WX11008<=WX10532 and RESET;
	WX11010<=WX10546 and RESET;
	WX11012<=WX10560 and RESET;
	WX11014<=WX10574 and RESET;
	WX11016<=WX10588 and RESET;
	WX11018<=WX10602 and RESET;
	WX11020<=WX10616 and RESET;
	WX11022<=WX10630 and RESET;
	WX11024<=WX10644 and RESET;
	WX11026<=WX10658 and RESET;
	WX11028<=WX10672 and RESET;
	WX11030<=WX10686 and RESET;
	WX11032<=WX10700 and RESET;
	WX11034<=WX10714 and RESET;
	WX11036<=WX10728 and RESET;
	WX11038<=WX10742 and RESET;
	WX11040<=WX10756 and RESET;
	WX11042<=WX10770 and RESET;
	WX11044<=WX10784 and RESET;
	WX11046<=WX10798 and RESET;
	WX11048<=WX10812 and RESET;
	WX11050<=WX10826 and RESET;
	WX11052<=WX10989 and RESET;
	WX11054<=WX10991 and RESET;
	WX11056<=WX10993 and RESET;
	WX11058<=WX10995 and RESET;
	WX11060<=WX10997 and RESET;
	WX11062<=WX10999 and RESET;
	WX11064<=WX11001 and RESET;
	WX11066<=WX11003 and RESET;
	WX11068<=WX11005 and RESET;
	WX11070<=WX11007 and RESET;
	WX11072<=WX11009 and RESET;
	WX11074<=WX11011 and RESET;
	WX11076<=WX11013 and RESET;
	WX11078<=WX11015 and RESET;
	WX11080<=WX11017 and RESET;
	WX11082<=WX11019 and RESET;
	WX11084<=WX11021 and RESET;
	WX11086<=WX11023 and RESET;
	WX11088<=WX11025 and RESET;
	WX11090<=WX11027 and RESET;
	WX11092<=WX11029 and RESET;
	WX11094<=WX11031 and RESET;
	WX11096<=WX11033 and RESET;
	WX11098<=WX11035 and RESET;
	WX11100<=WX11037 and RESET;
	WX11102<=WX11039 and RESET;
	WX11104<=WX11041 and RESET;
	WX11106<=WX11043 and RESET;
	WX11108<=WX11045 and RESET;
	WX11110<=WX11047 and RESET;
	WX11112<=WX11049 and RESET;
	WX11114<=WX11051 and RESET;
	WX11116<=WX11053 and RESET;
	WX11118<=WX11055 and RESET;
	WX11120<=WX11057 and RESET;
	WX11122<=WX11059 and RESET;
	WX11124<=WX11061 and RESET;
	WX11126<=WX11063 and RESET;
	WX11128<=WX11065 and RESET;
	WX11130<=WX11067 and RESET;
	WX11132<=WX11069 and RESET;
	WX11134<=WX11071 and RESET;
	WX11136<=WX11073 and RESET;
	WX11138<=WX11075 and RESET;
	WX11140<=WX11077 and RESET;
	WX11142<=WX11079 and RESET;
	WX11144<=WX11081 and RESET;
	WX11146<=WX11083 and RESET;
	WX11148<=WX11085 and RESET;
	WX11150<=WX11087 and RESET;
	WX11152<=WX11089 and RESET;
	WX11154<=WX11091 and RESET;
	WX11156<=WX11093 and RESET;
	WX11158<=WX11095 and RESET;
	WX11160<=WX11097 and RESET;
	WX11162<=WX11099 and RESET;
	WX11164<=WX11101 and RESET;
	WX11166<=WX11103 and RESET;
	WX11168<=WX11105 and RESET;
	WX11170<=WX11107 and RESET;
	WX11172<=WX11109 and RESET;
	WX11174<=WX11111 and RESET;
	WX11176<=WX11113 and RESET;
	WX11178<=WX11115 and RESET;
	WX11180<=WX11117 and RESET;
	WX11182<=WX11119 and RESET;
	WX11184<=WX11121 and RESET;
	WX11186<=WX11123 and RESET;
	WX11188<=WX11125 and RESET;
	WX11190<=WX11127 and RESET;
	WX11192<=WX11129 and RESET;
	WX11194<=WX11131 and RESET;
	WX11196<=WX11133 and RESET;
	WX11198<=WX11135 and RESET;
	WX11200<=WX11137 and RESET;
	WX11202<=WX11139 and RESET;
	WX11204<=WX11141 and RESET;
	WX11206<=WX11143 and RESET;
	WX11208<=WX11145 and RESET;
	WX11210<=WX11147 and RESET;
	WX11212<=WX11149 and RESET;
	WX11214<=WX11151 and RESET;
	WX11216<=WX11153 and RESET;
	WX11218<=WX11155 and RESET;
	WX11220<=WX11157 and RESET;
	WX11222<=WX11159 and RESET;
	WX11224<=WX11161 and RESET;
	WX11226<=WX11163 and RESET;
	WX11228<=WX11165 and RESET;
	WX11230<=WX11167 and RESET;
	WX11232<=WX11169 and RESET;
	WX11234<=WX11171 and RESET;
	WX11236<=WX11173 and RESET;
	WX11238<=WX11175 and RESET;
	WX11240<=WX11177 and RESET;
	WX11242<=WX11179 and RESET;
	WX11351<=WX11350 and WX11349;
	WX11352<=WX10924 and WX11353;
	WX11358<=WX11357 and WX11349;
	WX11359<=WX10925 and WX11360;
	WX11365<=WX11364 and WX11349;
	WX11366<=WX10926 and WX11367;
	WX11372<=WX11371 and WX11349;
	WX11373<=WX10927 and WX11374;
	WX11379<=WX11378 and WX11349;
	WX11380<=WX10928 and WX11381;
	WX11386<=WX11385 and WX11349;
	WX11387<=WX10929 and WX11388;
	WX11393<=WX11392 and WX11349;
	WX11394<=WX10930 and WX11395;
	WX11400<=WX11399 and WX11349;
	WX11401<=WX10931 and WX11402;
	WX11407<=WX11406 and WX11349;
	WX11408<=WX10932 and WX11409;
	WX11414<=WX11413 and WX11349;
	WX11415<=WX10933 and WX11416;
	WX11421<=WX11420 and WX11349;
	WX11422<=WX10934 and WX11423;
	WX11428<=WX11427 and WX11349;
	WX11429<=WX10935 and WX11430;
	WX11435<=WX11434 and WX11349;
	WX11436<=WX10936 and WX11437;
	WX11442<=WX11441 and WX11349;
	WX11443<=WX10937 and WX11444;
	WX11449<=WX11448 and WX11349;
	WX11450<=WX10938 and WX11451;
	WX11456<=WX11455 and WX11349;
	WX11457<=WX10939 and WX11458;
	WX11463<=WX11462 and WX11349;
	WX11464<=WX10940 and WX11465;
	WX11470<=WX11469 and WX11349;
	WX11471<=WX10941 and WX11472;
	WX11477<=WX11476 and WX11349;
	WX11478<=WX10942 and WX11479;
	WX11484<=WX11483 and WX11349;
	WX11485<=WX10943 and WX11486;
	WX11491<=WX11490 and WX11349;
	WX11492<=WX10944 and WX11493;
	WX11498<=WX11497 and WX11349;
	WX11499<=WX10945 and WX11500;
	WX11505<=WX11504 and WX11349;
	WX11506<=WX10946 and WX11507;
	WX11512<=WX11511 and WX11349;
	WX11513<=WX10947 and WX11514;
	WX11519<=WX11518 and WX11349;
	WX11520<=WX10948 and WX11521;
	WX11526<=WX11525 and WX11349;
	WX11527<=WX10949 and WX11528;
	WX11533<=WX11532 and WX11349;
	WX11534<=WX10950 and WX11535;
	WX11540<=WX11539 and WX11349;
	WX11541<=WX10951 and WX11542;
	WX11547<=WX11546 and WX11349;
	WX11548<=WX10952 and WX11549;
	WX11554<=WX11553 and WX11349;
	WX11555<=WX10953 and WX11556;
	WX11561<=WX11560 and WX11349;
	WX11562<=WX10954 and WX11563;
	WX11568<=WX11567 and WX11349;
	WX11569<=WX10955 and WX11570;
	WX11608<=WX11578 and WX11607;
	WX11610<=WX11606 and WX11607;
	WX11612<=WX11605 and WX11607;
	WX11614<=WX11604 and WX11607;
	WX11616<=WX11577 and WX11607;
	WX11618<=WX11603 and WX11607;
	WX11620<=WX11602 and WX11607;
	WX11622<=WX11601 and WX11607;
	WX11624<=WX11600 and WX11607;
	WX11626<=WX11599 and WX11607;
	WX11628<=WX11598 and WX11607;
	WX11630<=WX11576 and WX11607;
	WX11632<=WX11597 and WX11607;
	WX11634<=WX11596 and WX11607;
	WX11636<=WX11595 and WX11607;
	WX11638<=WX11594 and WX11607;
	WX11640<=WX11575 and WX11607;
	WX11642<=WX11593 and WX11607;
	WX11644<=WX11592 and WX11607;
	WX11646<=WX11591 and WX11607;
	WX11648<=WX11590 and WX11607;
	WX11650<=WX11589 and WX11607;
	WX11652<=WX11588 and WX11607;
	WX11654<=WX11587 and WX11607;
	WX11656<=WX11586 and WX11607;
	WX11658<=WX11585 and WX11607;
	WX11660<=WX11584 and WX11607;
	WX11662<=WX11583 and WX11607;
	WX11664<=WX11582 and WX11607;
	WX11666<=WX11581 and WX11607;
	WX11668<=WX11580 and WX11607;
	WX11670<=WX11579 and WX11607;
	I1986<= not (I1996 and I1997);
	I1987<= not (I1989 and I1990);
	I1988<= not (WX1001 and WX645);
	I1989<= not (WX1001 and I1988);
	I1990<= not (WX645 and I1988);
	I1995<= not (WX709 and I1987);
	I1996<= not (WX709 and I1995);
	I1997<= not (I1987 and I1995);
	I2002<= not (I2004 and I2005);
	I2003<= not (WX773 and WX837);
	I2004<= not (WX773 and I2003);
	I2005<= not (WX837 and I2003);
	I2010<= not (I1986 and I2002);
	I2011<= not (I1986 and I2010);
	I2012<= not (I2002 and I2010);
	I2017<= not (I2027 and I2028);
	I2018<= not (I2020 and I2021);
	I2019<= not (WX1001 and WX647);
	I2020<= not (WX1001 and I2019);
	I2021<= not (WX647 and I2019);
	I2026<= not (WX711 and I2018);
	I2027<= not (WX711 and I2026);
	I2028<= not (I2018 and I2026);
	I2033<= not (I2035 and I2036);
	I2034<= not (WX775 and WX839);
	I2035<= not (WX775 and I2034);
	I2036<= not (WX839 and I2034);
	I2041<= not (I2017 and I2033);
	I2042<= not (I2017 and I2041);
	I2043<= not (I2033 and I2041);
	I2048<= not (I2058 and I2059);
	I2049<= not (I2051 and I2052);
	I2050<= not (WX1001 and WX649);
	I2051<= not (WX1001 and I2050);
	I2052<= not (WX649 and I2050);
	I2057<= not (WX713 and I2049);
	I2058<= not (WX713 and I2057);
	I2059<= not (I2049 and I2057);
	I2064<= not (I2066 and I2067);
	I2065<= not (WX777 and WX841);
	I2066<= not (WX777 and I2065);
	I2067<= not (WX841 and I2065);
	I2072<= not (I2048 and I2064);
	I2073<= not (I2048 and I2072);
	I2074<= not (I2064 and I2072);
	I2079<= not (I2089 and I2090);
	I2080<= not (I2082 and I2083);
	I2081<= not (WX1001 and WX651);
	I2082<= not (WX1001 and I2081);
	I2083<= not (WX651 and I2081);
	I2088<= not (WX715 and I2080);
	I2089<= not (WX715 and I2088);
	I2090<= not (I2080 and I2088);
	I2095<= not (I2097 and I2098);
	I2096<= not (WX779 and WX843);
	I2097<= not (WX779 and I2096);
	I2098<= not (WX843 and I2096);
	I2103<= not (I2079 and I2095);
	I2104<= not (I2079 and I2103);
	I2105<= not (I2095 and I2103);
	I2110<= not (I2120 and I2121);
	I2111<= not (I2113 and I2114);
	I2112<= not (WX1001 and WX653);
	I2113<= not (WX1001 and I2112);
	I2114<= not (WX653 and I2112);
	I2119<= not (WX717 and I2111);
	I2120<= not (WX717 and I2119);
	I2121<= not (I2111 and I2119);
	I2126<= not (I2128 and I2129);
	I2127<= not (WX781 and WX845);
	I2128<= not (WX781 and I2127);
	I2129<= not (WX845 and I2127);
	I2134<= not (I2110 and I2126);
	I2135<= not (I2110 and I2134);
	I2136<= not (I2126 and I2134);
	I2141<= not (I2151 and I2152);
	I2142<= not (I2144 and I2145);
	I2143<= not (WX1001 and WX655);
	I2144<= not (WX1001 and I2143);
	I2145<= not (WX655 and I2143);
	I2150<= not (WX719 and I2142);
	I2151<= not (WX719 and I2150);
	I2152<= not (I2142 and I2150);
	I2157<= not (I2159 and I2160);
	I2158<= not (WX783 and WX847);
	I2159<= not (WX783 and I2158);
	I2160<= not (WX847 and I2158);
	I2165<= not (I2141 and I2157);
	I2166<= not (I2141 and I2165);
	I2167<= not (I2157 and I2165);
	I2172<= not (I2182 and I2183);
	I2173<= not (I2175 and I2176);
	I2174<= not (WX1001 and WX657);
	I2175<= not (WX1001 and I2174);
	I2176<= not (WX657 and I2174);
	I2181<= not (WX721 and I2173);
	I2182<= not (WX721 and I2181);
	I2183<= not (I2173 and I2181);
	I2188<= not (I2190 and I2191);
	I2189<= not (WX785 and WX849);
	I2190<= not (WX785 and I2189);
	I2191<= not (WX849 and I2189);
	I2196<= not (I2172 and I2188);
	I2197<= not (I2172 and I2196);
	I2198<= not (I2188 and I2196);
	I2203<= not (I2213 and I2214);
	I2204<= not (I2206 and I2207);
	I2205<= not (WX1001 and WX659);
	I2206<= not (WX1001 and I2205);
	I2207<= not (WX659 and I2205);
	I2212<= not (WX723 and I2204);
	I2213<= not (WX723 and I2212);
	I2214<= not (I2204 and I2212);
	I2219<= not (I2221 and I2222);
	I2220<= not (WX787 and WX851);
	I2221<= not (WX787 and I2220);
	I2222<= not (WX851 and I2220);
	I2227<= not (I2203 and I2219);
	I2228<= not (I2203 and I2227);
	I2229<= not (I2219 and I2227);
	I2234<= not (I2244 and I2245);
	I2235<= not (I2237 and I2238);
	I2236<= not (WX1001 and WX661);
	I2237<= not (WX1001 and I2236);
	I2238<= not (WX661 and I2236);
	I2243<= not (WX725 and I2235);
	I2244<= not (WX725 and I2243);
	I2245<= not (I2235 and I2243);
	I2250<= not (I2252 and I2253);
	I2251<= not (WX789 and WX853);
	I2252<= not (WX789 and I2251);
	I2253<= not (WX853 and I2251);
	I2258<= not (I2234 and I2250);
	I2259<= not (I2234 and I2258);
	I2260<= not (I2250 and I2258);
	I2265<= not (I2275 and I2276);
	I2266<= not (I2268 and I2269);
	I2267<= not (WX1001 and WX663);
	I2268<= not (WX1001 and I2267);
	I2269<= not (WX663 and I2267);
	I2274<= not (WX727 and I2266);
	I2275<= not (WX727 and I2274);
	I2276<= not (I2266 and I2274);
	I2281<= not (I2283 and I2284);
	I2282<= not (WX791 and WX855);
	I2283<= not (WX791 and I2282);
	I2284<= not (WX855 and I2282);
	I2289<= not (I2265 and I2281);
	I2290<= not (I2265 and I2289);
	I2291<= not (I2281 and I2289);
	I2296<= not (I2306 and I2307);
	I2297<= not (I2299 and I2300);
	I2298<= not (WX1001 and WX665);
	I2299<= not (WX1001 and I2298);
	I2300<= not (WX665 and I2298);
	I2305<= not (WX729 and I2297);
	I2306<= not (WX729 and I2305);
	I2307<= not (I2297 and I2305);
	I2312<= not (I2314 and I2315);
	I2313<= not (WX793 and WX857);
	I2314<= not (WX793 and I2313);
	I2315<= not (WX857 and I2313);
	I2320<= not (I2296 and I2312);
	I2321<= not (I2296 and I2320);
	I2322<= not (I2312 and I2320);
	I2327<= not (I2337 and I2338);
	I2328<= not (I2330 and I2331);
	I2329<= not (WX1001 and WX667);
	I2330<= not (WX1001 and I2329);
	I2331<= not (WX667 and I2329);
	I2336<= not (WX731 and I2328);
	I2337<= not (WX731 and I2336);
	I2338<= not (I2328 and I2336);
	I2343<= not (I2345 and I2346);
	I2344<= not (WX795 and WX859);
	I2345<= not (WX795 and I2344);
	I2346<= not (WX859 and I2344);
	I2351<= not (I2327 and I2343);
	I2352<= not (I2327 and I2351);
	I2353<= not (I2343 and I2351);
	I2358<= not (I2368 and I2369);
	I2359<= not (I2361 and I2362);
	I2360<= not (WX1001 and WX669);
	I2361<= not (WX1001 and I2360);
	I2362<= not (WX669 and I2360);
	I2367<= not (WX733 and I2359);
	I2368<= not (WX733 and I2367);
	I2369<= not (I2359 and I2367);
	I2374<= not (I2376 and I2377);
	I2375<= not (WX797 and WX861);
	I2376<= not (WX797 and I2375);
	I2377<= not (WX861 and I2375);
	I2382<= not (I2358 and I2374);
	I2383<= not (I2358 and I2382);
	I2384<= not (I2374 and I2382);
	I2389<= not (I2399 and I2400);
	I2390<= not (I2392 and I2393);
	I2391<= not (WX1001 and WX671);
	I2392<= not (WX1001 and I2391);
	I2393<= not (WX671 and I2391);
	I2398<= not (WX735 and I2390);
	I2399<= not (WX735 and I2398);
	I2400<= not (I2390 and I2398);
	I2405<= not (I2407 and I2408);
	I2406<= not (WX799 and WX863);
	I2407<= not (WX799 and I2406);
	I2408<= not (WX863 and I2406);
	I2413<= not (I2389 and I2405);
	I2414<= not (I2389 and I2413);
	I2415<= not (I2405 and I2413);
	I2420<= not (I2430 and I2431);
	I2421<= not (I2423 and I2424);
	I2422<= not (WX1001 and WX673);
	I2423<= not (WX1001 and I2422);
	I2424<= not (WX673 and I2422);
	I2429<= not (WX737 and I2421);
	I2430<= not (WX737 and I2429);
	I2431<= not (I2421 and I2429);
	I2436<= not (I2438 and I2439);
	I2437<= not (WX801 and WX865);
	I2438<= not (WX801 and I2437);
	I2439<= not (WX865 and I2437);
	I2444<= not (I2420 and I2436);
	I2445<= not (I2420 and I2444);
	I2446<= not (I2436 and I2444);
	I2451<= not (I2461 and I2462);
	I2452<= not (I2454 and I2455);
	I2453<= not (WX1001 and WX675);
	I2454<= not (WX1001 and I2453);
	I2455<= not (WX675 and I2453);
	I2460<= not (WX739 and I2452);
	I2461<= not (WX739 and I2460);
	I2462<= not (I2452 and I2460);
	I2467<= not (I2469 and I2470);
	I2468<= not (WX803 and WX867);
	I2469<= not (WX803 and I2468);
	I2470<= not (WX867 and I2468);
	I2475<= not (I2451 and I2467);
	I2476<= not (I2451 and I2475);
	I2477<= not (I2467 and I2475);
	I2482<= not (I2492 and I2493);
	I2483<= not (I2485 and I2486);
	I2484<= not (WX1002 and WX677);
	I2485<= not (WX1002 and I2484);
	I2486<= not (WX677 and I2484);
	I2491<= not (WX741 and I2483);
	I2492<= not (WX741 and I2491);
	I2493<= not (I2483 and I2491);
	I2498<= not (I2500 and I2501);
	I2499<= not (WX805 and WX869);
	I2500<= not (WX805 and I2499);
	I2501<= not (WX869 and I2499);
	I2506<= not (I2482 and I2498);
	I2507<= not (I2482 and I2506);
	I2508<= not (I2498 and I2506);
	I2513<= not (I2523 and I2524);
	I2514<= not (I2516 and I2517);
	I2515<= not (WX1002 and WX679);
	I2516<= not (WX1002 and I2515);
	I2517<= not (WX679 and I2515);
	I2522<= not (WX743 and I2514);
	I2523<= not (WX743 and I2522);
	I2524<= not (I2514 and I2522);
	I2529<= not (I2531 and I2532);
	I2530<= not (WX807 and WX871);
	I2531<= not (WX807 and I2530);
	I2532<= not (WX871 and I2530);
	I2537<= not (I2513 and I2529);
	I2538<= not (I2513 and I2537);
	I2539<= not (I2529 and I2537);
	I2544<= not (I2554 and I2555);
	I2545<= not (I2547 and I2548);
	I2546<= not (WX1002 and WX681);
	I2547<= not (WX1002 and I2546);
	I2548<= not (WX681 and I2546);
	I2553<= not (WX745 and I2545);
	I2554<= not (WX745 and I2553);
	I2555<= not (I2545 and I2553);
	I2560<= not (I2562 and I2563);
	I2561<= not (WX809 and WX873);
	I2562<= not (WX809 and I2561);
	I2563<= not (WX873 and I2561);
	I2568<= not (I2544 and I2560);
	I2569<= not (I2544 and I2568);
	I2570<= not (I2560 and I2568);
	I2575<= not (I2585 and I2586);
	I2576<= not (I2578 and I2579);
	I2577<= not (WX1002 and WX683);
	I2578<= not (WX1002 and I2577);
	I2579<= not (WX683 and I2577);
	I2584<= not (WX747 and I2576);
	I2585<= not (WX747 and I2584);
	I2586<= not (I2576 and I2584);
	I2591<= not (I2593 and I2594);
	I2592<= not (WX811 and WX875);
	I2593<= not (WX811 and I2592);
	I2594<= not (WX875 and I2592);
	I2599<= not (I2575 and I2591);
	I2600<= not (I2575 and I2599);
	I2601<= not (I2591 and I2599);
	I2606<= not (I2616 and I2617);
	I2607<= not (I2609 and I2610);
	I2608<= not (WX1002 and WX685);
	I2609<= not (WX1002 and I2608);
	I2610<= not (WX685 and I2608);
	I2615<= not (WX749 and I2607);
	I2616<= not (WX749 and I2615);
	I2617<= not (I2607 and I2615);
	I2622<= not (I2624 and I2625);
	I2623<= not (WX813 and WX877);
	I2624<= not (WX813 and I2623);
	I2625<= not (WX877 and I2623);
	I2630<= not (I2606 and I2622);
	I2631<= not (I2606 and I2630);
	I2632<= not (I2622 and I2630);
	I2637<= not (I2647 and I2648);
	I2638<= not (I2640 and I2641);
	I2639<= not (WX1002 and WX687);
	I2640<= not (WX1002 and I2639);
	I2641<= not (WX687 and I2639);
	I2646<= not (WX751 and I2638);
	I2647<= not (WX751 and I2646);
	I2648<= not (I2638 and I2646);
	I2653<= not (I2655 and I2656);
	I2654<= not (WX815 and WX879);
	I2655<= not (WX815 and I2654);
	I2656<= not (WX879 and I2654);
	I2661<= not (I2637 and I2653);
	I2662<= not (I2637 and I2661);
	I2663<= not (I2653 and I2661);
	I2668<= not (I2678 and I2679);
	I2669<= not (I2671 and I2672);
	I2670<= not (WX1002 and WX689);
	I2671<= not (WX1002 and I2670);
	I2672<= not (WX689 and I2670);
	I2677<= not (WX753 and I2669);
	I2678<= not (WX753 and I2677);
	I2679<= not (I2669 and I2677);
	I2684<= not (I2686 and I2687);
	I2685<= not (WX817 and WX881);
	I2686<= not (WX817 and I2685);
	I2687<= not (WX881 and I2685);
	I2692<= not (I2668 and I2684);
	I2693<= not (I2668 and I2692);
	I2694<= not (I2684 and I2692);
	I2699<= not (I2709 and I2710);
	I2700<= not (I2702 and I2703);
	I2701<= not (WX1002 and WX691);
	I2702<= not (WX1002 and I2701);
	I2703<= not (WX691 and I2701);
	I2708<= not (WX755 and I2700);
	I2709<= not (WX755 and I2708);
	I2710<= not (I2700 and I2708);
	I2715<= not (I2717 and I2718);
	I2716<= not (WX819 and WX883);
	I2717<= not (WX819 and I2716);
	I2718<= not (WX883 and I2716);
	I2723<= not (I2699 and I2715);
	I2724<= not (I2699 and I2723);
	I2725<= not (I2715 and I2723);
	I2730<= not (I2740 and I2741);
	I2731<= not (I2733 and I2734);
	I2732<= not (WX1002 and WX693);
	I2733<= not (WX1002 and I2732);
	I2734<= not (WX693 and I2732);
	I2739<= not (WX757 and I2731);
	I2740<= not (WX757 and I2739);
	I2741<= not (I2731 and I2739);
	I2746<= not (I2748 and I2749);
	I2747<= not (WX821 and WX885);
	I2748<= not (WX821 and I2747);
	I2749<= not (WX885 and I2747);
	I2754<= not (I2730 and I2746);
	I2755<= not (I2730 and I2754);
	I2756<= not (I2746 and I2754);
	I2761<= not (I2771 and I2772);
	I2762<= not (I2764 and I2765);
	I2763<= not (WX1002 and WX695);
	I2764<= not (WX1002 and I2763);
	I2765<= not (WX695 and I2763);
	I2770<= not (WX759 and I2762);
	I2771<= not (WX759 and I2770);
	I2772<= not (I2762 and I2770);
	I2777<= not (I2779 and I2780);
	I2778<= not (WX823 and WX887);
	I2779<= not (WX823 and I2778);
	I2780<= not (WX887 and I2778);
	I2785<= not (I2761 and I2777);
	I2786<= not (I2761 and I2785);
	I2787<= not (I2777 and I2785);
	I2792<= not (I2802 and I2803);
	I2793<= not (I2795 and I2796);
	I2794<= not (WX1002 and WX697);
	I2795<= not (WX1002 and I2794);
	I2796<= not (WX697 and I2794);
	I2801<= not (WX761 and I2793);
	I2802<= not (WX761 and I2801);
	I2803<= not (I2793 and I2801);
	I2808<= not (I2810 and I2811);
	I2809<= not (WX825 and WX889);
	I2810<= not (WX825 and I2809);
	I2811<= not (WX889 and I2809);
	I2816<= not (I2792 and I2808);
	I2817<= not (I2792 and I2816);
	I2818<= not (I2808 and I2816);
	I2823<= not (I2833 and I2834);
	I2824<= not (I2826 and I2827);
	I2825<= not (WX1002 and WX699);
	I2826<= not (WX1002 and I2825);
	I2827<= not (WX699 and I2825);
	I2832<= not (WX763 and I2824);
	I2833<= not (WX763 and I2832);
	I2834<= not (I2824 and I2832);
	I2839<= not (I2841 and I2842);
	I2840<= not (WX827 and WX891);
	I2841<= not (WX827 and I2840);
	I2842<= not (WX891 and I2840);
	I2847<= not (I2823 and I2839);
	I2848<= not (I2823 and I2847);
	I2849<= not (I2839 and I2847);
	I2854<= not (I2864 and I2865);
	I2855<= not (I2857 and I2858);
	I2856<= not (WX1002 and WX701);
	I2857<= not (WX1002 and I2856);
	I2858<= not (WX701 and I2856);
	I2863<= not (WX765 and I2855);
	I2864<= not (WX765 and I2863);
	I2865<= not (I2855 and I2863);
	I2870<= not (I2872 and I2873);
	I2871<= not (WX829 and WX893);
	I2872<= not (WX829 and I2871);
	I2873<= not (WX893 and I2871);
	I2878<= not (I2854 and I2870);
	I2879<= not (I2854 and I2878);
	I2880<= not (I2870 and I2878);
	I2885<= not (I2895 and I2896);
	I2886<= not (I2888 and I2889);
	I2887<= not (WX1002 and WX703);
	I2888<= not (WX1002 and I2887);
	I2889<= not (WX703 and I2887);
	I2894<= not (WX767 and I2886);
	I2895<= not (WX767 and I2894);
	I2896<= not (I2886 and I2894);
	I2901<= not (I2903 and I2904);
	I2902<= not (WX831 and WX895);
	I2903<= not (WX831 and I2902);
	I2904<= not (WX895 and I2902);
	I2909<= not (I2885 and I2901);
	I2910<= not (I2885 and I2909);
	I2911<= not (I2901 and I2909);
	I2916<= not (I2926 and I2927);
	I2917<= not (I2919 and I2920);
	I2918<= not (WX1002 and WX705);
	I2919<= not (WX1002 and I2918);
	I2920<= not (WX705 and I2918);
	I2925<= not (WX769 and I2917);
	I2926<= not (WX769 and I2925);
	I2927<= not (I2917 and I2925);
	I2932<= not (I2934 and I2935);
	I2933<= not (WX833 and WX897);
	I2934<= not (WX833 and I2933);
	I2935<= not (WX897 and I2933);
	I2940<= not (I2916 and I2932);
	I2941<= not (I2916 and I2940);
	I2942<= not (I2932 and I2940);
	I2947<= not (I2957 and I2958);
	I2948<= not (I2950 and I2951);
	I2949<= not (WX1002 and WX707);
	I2950<= not (WX1002 and I2949);
	I2951<= not (WX707 and I2949);
	I2956<= not (WX771 and I2948);
	I2957<= not (WX771 and I2956);
	I2958<= not (I2948 and I2956);
	I2963<= not (I2965 and I2966);
	I2964<= not (WX835 and WX899);
	I2965<= not (WX835 and I2964);
	I2966<= not (WX899 and I2964);
	I2971<= not (I2947 and I2963);
	I2972<= not (I2947 and I2971);
	I2973<= not (I2963 and I2971);
	I3052<= not (WX580 and WX485);
	I3053<= not (WX580 and I3052);
	I3054<= not (WX485 and I3052);
	I3065<= not (WX581 and WX487);
	I3066<= not (WX581 and I3065);
	I3067<= not (WX487 and I3065);
	I3078<= not (WX582 and WX489);
	I3079<= not (WX582 and I3078);
	I3080<= not (WX489 and I3078);
	I3091<= not (WX583 and WX491);
	I3092<= not (WX583 and I3091);
	I3093<= not (WX491 and I3091);
	I3104<= not (WX584 and WX493);
	I3105<= not (WX584 and I3104);
	I3106<= not (WX493 and I3104);
	I3117<= not (WX585 and WX495);
	I3118<= not (WX585 and I3117);
	I3119<= not (WX495 and I3117);
	I3130<= not (WX586 and WX497);
	I3131<= not (WX586 and I3130);
	I3132<= not (WX497 and I3130);
	I3143<= not (WX587 and WX499);
	I3144<= not (WX587 and I3143);
	I3145<= not (WX499 and I3143);
	I3156<= not (WX588 and WX501);
	I3157<= not (WX588 and I3156);
	I3158<= not (WX501 and I3156);
	I3169<= not (WX589 and WX503);
	I3170<= not (WX589 and I3169);
	I3171<= not (WX503 and I3169);
	I3182<= not (WX590 and WX505);
	I3183<= not (WX590 and I3182);
	I3184<= not (WX505 and I3182);
	I3195<= not (WX591 and WX507);
	I3196<= not (WX591 and I3195);
	I3197<= not (WX507 and I3195);
	I3208<= not (WX592 and WX509);
	I3209<= not (WX592 and I3208);
	I3210<= not (WX509 and I3208);
	I3221<= not (WX593 and WX511);
	I3222<= not (WX593 and I3221);
	I3223<= not (WX511 and I3221);
	I3234<= not (WX594 and WX513);
	I3235<= not (WX594 and I3234);
	I3236<= not (WX513 and I3234);
	I3247<= not (WX595 and WX515);
	I3248<= not (WX595 and I3247);
	I3249<= not (WX515 and I3247);
	I3260<= not (WX596 and WX517);
	I3261<= not (WX596 and I3260);
	I3262<= not (WX517 and I3260);
	I3273<= not (WX597 and WX519);
	I3274<= not (WX597 and I3273);
	I3275<= not (WX519 and I3273);
	I3286<= not (WX598 and WX521);
	I3287<= not (WX598 and I3286);
	I3288<= not (WX521 and I3286);
	I3299<= not (WX599 and WX523);
	I3300<= not (WX599 and I3299);
	I3301<= not (WX523 and I3299);
	I3312<= not (WX600 and WX525);
	I3313<= not (WX600 and I3312);
	I3314<= not (WX525 and I3312);
	I3325<= not (WX601 and WX527);
	I3326<= not (WX601 and I3325);
	I3327<= not (WX527 and I3325);
	I3338<= not (WX602 and WX529);
	I3339<= not (WX602 and I3338);
	I3340<= not (WX529 and I3338);
	I3351<= not (WX603 and WX531);
	I3352<= not (WX603 and I3351);
	I3353<= not (WX531 and I3351);
	I3364<= not (WX604 and WX533);
	I3365<= not (WX604 and I3364);
	I3366<= not (WX533 and I3364);
	I3377<= not (WX605 and WX535);
	I3378<= not (WX605 and I3377);
	I3379<= not (WX535 and I3377);
	I3390<= not (WX606 and WX537);
	I3391<= not (WX606 and I3390);
	I3392<= not (WX537 and I3390);
	I3403<= not (WX607 and WX539);
	I3404<= not (WX607 and I3403);
	I3405<= not (WX539 and I3403);
	I3416<= not (WX608 and WX541);
	I3417<= not (WX608 and I3416);
	I3418<= not (WX541 and I3416);
	I3429<= not (WX609 and WX543);
	I3430<= not (WX609 and I3429);
	I3431<= not (WX543 and I3429);
	I3442<= not (WX610 and WX545);
	I3443<= not (WX610 and I3442);
	I3444<= not (WX545 and I3442);
	I3455<= not (WX611 and WX547);
	I3456<= not (WX611 and I3455);
	I3457<= not (WX547 and I3455);
	I3469<= not (I3471 and I3472);
	I3470<= not (WX627 and CRC_OUT_9_31);
	I3471<= not (WX627 and I3470);
	I3472<= not (CRC_OUT_9_31 and I3470);
	I3477<= not (CRC_OUT_9_15 and I3469);
	I3478<= not (CRC_OUT_9_15 and I3477);
	I3479<= not (I3469 and I3477);
	I3484<= not (I3486 and I3487);
	I3485<= not (WX632 and CRC_OUT_9_31);
	I3486<= not (WX632 and I3485);
	I3487<= not (CRC_OUT_9_31 and I3485);
	I3492<= not (CRC_OUT_9_10 and I3484);
	I3493<= not (CRC_OUT_9_10 and I3492);
	I3494<= not (I3484 and I3492);
	I3499<= not (I3501 and I3502);
	I3500<= not (WX639 and CRC_OUT_9_31);
	I3501<= not (WX639 and I3500);
	I3502<= not (CRC_OUT_9_31 and I3500);
	I3507<= not (CRC_OUT_9_3 and I3499);
	I3508<= not (CRC_OUT_9_3 and I3507);
	I3509<= not (I3499 and I3507);
	I3514<= not (WX643 and CRC_OUT_9_31);
	I3515<= not (WX643 and I3514);
	I3516<= not (CRC_OUT_9_31 and I3514);
	I3521<= not (WX612 and CRC_OUT_9_30);
	I3522<= not (WX612 and I3521);
	I3523<= not (CRC_OUT_9_30 and I3521);
	I3528<= not (WX613 and CRC_OUT_9_29);
	I3529<= not (WX613 and I3528);
	I3530<= not (CRC_OUT_9_29 and I3528);
	I3535<= not (WX614 and CRC_OUT_9_28);
	I3536<= not (WX614 and I3535);
	I3537<= not (CRC_OUT_9_28 and I3535);
	I3542<= not (WX615 and CRC_OUT_9_27);
	I3543<= not (WX615 and I3542);
	I3544<= not (CRC_OUT_9_27 and I3542);
	I3549<= not (WX616 and CRC_OUT_9_26);
	I3550<= not (WX616 and I3549);
	I3551<= not (CRC_OUT_9_26 and I3549);
	I3556<= not (WX617 and CRC_OUT_9_25);
	I3557<= not (WX617 and I3556);
	I3558<= not (CRC_OUT_9_25 and I3556);
	I3563<= not (WX618 and CRC_OUT_9_24);
	I3564<= not (WX618 and I3563);
	I3565<= not (CRC_OUT_9_24 and I3563);
	I3570<= not (WX619 and CRC_OUT_9_23);
	I3571<= not (WX619 and I3570);
	I3572<= not (CRC_OUT_9_23 and I3570);
	I3577<= not (WX620 and CRC_OUT_9_22);
	I3578<= not (WX620 and I3577);
	I3579<= not (CRC_OUT_9_22 and I3577);
	I3584<= not (WX621 and CRC_OUT_9_21);
	I3585<= not (WX621 and I3584);
	I3586<= not (CRC_OUT_9_21 and I3584);
	I3591<= not (WX622 and CRC_OUT_9_20);
	I3592<= not (WX622 and I3591);
	I3593<= not (CRC_OUT_9_20 and I3591);
	I3598<= not (WX623 and CRC_OUT_9_19);
	I3599<= not (WX623 and I3598);
	I3600<= not (CRC_OUT_9_19 and I3598);
	I3605<= not (WX624 and CRC_OUT_9_18);
	I3606<= not (WX624 and I3605);
	I3607<= not (CRC_OUT_9_18 and I3605);
	I3612<= not (WX625 and CRC_OUT_9_17);
	I3613<= not (WX625 and I3612);
	I3614<= not (CRC_OUT_9_17 and I3612);
	I3619<= not (WX626 and CRC_OUT_9_16);
	I3620<= not (WX626 and I3619);
	I3621<= not (CRC_OUT_9_16 and I3619);
	I3626<= not (WX628 and CRC_OUT_9_14);
	I3627<= not (WX628 and I3626);
	I3628<= not (CRC_OUT_9_14 and I3626);
	I3633<= not (WX629 and CRC_OUT_9_13);
	I3634<= not (WX629 and I3633);
	I3635<= not (CRC_OUT_9_13 and I3633);
	I3640<= not (WX630 and CRC_OUT_9_12);
	I3641<= not (WX630 and I3640);
	I3642<= not (CRC_OUT_9_12 and I3640);
	I3647<= not (WX631 and CRC_OUT_9_11);
	I3648<= not (WX631 and I3647);
	I3649<= not (CRC_OUT_9_11 and I3647);
	I3654<= not (WX633 and CRC_OUT_9_9);
	I3655<= not (WX633 and I3654);
	I3656<= not (CRC_OUT_9_9 and I3654);
	I3661<= not (WX634 and CRC_OUT_9_8);
	I3662<= not (WX634 and I3661);
	I3663<= not (CRC_OUT_9_8 and I3661);
	I3668<= not (WX635 and CRC_OUT_9_7);
	I3669<= not (WX635 and I3668);
	I3670<= not (CRC_OUT_9_7 and I3668);
	I3675<= not (WX636 and CRC_OUT_9_6);
	I3676<= not (WX636 and I3675);
	I3677<= not (CRC_OUT_9_6 and I3675);
	I3682<= not (WX637 and CRC_OUT_9_5);
	I3683<= not (WX637 and I3682);
	I3684<= not (CRC_OUT_9_5 and I3682);
	I3689<= not (WX638 and CRC_OUT_9_4);
	I3690<= not (WX638 and I3689);
	I3691<= not (CRC_OUT_9_4 and I3689);
	I3696<= not (WX640 and CRC_OUT_9_2);
	I3697<= not (WX640 and I3696);
	I3698<= not (CRC_OUT_9_2 and I3696);
	I3703<= not (WX641 and CRC_OUT_9_1);
	I3704<= not (WX641 and I3703);
	I3705<= not (CRC_OUT_9_1 and I3703);
	I3710<= not (WX642 and CRC_OUT_9_0);
	I3711<= not (WX642 and I3710);
	I3712<= not (CRC_OUT_9_0 and I3710);
	I5991<= not (I6001 and I6002);
	I5992<= not (I5994 and I5995);
	I5993<= not (WX2294 and WX1938);
	I5994<= not (WX2294 and I5993);
	I5995<= not (WX1938 and I5993);
	I6000<= not (WX2002 and I5992);
	I6001<= not (WX2002 and I6000);
	I6002<= not (I5992 and I6000);
	I6007<= not (I6009 and I6010);
	I6008<= not (WX2066 and WX2130);
	I6009<= not (WX2066 and I6008);
	I6010<= not (WX2130 and I6008);
	I6015<= not (I5991 and I6007);
	I6016<= not (I5991 and I6015);
	I6017<= not (I6007 and I6015);
	I6022<= not (I6032 and I6033);
	I6023<= not (I6025 and I6026);
	I6024<= not (WX2294 and WX1940);
	I6025<= not (WX2294 and I6024);
	I6026<= not (WX1940 and I6024);
	I6031<= not (WX2004 and I6023);
	I6032<= not (WX2004 and I6031);
	I6033<= not (I6023 and I6031);
	I6038<= not (I6040 and I6041);
	I6039<= not (WX2068 and WX2132);
	I6040<= not (WX2068 and I6039);
	I6041<= not (WX2132 and I6039);
	I6046<= not (I6022 and I6038);
	I6047<= not (I6022 and I6046);
	I6048<= not (I6038 and I6046);
	I6053<= not (I6063 and I6064);
	I6054<= not (I6056 and I6057);
	I6055<= not (WX2294 and WX1942);
	I6056<= not (WX2294 and I6055);
	I6057<= not (WX1942 and I6055);
	I6062<= not (WX2006 and I6054);
	I6063<= not (WX2006 and I6062);
	I6064<= not (I6054 and I6062);
	I6069<= not (I6071 and I6072);
	I6070<= not (WX2070 and WX2134);
	I6071<= not (WX2070 and I6070);
	I6072<= not (WX2134 and I6070);
	I6077<= not (I6053 and I6069);
	I6078<= not (I6053 and I6077);
	I6079<= not (I6069 and I6077);
	I6084<= not (I6094 and I6095);
	I6085<= not (I6087 and I6088);
	I6086<= not (WX2294 and WX1944);
	I6087<= not (WX2294 and I6086);
	I6088<= not (WX1944 and I6086);
	I6093<= not (WX2008 and I6085);
	I6094<= not (WX2008 and I6093);
	I6095<= not (I6085 and I6093);
	I6100<= not (I6102 and I6103);
	I6101<= not (WX2072 and WX2136);
	I6102<= not (WX2072 and I6101);
	I6103<= not (WX2136 and I6101);
	I6108<= not (I6084 and I6100);
	I6109<= not (I6084 and I6108);
	I6110<= not (I6100 and I6108);
	I6115<= not (I6125 and I6126);
	I6116<= not (I6118 and I6119);
	I6117<= not (WX2294 and WX1946);
	I6118<= not (WX2294 and I6117);
	I6119<= not (WX1946 and I6117);
	I6124<= not (WX2010 and I6116);
	I6125<= not (WX2010 and I6124);
	I6126<= not (I6116 and I6124);
	I6131<= not (I6133 and I6134);
	I6132<= not (WX2074 and WX2138);
	I6133<= not (WX2074 and I6132);
	I6134<= not (WX2138 and I6132);
	I6139<= not (I6115 and I6131);
	I6140<= not (I6115 and I6139);
	I6141<= not (I6131 and I6139);
	I6146<= not (I6156 and I6157);
	I6147<= not (I6149 and I6150);
	I6148<= not (WX2294 and WX1948);
	I6149<= not (WX2294 and I6148);
	I6150<= not (WX1948 and I6148);
	I6155<= not (WX2012 and I6147);
	I6156<= not (WX2012 and I6155);
	I6157<= not (I6147 and I6155);
	I6162<= not (I6164 and I6165);
	I6163<= not (WX2076 and WX2140);
	I6164<= not (WX2076 and I6163);
	I6165<= not (WX2140 and I6163);
	I6170<= not (I6146 and I6162);
	I6171<= not (I6146 and I6170);
	I6172<= not (I6162 and I6170);
	I6177<= not (I6187 and I6188);
	I6178<= not (I6180 and I6181);
	I6179<= not (WX2294 and WX1950);
	I6180<= not (WX2294 and I6179);
	I6181<= not (WX1950 and I6179);
	I6186<= not (WX2014 and I6178);
	I6187<= not (WX2014 and I6186);
	I6188<= not (I6178 and I6186);
	I6193<= not (I6195 and I6196);
	I6194<= not (WX2078 and WX2142);
	I6195<= not (WX2078 and I6194);
	I6196<= not (WX2142 and I6194);
	I6201<= not (I6177 and I6193);
	I6202<= not (I6177 and I6201);
	I6203<= not (I6193 and I6201);
	I6208<= not (I6218 and I6219);
	I6209<= not (I6211 and I6212);
	I6210<= not (WX2294 and WX1952);
	I6211<= not (WX2294 and I6210);
	I6212<= not (WX1952 and I6210);
	I6217<= not (WX2016 and I6209);
	I6218<= not (WX2016 and I6217);
	I6219<= not (I6209 and I6217);
	I6224<= not (I6226 and I6227);
	I6225<= not (WX2080 and WX2144);
	I6226<= not (WX2080 and I6225);
	I6227<= not (WX2144 and I6225);
	I6232<= not (I6208 and I6224);
	I6233<= not (I6208 and I6232);
	I6234<= not (I6224 and I6232);
	I6239<= not (I6249 and I6250);
	I6240<= not (I6242 and I6243);
	I6241<= not (WX2294 and WX1954);
	I6242<= not (WX2294 and I6241);
	I6243<= not (WX1954 and I6241);
	I6248<= not (WX2018 and I6240);
	I6249<= not (WX2018 and I6248);
	I6250<= not (I6240 and I6248);
	I6255<= not (I6257 and I6258);
	I6256<= not (WX2082 and WX2146);
	I6257<= not (WX2082 and I6256);
	I6258<= not (WX2146 and I6256);
	I6263<= not (I6239 and I6255);
	I6264<= not (I6239 and I6263);
	I6265<= not (I6255 and I6263);
	I6270<= not (I6280 and I6281);
	I6271<= not (I6273 and I6274);
	I6272<= not (WX2294 and WX1956);
	I6273<= not (WX2294 and I6272);
	I6274<= not (WX1956 and I6272);
	I6279<= not (WX2020 and I6271);
	I6280<= not (WX2020 and I6279);
	I6281<= not (I6271 and I6279);
	I6286<= not (I6288 and I6289);
	I6287<= not (WX2084 and WX2148);
	I6288<= not (WX2084 and I6287);
	I6289<= not (WX2148 and I6287);
	I6294<= not (I6270 and I6286);
	I6295<= not (I6270 and I6294);
	I6296<= not (I6286 and I6294);
	I6301<= not (I6311 and I6312);
	I6302<= not (I6304 and I6305);
	I6303<= not (WX2294 and WX1958);
	I6304<= not (WX2294 and I6303);
	I6305<= not (WX1958 and I6303);
	I6310<= not (WX2022 and I6302);
	I6311<= not (WX2022 and I6310);
	I6312<= not (I6302 and I6310);
	I6317<= not (I6319 and I6320);
	I6318<= not (WX2086 and WX2150);
	I6319<= not (WX2086 and I6318);
	I6320<= not (WX2150 and I6318);
	I6325<= not (I6301 and I6317);
	I6326<= not (I6301 and I6325);
	I6327<= not (I6317 and I6325);
	I6332<= not (I6342 and I6343);
	I6333<= not (I6335 and I6336);
	I6334<= not (WX2294 and WX1960);
	I6335<= not (WX2294 and I6334);
	I6336<= not (WX1960 and I6334);
	I6341<= not (WX2024 and I6333);
	I6342<= not (WX2024 and I6341);
	I6343<= not (I6333 and I6341);
	I6348<= not (I6350 and I6351);
	I6349<= not (WX2088 and WX2152);
	I6350<= not (WX2088 and I6349);
	I6351<= not (WX2152 and I6349);
	I6356<= not (I6332 and I6348);
	I6357<= not (I6332 and I6356);
	I6358<= not (I6348 and I6356);
	I6363<= not (I6373 and I6374);
	I6364<= not (I6366 and I6367);
	I6365<= not (WX2294 and WX1962);
	I6366<= not (WX2294 and I6365);
	I6367<= not (WX1962 and I6365);
	I6372<= not (WX2026 and I6364);
	I6373<= not (WX2026 and I6372);
	I6374<= not (I6364 and I6372);
	I6379<= not (I6381 and I6382);
	I6380<= not (WX2090 and WX2154);
	I6381<= not (WX2090 and I6380);
	I6382<= not (WX2154 and I6380);
	I6387<= not (I6363 and I6379);
	I6388<= not (I6363 and I6387);
	I6389<= not (I6379 and I6387);
	I6394<= not (I6404 and I6405);
	I6395<= not (I6397 and I6398);
	I6396<= not (WX2294 and WX1964);
	I6397<= not (WX2294 and I6396);
	I6398<= not (WX1964 and I6396);
	I6403<= not (WX2028 and I6395);
	I6404<= not (WX2028 and I6403);
	I6405<= not (I6395 and I6403);
	I6410<= not (I6412 and I6413);
	I6411<= not (WX2092 and WX2156);
	I6412<= not (WX2092 and I6411);
	I6413<= not (WX2156 and I6411);
	I6418<= not (I6394 and I6410);
	I6419<= not (I6394 and I6418);
	I6420<= not (I6410 and I6418);
	I6425<= not (I6435 and I6436);
	I6426<= not (I6428 and I6429);
	I6427<= not (WX2294 and WX1966);
	I6428<= not (WX2294 and I6427);
	I6429<= not (WX1966 and I6427);
	I6434<= not (WX2030 and I6426);
	I6435<= not (WX2030 and I6434);
	I6436<= not (I6426 and I6434);
	I6441<= not (I6443 and I6444);
	I6442<= not (WX2094 and WX2158);
	I6443<= not (WX2094 and I6442);
	I6444<= not (WX2158 and I6442);
	I6449<= not (I6425 and I6441);
	I6450<= not (I6425 and I6449);
	I6451<= not (I6441 and I6449);
	I6456<= not (I6466 and I6467);
	I6457<= not (I6459 and I6460);
	I6458<= not (WX2294 and WX1968);
	I6459<= not (WX2294 and I6458);
	I6460<= not (WX1968 and I6458);
	I6465<= not (WX2032 and I6457);
	I6466<= not (WX2032 and I6465);
	I6467<= not (I6457 and I6465);
	I6472<= not (I6474 and I6475);
	I6473<= not (WX2096 and WX2160);
	I6474<= not (WX2096 and I6473);
	I6475<= not (WX2160 and I6473);
	I6480<= not (I6456 and I6472);
	I6481<= not (I6456 and I6480);
	I6482<= not (I6472 and I6480);
	I6487<= not (I6497 and I6498);
	I6488<= not (I6490 and I6491);
	I6489<= not (WX2295 and WX1970);
	I6490<= not (WX2295 and I6489);
	I6491<= not (WX1970 and I6489);
	I6496<= not (WX2034 and I6488);
	I6497<= not (WX2034 and I6496);
	I6498<= not (I6488 and I6496);
	I6503<= not (I6505 and I6506);
	I6504<= not (WX2098 and WX2162);
	I6505<= not (WX2098 and I6504);
	I6506<= not (WX2162 and I6504);
	I6511<= not (I6487 and I6503);
	I6512<= not (I6487 and I6511);
	I6513<= not (I6503 and I6511);
	I6518<= not (I6528 and I6529);
	I6519<= not (I6521 and I6522);
	I6520<= not (WX2295 and WX1972);
	I6521<= not (WX2295 and I6520);
	I6522<= not (WX1972 and I6520);
	I6527<= not (WX2036 and I6519);
	I6528<= not (WX2036 and I6527);
	I6529<= not (I6519 and I6527);
	I6534<= not (I6536 and I6537);
	I6535<= not (WX2100 and WX2164);
	I6536<= not (WX2100 and I6535);
	I6537<= not (WX2164 and I6535);
	I6542<= not (I6518 and I6534);
	I6543<= not (I6518 and I6542);
	I6544<= not (I6534 and I6542);
	I6549<= not (I6559 and I6560);
	I6550<= not (I6552 and I6553);
	I6551<= not (WX2295 and WX1974);
	I6552<= not (WX2295 and I6551);
	I6553<= not (WX1974 and I6551);
	I6558<= not (WX2038 and I6550);
	I6559<= not (WX2038 and I6558);
	I6560<= not (I6550 and I6558);
	I6565<= not (I6567 and I6568);
	I6566<= not (WX2102 and WX2166);
	I6567<= not (WX2102 and I6566);
	I6568<= not (WX2166 and I6566);
	I6573<= not (I6549 and I6565);
	I6574<= not (I6549 and I6573);
	I6575<= not (I6565 and I6573);
	I6580<= not (I6590 and I6591);
	I6581<= not (I6583 and I6584);
	I6582<= not (WX2295 and WX1976);
	I6583<= not (WX2295 and I6582);
	I6584<= not (WX1976 and I6582);
	I6589<= not (WX2040 and I6581);
	I6590<= not (WX2040 and I6589);
	I6591<= not (I6581 and I6589);
	I6596<= not (I6598 and I6599);
	I6597<= not (WX2104 and WX2168);
	I6598<= not (WX2104 and I6597);
	I6599<= not (WX2168 and I6597);
	I6604<= not (I6580 and I6596);
	I6605<= not (I6580 and I6604);
	I6606<= not (I6596 and I6604);
	I6611<= not (I6621 and I6622);
	I6612<= not (I6614 and I6615);
	I6613<= not (WX2295 and WX1978);
	I6614<= not (WX2295 and I6613);
	I6615<= not (WX1978 and I6613);
	I6620<= not (WX2042 and I6612);
	I6621<= not (WX2042 and I6620);
	I6622<= not (I6612 and I6620);
	I6627<= not (I6629 and I6630);
	I6628<= not (WX2106 and WX2170);
	I6629<= not (WX2106 and I6628);
	I6630<= not (WX2170 and I6628);
	I6635<= not (I6611 and I6627);
	I6636<= not (I6611 and I6635);
	I6637<= not (I6627 and I6635);
	I6642<= not (I6652 and I6653);
	I6643<= not (I6645 and I6646);
	I6644<= not (WX2295 and WX1980);
	I6645<= not (WX2295 and I6644);
	I6646<= not (WX1980 and I6644);
	I6651<= not (WX2044 and I6643);
	I6652<= not (WX2044 and I6651);
	I6653<= not (I6643 and I6651);
	I6658<= not (I6660 and I6661);
	I6659<= not (WX2108 and WX2172);
	I6660<= not (WX2108 and I6659);
	I6661<= not (WX2172 and I6659);
	I6666<= not (I6642 and I6658);
	I6667<= not (I6642 and I6666);
	I6668<= not (I6658 and I6666);
	I6673<= not (I6683 and I6684);
	I6674<= not (I6676 and I6677);
	I6675<= not (WX2295 and WX1982);
	I6676<= not (WX2295 and I6675);
	I6677<= not (WX1982 and I6675);
	I6682<= not (WX2046 and I6674);
	I6683<= not (WX2046 and I6682);
	I6684<= not (I6674 and I6682);
	I6689<= not (I6691 and I6692);
	I6690<= not (WX2110 and WX2174);
	I6691<= not (WX2110 and I6690);
	I6692<= not (WX2174 and I6690);
	I6697<= not (I6673 and I6689);
	I6698<= not (I6673 and I6697);
	I6699<= not (I6689 and I6697);
	I6704<= not (I6714 and I6715);
	I6705<= not (I6707 and I6708);
	I6706<= not (WX2295 and WX1984);
	I6707<= not (WX2295 and I6706);
	I6708<= not (WX1984 and I6706);
	I6713<= not (WX2048 and I6705);
	I6714<= not (WX2048 and I6713);
	I6715<= not (I6705 and I6713);
	I6720<= not (I6722 and I6723);
	I6721<= not (WX2112 and WX2176);
	I6722<= not (WX2112 and I6721);
	I6723<= not (WX2176 and I6721);
	I6728<= not (I6704 and I6720);
	I6729<= not (I6704 and I6728);
	I6730<= not (I6720 and I6728);
	I6735<= not (I6745 and I6746);
	I6736<= not (I6738 and I6739);
	I6737<= not (WX2295 and WX1986);
	I6738<= not (WX2295 and I6737);
	I6739<= not (WX1986 and I6737);
	I6744<= not (WX2050 and I6736);
	I6745<= not (WX2050 and I6744);
	I6746<= not (I6736 and I6744);
	I6751<= not (I6753 and I6754);
	I6752<= not (WX2114 and WX2178);
	I6753<= not (WX2114 and I6752);
	I6754<= not (WX2178 and I6752);
	I6759<= not (I6735 and I6751);
	I6760<= not (I6735 and I6759);
	I6761<= not (I6751 and I6759);
	I6766<= not (I6776 and I6777);
	I6767<= not (I6769 and I6770);
	I6768<= not (WX2295 and WX1988);
	I6769<= not (WX2295 and I6768);
	I6770<= not (WX1988 and I6768);
	I6775<= not (WX2052 and I6767);
	I6776<= not (WX2052 and I6775);
	I6777<= not (I6767 and I6775);
	I6782<= not (I6784 and I6785);
	I6783<= not (WX2116 and WX2180);
	I6784<= not (WX2116 and I6783);
	I6785<= not (WX2180 and I6783);
	I6790<= not (I6766 and I6782);
	I6791<= not (I6766 and I6790);
	I6792<= not (I6782 and I6790);
	I6797<= not (I6807 and I6808);
	I6798<= not (I6800 and I6801);
	I6799<= not (WX2295 and WX1990);
	I6800<= not (WX2295 and I6799);
	I6801<= not (WX1990 and I6799);
	I6806<= not (WX2054 and I6798);
	I6807<= not (WX2054 and I6806);
	I6808<= not (I6798 and I6806);
	I6813<= not (I6815 and I6816);
	I6814<= not (WX2118 and WX2182);
	I6815<= not (WX2118 and I6814);
	I6816<= not (WX2182 and I6814);
	I6821<= not (I6797 and I6813);
	I6822<= not (I6797 and I6821);
	I6823<= not (I6813 and I6821);
	I6828<= not (I6838 and I6839);
	I6829<= not (I6831 and I6832);
	I6830<= not (WX2295 and WX1992);
	I6831<= not (WX2295 and I6830);
	I6832<= not (WX1992 and I6830);
	I6837<= not (WX2056 and I6829);
	I6838<= not (WX2056 and I6837);
	I6839<= not (I6829 and I6837);
	I6844<= not (I6846 and I6847);
	I6845<= not (WX2120 and WX2184);
	I6846<= not (WX2120 and I6845);
	I6847<= not (WX2184 and I6845);
	I6852<= not (I6828 and I6844);
	I6853<= not (I6828 and I6852);
	I6854<= not (I6844 and I6852);
	I6859<= not (I6869 and I6870);
	I6860<= not (I6862 and I6863);
	I6861<= not (WX2295 and WX1994);
	I6862<= not (WX2295 and I6861);
	I6863<= not (WX1994 and I6861);
	I6868<= not (WX2058 and I6860);
	I6869<= not (WX2058 and I6868);
	I6870<= not (I6860 and I6868);
	I6875<= not (I6877 and I6878);
	I6876<= not (WX2122 and WX2186);
	I6877<= not (WX2122 and I6876);
	I6878<= not (WX2186 and I6876);
	I6883<= not (I6859 and I6875);
	I6884<= not (I6859 and I6883);
	I6885<= not (I6875 and I6883);
	I6890<= not (I6900 and I6901);
	I6891<= not (I6893 and I6894);
	I6892<= not (WX2295 and WX1996);
	I6893<= not (WX2295 and I6892);
	I6894<= not (WX1996 and I6892);
	I6899<= not (WX2060 and I6891);
	I6900<= not (WX2060 and I6899);
	I6901<= not (I6891 and I6899);
	I6906<= not (I6908 and I6909);
	I6907<= not (WX2124 and WX2188);
	I6908<= not (WX2124 and I6907);
	I6909<= not (WX2188 and I6907);
	I6914<= not (I6890 and I6906);
	I6915<= not (I6890 and I6914);
	I6916<= not (I6906 and I6914);
	I6921<= not (I6931 and I6932);
	I6922<= not (I6924 and I6925);
	I6923<= not (WX2295 and WX1998);
	I6924<= not (WX2295 and I6923);
	I6925<= not (WX1998 and I6923);
	I6930<= not (WX2062 and I6922);
	I6931<= not (WX2062 and I6930);
	I6932<= not (I6922 and I6930);
	I6937<= not (I6939 and I6940);
	I6938<= not (WX2126 and WX2190);
	I6939<= not (WX2126 and I6938);
	I6940<= not (WX2190 and I6938);
	I6945<= not (I6921 and I6937);
	I6946<= not (I6921 and I6945);
	I6947<= not (I6937 and I6945);
	I6952<= not (I6962 and I6963);
	I6953<= not (I6955 and I6956);
	I6954<= not (WX2295 and WX2000);
	I6955<= not (WX2295 and I6954);
	I6956<= not (WX2000 and I6954);
	I6961<= not (WX2064 and I6953);
	I6962<= not (WX2064 and I6961);
	I6963<= not (I6953 and I6961);
	I6968<= not (I6970 and I6971);
	I6969<= not (WX2128 and WX2192);
	I6970<= not (WX2128 and I6969);
	I6971<= not (WX2192 and I6969);
	I6976<= not (I6952 and I6968);
	I6977<= not (I6952 and I6976);
	I6978<= not (I6968 and I6976);
	I7057<= not (WX1873 and WX1778);
	I7058<= not (WX1873 and I7057);
	I7059<= not (WX1778 and I7057);
	I7070<= not (WX1874 and WX1780);
	I7071<= not (WX1874 and I7070);
	I7072<= not (WX1780 and I7070);
	I7083<= not (WX1875 and WX1782);
	I7084<= not (WX1875 and I7083);
	I7085<= not (WX1782 and I7083);
	I7096<= not (WX1876 and WX1784);
	I7097<= not (WX1876 and I7096);
	I7098<= not (WX1784 and I7096);
	I7109<= not (WX1877 and WX1786);
	I7110<= not (WX1877 and I7109);
	I7111<= not (WX1786 and I7109);
	I7122<= not (WX1878 and WX1788);
	I7123<= not (WX1878 and I7122);
	I7124<= not (WX1788 and I7122);
	I7135<= not (WX1879 and WX1790);
	I7136<= not (WX1879 and I7135);
	I7137<= not (WX1790 and I7135);
	I7148<= not (WX1880 and WX1792);
	I7149<= not (WX1880 and I7148);
	I7150<= not (WX1792 and I7148);
	I7161<= not (WX1881 and WX1794);
	I7162<= not (WX1881 and I7161);
	I7163<= not (WX1794 and I7161);
	I7174<= not (WX1882 and WX1796);
	I7175<= not (WX1882 and I7174);
	I7176<= not (WX1796 and I7174);
	I7187<= not (WX1883 and WX1798);
	I7188<= not (WX1883 and I7187);
	I7189<= not (WX1798 and I7187);
	I7200<= not (WX1884 and WX1800);
	I7201<= not (WX1884 and I7200);
	I7202<= not (WX1800 and I7200);
	I7213<= not (WX1885 and WX1802);
	I7214<= not (WX1885 and I7213);
	I7215<= not (WX1802 and I7213);
	I7226<= not (WX1886 and WX1804);
	I7227<= not (WX1886 and I7226);
	I7228<= not (WX1804 and I7226);
	I7239<= not (WX1887 and WX1806);
	I7240<= not (WX1887 and I7239);
	I7241<= not (WX1806 and I7239);
	I7252<= not (WX1888 and WX1808);
	I7253<= not (WX1888 and I7252);
	I7254<= not (WX1808 and I7252);
	I7265<= not (WX1889 and WX1810);
	I7266<= not (WX1889 and I7265);
	I7267<= not (WX1810 and I7265);
	I7278<= not (WX1890 and WX1812);
	I7279<= not (WX1890 and I7278);
	I7280<= not (WX1812 and I7278);
	I7291<= not (WX1891 and WX1814);
	I7292<= not (WX1891 and I7291);
	I7293<= not (WX1814 and I7291);
	I7304<= not (WX1892 and WX1816);
	I7305<= not (WX1892 and I7304);
	I7306<= not (WX1816 and I7304);
	I7317<= not (WX1893 and WX1818);
	I7318<= not (WX1893 and I7317);
	I7319<= not (WX1818 and I7317);
	I7330<= not (WX1894 and WX1820);
	I7331<= not (WX1894 and I7330);
	I7332<= not (WX1820 and I7330);
	I7343<= not (WX1895 and WX1822);
	I7344<= not (WX1895 and I7343);
	I7345<= not (WX1822 and I7343);
	I7356<= not (WX1896 and WX1824);
	I7357<= not (WX1896 and I7356);
	I7358<= not (WX1824 and I7356);
	I7369<= not (WX1897 and WX1826);
	I7370<= not (WX1897 and I7369);
	I7371<= not (WX1826 and I7369);
	I7382<= not (WX1898 and WX1828);
	I7383<= not (WX1898 and I7382);
	I7384<= not (WX1828 and I7382);
	I7395<= not (WX1899 and WX1830);
	I7396<= not (WX1899 and I7395);
	I7397<= not (WX1830 and I7395);
	I7408<= not (WX1900 and WX1832);
	I7409<= not (WX1900 and I7408);
	I7410<= not (WX1832 and I7408);
	I7421<= not (WX1901 and WX1834);
	I7422<= not (WX1901 and I7421);
	I7423<= not (WX1834 and I7421);
	I7434<= not (WX1902 and WX1836);
	I7435<= not (WX1902 and I7434);
	I7436<= not (WX1836 and I7434);
	I7447<= not (WX1903 and WX1838);
	I7448<= not (WX1903 and I7447);
	I7449<= not (WX1838 and I7447);
	I7460<= not (WX1904 and WX1840);
	I7461<= not (WX1904 and I7460);
	I7462<= not (WX1840 and I7460);
	I7474<= not (I7476 and I7477);
	I7475<= not (WX1920 and CRC_OUT_8_31);
	I7476<= not (WX1920 and I7475);
	I7477<= not (CRC_OUT_8_31 and I7475);
	I7482<= not (CRC_OUT_8_15 and I7474);
	I7483<= not (CRC_OUT_8_15 and I7482);
	I7484<= not (I7474 and I7482);
	I7489<= not (I7491 and I7492);
	I7490<= not (WX1925 and CRC_OUT_8_31);
	I7491<= not (WX1925 and I7490);
	I7492<= not (CRC_OUT_8_31 and I7490);
	I7497<= not (CRC_OUT_8_10 and I7489);
	I7498<= not (CRC_OUT_8_10 and I7497);
	I7499<= not (I7489 and I7497);
	I7504<= not (I7506 and I7507);
	I7505<= not (WX1932 and CRC_OUT_8_31);
	I7506<= not (WX1932 and I7505);
	I7507<= not (CRC_OUT_8_31 and I7505);
	I7512<= not (CRC_OUT_8_3 and I7504);
	I7513<= not (CRC_OUT_8_3 and I7512);
	I7514<= not (I7504 and I7512);
	I7519<= not (WX1936 and CRC_OUT_8_31);
	I7520<= not (WX1936 and I7519);
	I7521<= not (CRC_OUT_8_31 and I7519);
	I7526<= not (WX1905 and CRC_OUT_8_30);
	I7527<= not (WX1905 and I7526);
	I7528<= not (CRC_OUT_8_30 and I7526);
	I7533<= not (WX1906 and CRC_OUT_8_29);
	I7534<= not (WX1906 and I7533);
	I7535<= not (CRC_OUT_8_29 and I7533);
	I7540<= not (WX1907 and CRC_OUT_8_28);
	I7541<= not (WX1907 and I7540);
	I7542<= not (CRC_OUT_8_28 and I7540);
	I7547<= not (WX1908 and CRC_OUT_8_27);
	I7548<= not (WX1908 and I7547);
	I7549<= not (CRC_OUT_8_27 and I7547);
	I7554<= not (WX1909 and CRC_OUT_8_26);
	I7555<= not (WX1909 and I7554);
	I7556<= not (CRC_OUT_8_26 and I7554);
	I7561<= not (WX1910 and CRC_OUT_8_25);
	I7562<= not (WX1910 and I7561);
	I7563<= not (CRC_OUT_8_25 and I7561);
	I7568<= not (WX1911 and CRC_OUT_8_24);
	I7569<= not (WX1911 and I7568);
	I7570<= not (CRC_OUT_8_24 and I7568);
	I7575<= not (WX1912 and CRC_OUT_8_23);
	I7576<= not (WX1912 and I7575);
	I7577<= not (CRC_OUT_8_23 and I7575);
	I7582<= not (WX1913 and CRC_OUT_8_22);
	I7583<= not (WX1913 and I7582);
	I7584<= not (CRC_OUT_8_22 and I7582);
	I7589<= not (WX1914 and CRC_OUT_8_21);
	I7590<= not (WX1914 and I7589);
	I7591<= not (CRC_OUT_8_21 and I7589);
	I7596<= not (WX1915 and CRC_OUT_8_20);
	I7597<= not (WX1915 and I7596);
	I7598<= not (CRC_OUT_8_20 and I7596);
	I7603<= not (WX1916 and CRC_OUT_8_19);
	I7604<= not (WX1916 and I7603);
	I7605<= not (CRC_OUT_8_19 and I7603);
	I7610<= not (WX1917 and CRC_OUT_8_18);
	I7611<= not (WX1917 and I7610);
	I7612<= not (CRC_OUT_8_18 and I7610);
	I7617<= not (WX1918 and CRC_OUT_8_17);
	I7618<= not (WX1918 and I7617);
	I7619<= not (CRC_OUT_8_17 and I7617);
	I7624<= not (WX1919 and CRC_OUT_8_16);
	I7625<= not (WX1919 and I7624);
	I7626<= not (CRC_OUT_8_16 and I7624);
	I7631<= not (WX1921 and CRC_OUT_8_14);
	I7632<= not (WX1921 and I7631);
	I7633<= not (CRC_OUT_8_14 and I7631);
	I7638<= not (WX1922 and CRC_OUT_8_13);
	I7639<= not (WX1922 and I7638);
	I7640<= not (CRC_OUT_8_13 and I7638);
	I7645<= not (WX1923 and CRC_OUT_8_12);
	I7646<= not (WX1923 and I7645);
	I7647<= not (CRC_OUT_8_12 and I7645);
	I7652<= not (WX1924 and CRC_OUT_8_11);
	I7653<= not (WX1924 and I7652);
	I7654<= not (CRC_OUT_8_11 and I7652);
	I7659<= not (WX1926 and CRC_OUT_8_9);
	I7660<= not (WX1926 and I7659);
	I7661<= not (CRC_OUT_8_9 and I7659);
	I7666<= not (WX1927 and CRC_OUT_8_8);
	I7667<= not (WX1927 and I7666);
	I7668<= not (CRC_OUT_8_8 and I7666);
	I7673<= not (WX1928 and CRC_OUT_8_7);
	I7674<= not (WX1928 and I7673);
	I7675<= not (CRC_OUT_8_7 and I7673);
	I7680<= not (WX1929 and CRC_OUT_8_6);
	I7681<= not (WX1929 and I7680);
	I7682<= not (CRC_OUT_8_6 and I7680);
	I7687<= not (WX1930 and CRC_OUT_8_5);
	I7688<= not (WX1930 and I7687);
	I7689<= not (CRC_OUT_8_5 and I7687);
	I7694<= not (WX1931 and CRC_OUT_8_4);
	I7695<= not (WX1931 and I7694);
	I7696<= not (CRC_OUT_8_4 and I7694);
	I7701<= not (WX1933 and CRC_OUT_8_2);
	I7702<= not (WX1933 and I7701);
	I7703<= not (CRC_OUT_8_2 and I7701);
	I7708<= not (WX1934 and CRC_OUT_8_1);
	I7709<= not (WX1934 and I7708);
	I7710<= not (CRC_OUT_8_1 and I7708);
	I7715<= not (WX1935 and CRC_OUT_8_0);
	I7716<= not (WX1935 and I7715);
	I7717<= not (CRC_OUT_8_0 and I7715);
	I9996<= not (I10006 and I10007);
	I9997<= not (I9999 and I10000);
	I9998<= not (WX3587 and WX3231);
	I9999<= not (WX3587 and I9998);
	I10000<= not (WX3231 and I9998);
	I10005<= not (WX3295 and I9997);
	I10006<= not (WX3295 and I10005);
	I10007<= not (I9997 and I10005);
	I10012<= not (I10014 and I10015);
	I10013<= not (WX3359 and WX3423);
	I10014<= not (WX3359 and I10013);
	I10015<= not (WX3423 and I10013);
	I10020<= not (I9996 and I10012);
	I10021<= not (I9996 and I10020);
	I10022<= not (I10012 and I10020);
	I10027<= not (I10037 and I10038);
	I10028<= not (I10030 and I10031);
	I10029<= not (WX3587 and WX3233);
	I10030<= not (WX3587 and I10029);
	I10031<= not (WX3233 and I10029);
	I10036<= not (WX3297 and I10028);
	I10037<= not (WX3297 and I10036);
	I10038<= not (I10028 and I10036);
	I10043<= not (I10045 and I10046);
	I10044<= not (WX3361 and WX3425);
	I10045<= not (WX3361 and I10044);
	I10046<= not (WX3425 and I10044);
	I10051<= not (I10027 and I10043);
	I10052<= not (I10027 and I10051);
	I10053<= not (I10043 and I10051);
	I10058<= not (I10068 and I10069);
	I10059<= not (I10061 and I10062);
	I10060<= not (WX3587 and WX3235);
	I10061<= not (WX3587 and I10060);
	I10062<= not (WX3235 and I10060);
	I10067<= not (WX3299 and I10059);
	I10068<= not (WX3299 and I10067);
	I10069<= not (I10059 and I10067);
	I10074<= not (I10076 and I10077);
	I10075<= not (WX3363 and WX3427);
	I10076<= not (WX3363 and I10075);
	I10077<= not (WX3427 and I10075);
	I10082<= not (I10058 and I10074);
	I10083<= not (I10058 and I10082);
	I10084<= not (I10074 and I10082);
	I10089<= not (I10099 and I10100);
	I10090<= not (I10092 and I10093);
	I10091<= not (WX3587 and WX3237);
	I10092<= not (WX3587 and I10091);
	I10093<= not (WX3237 and I10091);
	I10098<= not (WX3301 and I10090);
	I10099<= not (WX3301 and I10098);
	I10100<= not (I10090 and I10098);
	I10105<= not (I10107 and I10108);
	I10106<= not (WX3365 and WX3429);
	I10107<= not (WX3365 and I10106);
	I10108<= not (WX3429 and I10106);
	I10113<= not (I10089 and I10105);
	I10114<= not (I10089 and I10113);
	I10115<= not (I10105 and I10113);
	I10120<= not (I10130 and I10131);
	I10121<= not (I10123 and I10124);
	I10122<= not (WX3587 and WX3239);
	I10123<= not (WX3587 and I10122);
	I10124<= not (WX3239 and I10122);
	I10129<= not (WX3303 and I10121);
	I10130<= not (WX3303 and I10129);
	I10131<= not (I10121 and I10129);
	I10136<= not (I10138 and I10139);
	I10137<= not (WX3367 and WX3431);
	I10138<= not (WX3367 and I10137);
	I10139<= not (WX3431 and I10137);
	I10144<= not (I10120 and I10136);
	I10145<= not (I10120 and I10144);
	I10146<= not (I10136 and I10144);
	I10151<= not (I10161 and I10162);
	I10152<= not (I10154 and I10155);
	I10153<= not (WX3587 and WX3241);
	I10154<= not (WX3587 and I10153);
	I10155<= not (WX3241 and I10153);
	I10160<= not (WX3305 and I10152);
	I10161<= not (WX3305 and I10160);
	I10162<= not (I10152 and I10160);
	I10167<= not (I10169 and I10170);
	I10168<= not (WX3369 and WX3433);
	I10169<= not (WX3369 and I10168);
	I10170<= not (WX3433 and I10168);
	I10175<= not (I10151 and I10167);
	I10176<= not (I10151 and I10175);
	I10177<= not (I10167 and I10175);
	I10182<= not (I10192 and I10193);
	I10183<= not (I10185 and I10186);
	I10184<= not (WX3587 and WX3243);
	I10185<= not (WX3587 and I10184);
	I10186<= not (WX3243 and I10184);
	I10191<= not (WX3307 and I10183);
	I10192<= not (WX3307 and I10191);
	I10193<= not (I10183 and I10191);
	I10198<= not (I10200 and I10201);
	I10199<= not (WX3371 and WX3435);
	I10200<= not (WX3371 and I10199);
	I10201<= not (WX3435 and I10199);
	I10206<= not (I10182 and I10198);
	I10207<= not (I10182 and I10206);
	I10208<= not (I10198 and I10206);
	I10213<= not (I10223 and I10224);
	I10214<= not (I10216 and I10217);
	I10215<= not (WX3587 and WX3245);
	I10216<= not (WX3587 and I10215);
	I10217<= not (WX3245 and I10215);
	I10222<= not (WX3309 and I10214);
	I10223<= not (WX3309 and I10222);
	I10224<= not (I10214 and I10222);
	I10229<= not (I10231 and I10232);
	I10230<= not (WX3373 and WX3437);
	I10231<= not (WX3373 and I10230);
	I10232<= not (WX3437 and I10230);
	I10237<= not (I10213 and I10229);
	I10238<= not (I10213 and I10237);
	I10239<= not (I10229 and I10237);
	I10244<= not (I10254 and I10255);
	I10245<= not (I10247 and I10248);
	I10246<= not (WX3587 and WX3247);
	I10247<= not (WX3587 and I10246);
	I10248<= not (WX3247 and I10246);
	I10253<= not (WX3311 and I10245);
	I10254<= not (WX3311 and I10253);
	I10255<= not (I10245 and I10253);
	I10260<= not (I10262 and I10263);
	I10261<= not (WX3375 and WX3439);
	I10262<= not (WX3375 and I10261);
	I10263<= not (WX3439 and I10261);
	I10268<= not (I10244 and I10260);
	I10269<= not (I10244 and I10268);
	I10270<= not (I10260 and I10268);
	I10275<= not (I10285 and I10286);
	I10276<= not (I10278 and I10279);
	I10277<= not (WX3587 and WX3249);
	I10278<= not (WX3587 and I10277);
	I10279<= not (WX3249 and I10277);
	I10284<= not (WX3313 and I10276);
	I10285<= not (WX3313 and I10284);
	I10286<= not (I10276 and I10284);
	I10291<= not (I10293 and I10294);
	I10292<= not (WX3377 and WX3441);
	I10293<= not (WX3377 and I10292);
	I10294<= not (WX3441 and I10292);
	I10299<= not (I10275 and I10291);
	I10300<= not (I10275 and I10299);
	I10301<= not (I10291 and I10299);
	I10306<= not (I10316 and I10317);
	I10307<= not (I10309 and I10310);
	I10308<= not (WX3587 and WX3251);
	I10309<= not (WX3587 and I10308);
	I10310<= not (WX3251 and I10308);
	I10315<= not (WX3315 and I10307);
	I10316<= not (WX3315 and I10315);
	I10317<= not (I10307 and I10315);
	I10322<= not (I10324 and I10325);
	I10323<= not (WX3379 and WX3443);
	I10324<= not (WX3379 and I10323);
	I10325<= not (WX3443 and I10323);
	I10330<= not (I10306 and I10322);
	I10331<= not (I10306 and I10330);
	I10332<= not (I10322 and I10330);
	I10337<= not (I10347 and I10348);
	I10338<= not (I10340 and I10341);
	I10339<= not (WX3587 and WX3253);
	I10340<= not (WX3587 and I10339);
	I10341<= not (WX3253 and I10339);
	I10346<= not (WX3317 and I10338);
	I10347<= not (WX3317 and I10346);
	I10348<= not (I10338 and I10346);
	I10353<= not (I10355 and I10356);
	I10354<= not (WX3381 and WX3445);
	I10355<= not (WX3381 and I10354);
	I10356<= not (WX3445 and I10354);
	I10361<= not (I10337 and I10353);
	I10362<= not (I10337 and I10361);
	I10363<= not (I10353 and I10361);
	I10368<= not (I10378 and I10379);
	I10369<= not (I10371 and I10372);
	I10370<= not (WX3587 and WX3255);
	I10371<= not (WX3587 and I10370);
	I10372<= not (WX3255 and I10370);
	I10377<= not (WX3319 and I10369);
	I10378<= not (WX3319 and I10377);
	I10379<= not (I10369 and I10377);
	I10384<= not (I10386 and I10387);
	I10385<= not (WX3383 and WX3447);
	I10386<= not (WX3383 and I10385);
	I10387<= not (WX3447 and I10385);
	I10392<= not (I10368 and I10384);
	I10393<= not (I10368 and I10392);
	I10394<= not (I10384 and I10392);
	I10399<= not (I10409 and I10410);
	I10400<= not (I10402 and I10403);
	I10401<= not (WX3587 and WX3257);
	I10402<= not (WX3587 and I10401);
	I10403<= not (WX3257 and I10401);
	I10408<= not (WX3321 and I10400);
	I10409<= not (WX3321 and I10408);
	I10410<= not (I10400 and I10408);
	I10415<= not (I10417 and I10418);
	I10416<= not (WX3385 and WX3449);
	I10417<= not (WX3385 and I10416);
	I10418<= not (WX3449 and I10416);
	I10423<= not (I10399 and I10415);
	I10424<= not (I10399 and I10423);
	I10425<= not (I10415 and I10423);
	I10430<= not (I10440 and I10441);
	I10431<= not (I10433 and I10434);
	I10432<= not (WX3587 and WX3259);
	I10433<= not (WX3587 and I10432);
	I10434<= not (WX3259 and I10432);
	I10439<= not (WX3323 and I10431);
	I10440<= not (WX3323 and I10439);
	I10441<= not (I10431 and I10439);
	I10446<= not (I10448 and I10449);
	I10447<= not (WX3387 and WX3451);
	I10448<= not (WX3387 and I10447);
	I10449<= not (WX3451 and I10447);
	I10454<= not (I10430 and I10446);
	I10455<= not (I10430 and I10454);
	I10456<= not (I10446 and I10454);
	I10461<= not (I10471 and I10472);
	I10462<= not (I10464 and I10465);
	I10463<= not (WX3587 and WX3261);
	I10464<= not (WX3587 and I10463);
	I10465<= not (WX3261 and I10463);
	I10470<= not (WX3325 and I10462);
	I10471<= not (WX3325 and I10470);
	I10472<= not (I10462 and I10470);
	I10477<= not (I10479 and I10480);
	I10478<= not (WX3389 and WX3453);
	I10479<= not (WX3389 and I10478);
	I10480<= not (WX3453 and I10478);
	I10485<= not (I10461 and I10477);
	I10486<= not (I10461 and I10485);
	I10487<= not (I10477 and I10485);
	I10492<= not (I10502 and I10503);
	I10493<= not (I10495 and I10496);
	I10494<= not (WX3588 and WX3263);
	I10495<= not (WX3588 and I10494);
	I10496<= not (WX3263 and I10494);
	I10501<= not (WX3327 and I10493);
	I10502<= not (WX3327 and I10501);
	I10503<= not (I10493 and I10501);
	I10508<= not (I10510 and I10511);
	I10509<= not (WX3391 and WX3455);
	I10510<= not (WX3391 and I10509);
	I10511<= not (WX3455 and I10509);
	I10516<= not (I10492 and I10508);
	I10517<= not (I10492 and I10516);
	I10518<= not (I10508 and I10516);
	I10523<= not (I10533 and I10534);
	I10524<= not (I10526 and I10527);
	I10525<= not (WX3588 and WX3265);
	I10526<= not (WX3588 and I10525);
	I10527<= not (WX3265 and I10525);
	I10532<= not (WX3329 and I10524);
	I10533<= not (WX3329 and I10532);
	I10534<= not (I10524 and I10532);
	I10539<= not (I10541 and I10542);
	I10540<= not (WX3393 and WX3457);
	I10541<= not (WX3393 and I10540);
	I10542<= not (WX3457 and I10540);
	I10547<= not (I10523 and I10539);
	I10548<= not (I10523 and I10547);
	I10549<= not (I10539 and I10547);
	I10554<= not (I10564 and I10565);
	I10555<= not (I10557 and I10558);
	I10556<= not (WX3588 and WX3267);
	I10557<= not (WX3588 and I10556);
	I10558<= not (WX3267 and I10556);
	I10563<= not (WX3331 and I10555);
	I10564<= not (WX3331 and I10563);
	I10565<= not (I10555 and I10563);
	I10570<= not (I10572 and I10573);
	I10571<= not (WX3395 and WX3459);
	I10572<= not (WX3395 and I10571);
	I10573<= not (WX3459 and I10571);
	I10578<= not (I10554 and I10570);
	I10579<= not (I10554 and I10578);
	I10580<= not (I10570 and I10578);
	I10585<= not (I10595 and I10596);
	I10586<= not (I10588 and I10589);
	I10587<= not (WX3588 and WX3269);
	I10588<= not (WX3588 and I10587);
	I10589<= not (WX3269 and I10587);
	I10594<= not (WX3333 and I10586);
	I10595<= not (WX3333 and I10594);
	I10596<= not (I10586 and I10594);
	I10601<= not (I10603 and I10604);
	I10602<= not (WX3397 and WX3461);
	I10603<= not (WX3397 and I10602);
	I10604<= not (WX3461 and I10602);
	I10609<= not (I10585 and I10601);
	I10610<= not (I10585 and I10609);
	I10611<= not (I10601 and I10609);
	I10616<= not (I10626 and I10627);
	I10617<= not (I10619 and I10620);
	I10618<= not (WX3588 and WX3271);
	I10619<= not (WX3588 and I10618);
	I10620<= not (WX3271 and I10618);
	I10625<= not (WX3335 and I10617);
	I10626<= not (WX3335 and I10625);
	I10627<= not (I10617 and I10625);
	I10632<= not (I10634 and I10635);
	I10633<= not (WX3399 and WX3463);
	I10634<= not (WX3399 and I10633);
	I10635<= not (WX3463 and I10633);
	I10640<= not (I10616 and I10632);
	I10641<= not (I10616 and I10640);
	I10642<= not (I10632 and I10640);
	I10647<= not (I10657 and I10658);
	I10648<= not (I10650 and I10651);
	I10649<= not (WX3588 and WX3273);
	I10650<= not (WX3588 and I10649);
	I10651<= not (WX3273 and I10649);
	I10656<= not (WX3337 and I10648);
	I10657<= not (WX3337 and I10656);
	I10658<= not (I10648 and I10656);
	I10663<= not (I10665 and I10666);
	I10664<= not (WX3401 and WX3465);
	I10665<= not (WX3401 and I10664);
	I10666<= not (WX3465 and I10664);
	I10671<= not (I10647 and I10663);
	I10672<= not (I10647 and I10671);
	I10673<= not (I10663 and I10671);
	I10678<= not (I10688 and I10689);
	I10679<= not (I10681 and I10682);
	I10680<= not (WX3588 and WX3275);
	I10681<= not (WX3588 and I10680);
	I10682<= not (WX3275 and I10680);
	I10687<= not (WX3339 and I10679);
	I10688<= not (WX3339 and I10687);
	I10689<= not (I10679 and I10687);
	I10694<= not (I10696 and I10697);
	I10695<= not (WX3403 and WX3467);
	I10696<= not (WX3403 and I10695);
	I10697<= not (WX3467 and I10695);
	I10702<= not (I10678 and I10694);
	I10703<= not (I10678 and I10702);
	I10704<= not (I10694 and I10702);
	I10709<= not (I10719 and I10720);
	I10710<= not (I10712 and I10713);
	I10711<= not (WX3588 and WX3277);
	I10712<= not (WX3588 and I10711);
	I10713<= not (WX3277 and I10711);
	I10718<= not (WX3341 and I10710);
	I10719<= not (WX3341 and I10718);
	I10720<= not (I10710 and I10718);
	I10725<= not (I10727 and I10728);
	I10726<= not (WX3405 and WX3469);
	I10727<= not (WX3405 and I10726);
	I10728<= not (WX3469 and I10726);
	I10733<= not (I10709 and I10725);
	I10734<= not (I10709 and I10733);
	I10735<= not (I10725 and I10733);
	I10740<= not (I10750 and I10751);
	I10741<= not (I10743 and I10744);
	I10742<= not (WX3588 and WX3279);
	I10743<= not (WX3588 and I10742);
	I10744<= not (WX3279 and I10742);
	I10749<= not (WX3343 and I10741);
	I10750<= not (WX3343 and I10749);
	I10751<= not (I10741 and I10749);
	I10756<= not (I10758 and I10759);
	I10757<= not (WX3407 and WX3471);
	I10758<= not (WX3407 and I10757);
	I10759<= not (WX3471 and I10757);
	I10764<= not (I10740 and I10756);
	I10765<= not (I10740 and I10764);
	I10766<= not (I10756 and I10764);
	I10771<= not (I10781 and I10782);
	I10772<= not (I10774 and I10775);
	I10773<= not (WX3588 and WX3281);
	I10774<= not (WX3588 and I10773);
	I10775<= not (WX3281 and I10773);
	I10780<= not (WX3345 and I10772);
	I10781<= not (WX3345 and I10780);
	I10782<= not (I10772 and I10780);
	I10787<= not (I10789 and I10790);
	I10788<= not (WX3409 and WX3473);
	I10789<= not (WX3409 and I10788);
	I10790<= not (WX3473 and I10788);
	I10795<= not (I10771 and I10787);
	I10796<= not (I10771 and I10795);
	I10797<= not (I10787 and I10795);
	I10802<= not (I10812 and I10813);
	I10803<= not (I10805 and I10806);
	I10804<= not (WX3588 and WX3283);
	I10805<= not (WX3588 and I10804);
	I10806<= not (WX3283 and I10804);
	I10811<= not (WX3347 and I10803);
	I10812<= not (WX3347 and I10811);
	I10813<= not (I10803 and I10811);
	I10818<= not (I10820 and I10821);
	I10819<= not (WX3411 and WX3475);
	I10820<= not (WX3411 and I10819);
	I10821<= not (WX3475 and I10819);
	I10826<= not (I10802 and I10818);
	I10827<= not (I10802 and I10826);
	I10828<= not (I10818 and I10826);
	I10833<= not (I10843 and I10844);
	I10834<= not (I10836 and I10837);
	I10835<= not (WX3588 and WX3285);
	I10836<= not (WX3588 and I10835);
	I10837<= not (WX3285 and I10835);
	I10842<= not (WX3349 and I10834);
	I10843<= not (WX3349 and I10842);
	I10844<= not (I10834 and I10842);
	I10849<= not (I10851 and I10852);
	I10850<= not (WX3413 and WX3477);
	I10851<= not (WX3413 and I10850);
	I10852<= not (WX3477 and I10850);
	I10857<= not (I10833 and I10849);
	I10858<= not (I10833 and I10857);
	I10859<= not (I10849 and I10857);
	I10864<= not (I10874 and I10875);
	I10865<= not (I10867 and I10868);
	I10866<= not (WX3588 and WX3287);
	I10867<= not (WX3588 and I10866);
	I10868<= not (WX3287 and I10866);
	I10873<= not (WX3351 and I10865);
	I10874<= not (WX3351 and I10873);
	I10875<= not (I10865 and I10873);
	I10880<= not (I10882 and I10883);
	I10881<= not (WX3415 and WX3479);
	I10882<= not (WX3415 and I10881);
	I10883<= not (WX3479 and I10881);
	I10888<= not (I10864 and I10880);
	I10889<= not (I10864 and I10888);
	I10890<= not (I10880 and I10888);
	I10895<= not (I10905 and I10906);
	I10896<= not (I10898 and I10899);
	I10897<= not (WX3588 and WX3289);
	I10898<= not (WX3588 and I10897);
	I10899<= not (WX3289 and I10897);
	I10904<= not (WX3353 and I10896);
	I10905<= not (WX3353 and I10904);
	I10906<= not (I10896 and I10904);
	I10911<= not (I10913 and I10914);
	I10912<= not (WX3417 and WX3481);
	I10913<= not (WX3417 and I10912);
	I10914<= not (WX3481 and I10912);
	I10919<= not (I10895 and I10911);
	I10920<= not (I10895 and I10919);
	I10921<= not (I10911 and I10919);
	I10926<= not (I10936 and I10937);
	I10927<= not (I10929 and I10930);
	I10928<= not (WX3588 and WX3291);
	I10929<= not (WX3588 and I10928);
	I10930<= not (WX3291 and I10928);
	I10935<= not (WX3355 and I10927);
	I10936<= not (WX3355 and I10935);
	I10937<= not (I10927 and I10935);
	I10942<= not (I10944 and I10945);
	I10943<= not (WX3419 and WX3483);
	I10944<= not (WX3419 and I10943);
	I10945<= not (WX3483 and I10943);
	I10950<= not (I10926 and I10942);
	I10951<= not (I10926 and I10950);
	I10952<= not (I10942 and I10950);
	I10957<= not (I10967 and I10968);
	I10958<= not (I10960 and I10961);
	I10959<= not (WX3588 and WX3293);
	I10960<= not (WX3588 and I10959);
	I10961<= not (WX3293 and I10959);
	I10966<= not (WX3357 and I10958);
	I10967<= not (WX3357 and I10966);
	I10968<= not (I10958 and I10966);
	I10973<= not (I10975 and I10976);
	I10974<= not (WX3421 and WX3485);
	I10975<= not (WX3421 and I10974);
	I10976<= not (WX3485 and I10974);
	I10981<= not (I10957 and I10973);
	I10982<= not (I10957 and I10981);
	I10983<= not (I10973 and I10981);
	I11062<= not (WX3166 and WX3071);
	I11063<= not (WX3166 and I11062);
	I11064<= not (WX3071 and I11062);
	I11075<= not (WX3167 and WX3073);
	I11076<= not (WX3167 and I11075);
	I11077<= not (WX3073 and I11075);
	I11088<= not (WX3168 and WX3075);
	I11089<= not (WX3168 and I11088);
	I11090<= not (WX3075 and I11088);
	I11101<= not (WX3169 and WX3077);
	I11102<= not (WX3169 and I11101);
	I11103<= not (WX3077 and I11101);
	I11114<= not (WX3170 and WX3079);
	I11115<= not (WX3170 and I11114);
	I11116<= not (WX3079 and I11114);
	I11127<= not (WX3171 and WX3081);
	I11128<= not (WX3171 and I11127);
	I11129<= not (WX3081 and I11127);
	I11140<= not (WX3172 and WX3083);
	I11141<= not (WX3172 and I11140);
	I11142<= not (WX3083 and I11140);
	I11153<= not (WX3173 and WX3085);
	I11154<= not (WX3173 and I11153);
	I11155<= not (WX3085 and I11153);
	I11166<= not (WX3174 and WX3087);
	I11167<= not (WX3174 and I11166);
	I11168<= not (WX3087 and I11166);
	I11179<= not (WX3175 and WX3089);
	I11180<= not (WX3175 and I11179);
	I11181<= not (WX3089 and I11179);
	I11192<= not (WX3176 and WX3091);
	I11193<= not (WX3176 and I11192);
	I11194<= not (WX3091 and I11192);
	I11205<= not (WX3177 and WX3093);
	I11206<= not (WX3177 and I11205);
	I11207<= not (WX3093 and I11205);
	I11218<= not (WX3178 and WX3095);
	I11219<= not (WX3178 and I11218);
	I11220<= not (WX3095 and I11218);
	I11231<= not (WX3179 and WX3097);
	I11232<= not (WX3179 and I11231);
	I11233<= not (WX3097 and I11231);
	I11244<= not (WX3180 and WX3099);
	I11245<= not (WX3180 and I11244);
	I11246<= not (WX3099 and I11244);
	I11257<= not (WX3181 and WX3101);
	I11258<= not (WX3181 and I11257);
	I11259<= not (WX3101 and I11257);
	I11270<= not (WX3182 and WX3103);
	I11271<= not (WX3182 and I11270);
	I11272<= not (WX3103 and I11270);
	I11283<= not (WX3183 and WX3105);
	I11284<= not (WX3183 and I11283);
	I11285<= not (WX3105 and I11283);
	I11296<= not (WX3184 and WX3107);
	I11297<= not (WX3184 and I11296);
	I11298<= not (WX3107 and I11296);
	I11309<= not (WX3185 and WX3109);
	I11310<= not (WX3185 and I11309);
	I11311<= not (WX3109 and I11309);
	I11322<= not (WX3186 and WX3111);
	I11323<= not (WX3186 and I11322);
	I11324<= not (WX3111 and I11322);
	I11335<= not (WX3187 and WX3113);
	I11336<= not (WX3187 and I11335);
	I11337<= not (WX3113 and I11335);
	I11348<= not (WX3188 and WX3115);
	I11349<= not (WX3188 and I11348);
	I11350<= not (WX3115 and I11348);
	I11361<= not (WX3189 and WX3117);
	I11362<= not (WX3189 and I11361);
	I11363<= not (WX3117 and I11361);
	I11374<= not (WX3190 and WX3119);
	I11375<= not (WX3190 and I11374);
	I11376<= not (WX3119 and I11374);
	I11387<= not (WX3191 and WX3121);
	I11388<= not (WX3191 and I11387);
	I11389<= not (WX3121 and I11387);
	I11400<= not (WX3192 and WX3123);
	I11401<= not (WX3192 and I11400);
	I11402<= not (WX3123 and I11400);
	I11413<= not (WX3193 and WX3125);
	I11414<= not (WX3193 and I11413);
	I11415<= not (WX3125 and I11413);
	I11426<= not (WX3194 and WX3127);
	I11427<= not (WX3194 and I11426);
	I11428<= not (WX3127 and I11426);
	I11439<= not (WX3195 and WX3129);
	I11440<= not (WX3195 and I11439);
	I11441<= not (WX3129 and I11439);
	I11452<= not (WX3196 and WX3131);
	I11453<= not (WX3196 and I11452);
	I11454<= not (WX3131 and I11452);
	I11465<= not (WX3197 and WX3133);
	I11466<= not (WX3197 and I11465);
	I11467<= not (WX3133 and I11465);
	I11479<= not (I11481 and I11482);
	I11480<= not (WX3213 and CRC_OUT_7_31);
	I11481<= not (WX3213 and I11480);
	I11482<= not (CRC_OUT_7_31 and I11480);
	I11487<= not (CRC_OUT_7_15 and I11479);
	I11488<= not (CRC_OUT_7_15 and I11487);
	I11489<= not (I11479 and I11487);
	I11494<= not (I11496 and I11497);
	I11495<= not (WX3218 and CRC_OUT_7_31);
	I11496<= not (WX3218 and I11495);
	I11497<= not (CRC_OUT_7_31 and I11495);
	I11502<= not (CRC_OUT_7_10 and I11494);
	I11503<= not (CRC_OUT_7_10 and I11502);
	I11504<= not (I11494 and I11502);
	I11509<= not (I11511 and I11512);
	I11510<= not (WX3225 and CRC_OUT_7_31);
	I11511<= not (WX3225 and I11510);
	I11512<= not (CRC_OUT_7_31 and I11510);
	I11517<= not (CRC_OUT_7_3 and I11509);
	I11518<= not (CRC_OUT_7_3 and I11517);
	I11519<= not (I11509 and I11517);
	I11524<= not (WX3229 and CRC_OUT_7_31);
	I11525<= not (WX3229 and I11524);
	I11526<= not (CRC_OUT_7_31 and I11524);
	I11531<= not (WX3198 and CRC_OUT_7_30);
	I11532<= not (WX3198 and I11531);
	I11533<= not (CRC_OUT_7_30 and I11531);
	I11538<= not (WX3199 and CRC_OUT_7_29);
	I11539<= not (WX3199 and I11538);
	I11540<= not (CRC_OUT_7_29 and I11538);
	I11545<= not (WX3200 and CRC_OUT_7_28);
	I11546<= not (WX3200 and I11545);
	I11547<= not (CRC_OUT_7_28 and I11545);
	I11552<= not (WX3201 and CRC_OUT_7_27);
	I11553<= not (WX3201 and I11552);
	I11554<= not (CRC_OUT_7_27 and I11552);
	I11559<= not (WX3202 and CRC_OUT_7_26);
	I11560<= not (WX3202 and I11559);
	I11561<= not (CRC_OUT_7_26 and I11559);
	I11566<= not (WX3203 and CRC_OUT_7_25);
	I11567<= not (WX3203 and I11566);
	I11568<= not (CRC_OUT_7_25 and I11566);
	I11573<= not (WX3204 and CRC_OUT_7_24);
	I11574<= not (WX3204 and I11573);
	I11575<= not (CRC_OUT_7_24 and I11573);
	I11580<= not (WX3205 and CRC_OUT_7_23);
	I11581<= not (WX3205 and I11580);
	I11582<= not (CRC_OUT_7_23 and I11580);
	I11587<= not (WX3206 and CRC_OUT_7_22);
	I11588<= not (WX3206 and I11587);
	I11589<= not (CRC_OUT_7_22 and I11587);
	I11594<= not (WX3207 and CRC_OUT_7_21);
	I11595<= not (WX3207 and I11594);
	I11596<= not (CRC_OUT_7_21 and I11594);
	I11601<= not (WX3208 and CRC_OUT_7_20);
	I11602<= not (WX3208 and I11601);
	I11603<= not (CRC_OUT_7_20 and I11601);
	I11608<= not (WX3209 and CRC_OUT_7_19);
	I11609<= not (WX3209 and I11608);
	I11610<= not (CRC_OUT_7_19 and I11608);
	I11615<= not (WX3210 and CRC_OUT_7_18);
	I11616<= not (WX3210 and I11615);
	I11617<= not (CRC_OUT_7_18 and I11615);
	I11622<= not (WX3211 and CRC_OUT_7_17);
	I11623<= not (WX3211 and I11622);
	I11624<= not (CRC_OUT_7_17 and I11622);
	I11629<= not (WX3212 and CRC_OUT_7_16);
	I11630<= not (WX3212 and I11629);
	I11631<= not (CRC_OUT_7_16 and I11629);
	I11636<= not (WX3214 and CRC_OUT_7_14);
	I11637<= not (WX3214 and I11636);
	I11638<= not (CRC_OUT_7_14 and I11636);
	I11643<= not (WX3215 and CRC_OUT_7_13);
	I11644<= not (WX3215 and I11643);
	I11645<= not (CRC_OUT_7_13 and I11643);
	I11650<= not (WX3216 and CRC_OUT_7_12);
	I11651<= not (WX3216 and I11650);
	I11652<= not (CRC_OUT_7_12 and I11650);
	I11657<= not (WX3217 and CRC_OUT_7_11);
	I11658<= not (WX3217 and I11657);
	I11659<= not (CRC_OUT_7_11 and I11657);
	I11664<= not (WX3219 and CRC_OUT_7_9);
	I11665<= not (WX3219 and I11664);
	I11666<= not (CRC_OUT_7_9 and I11664);
	I11671<= not (WX3220 and CRC_OUT_7_8);
	I11672<= not (WX3220 and I11671);
	I11673<= not (CRC_OUT_7_8 and I11671);
	I11678<= not (WX3221 and CRC_OUT_7_7);
	I11679<= not (WX3221 and I11678);
	I11680<= not (CRC_OUT_7_7 and I11678);
	I11685<= not (WX3222 and CRC_OUT_7_6);
	I11686<= not (WX3222 and I11685);
	I11687<= not (CRC_OUT_7_6 and I11685);
	I11692<= not (WX3223 and CRC_OUT_7_5);
	I11693<= not (WX3223 and I11692);
	I11694<= not (CRC_OUT_7_5 and I11692);
	I11699<= not (WX3224 and CRC_OUT_7_4);
	I11700<= not (WX3224 and I11699);
	I11701<= not (CRC_OUT_7_4 and I11699);
	I11706<= not (WX3226 and CRC_OUT_7_2);
	I11707<= not (WX3226 and I11706);
	I11708<= not (CRC_OUT_7_2 and I11706);
	I11713<= not (WX3227 and CRC_OUT_7_1);
	I11714<= not (WX3227 and I11713);
	I11715<= not (CRC_OUT_7_1 and I11713);
	I11720<= not (WX3228 and CRC_OUT_7_0);
	I11721<= not (WX3228 and I11720);
	I11722<= not (CRC_OUT_7_0 and I11720);
	I14001<= not (I14011 and I14012);
	I14002<= not (I14004 and I14005);
	I14003<= not (WX4880 and WX4524);
	I14004<= not (WX4880 and I14003);
	I14005<= not (WX4524 and I14003);
	I14010<= not (WX4588 and I14002);
	I14011<= not (WX4588 and I14010);
	I14012<= not (I14002 and I14010);
	I14017<= not (I14019 and I14020);
	I14018<= not (WX4652 and WX4716);
	I14019<= not (WX4652 and I14018);
	I14020<= not (WX4716 and I14018);
	I14025<= not (I14001 and I14017);
	I14026<= not (I14001 and I14025);
	I14027<= not (I14017 and I14025);
	I14032<= not (I14042 and I14043);
	I14033<= not (I14035 and I14036);
	I14034<= not (WX4880 and WX4526);
	I14035<= not (WX4880 and I14034);
	I14036<= not (WX4526 and I14034);
	I14041<= not (WX4590 and I14033);
	I14042<= not (WX4590 and I14041);
	I14043<= not (I14033 and I14041);
	I14048<= not (I14050 and I14051);
	I14049<= not (WX4654 and WX4718);
	I14050<= not (WX4654 and I14049);
	I14051<= not (WX4718 and I14049);
	I14056<= not (I14032 and I14048);
	I14057<= not (I14032 and I14056);
	I14058<= not (I14048 and I14056);
	I14063<= not (I14073 and I14074);
	I14064<= not (I14066 and I14067);
	I14065<= not (WX4880 and WX4528);
	I14066<= not (WX4880 and I14065);
	I14067<= not (WX4528 and I14065);
	I14072<= not (WX4592 and I14064);
	I14073<= not (WX4592 and I14072);
	I14074<= not (I14064 and I14072);
	I14079<= not (I14081 and I14082);
	I14080<= not (WX4656 and WX4720);
	I14081<= not (WX4656 and I14080);
	I14082<= not (WX4720 and I14080);
	I14087<= not (I14063 and I14079);
	I14088<= not (I14063 and I14087);
	I14089<= not (I14079 and I14087);
	I14094<= not (I14104 and I14105);
	I14095<= not (I14097 and I14098);
	I14096<= not (WX4880 and WX4530);
	I14097<= not (WX4880 and I14096);
	I14098<= not (WX4530 and I14096);
	I14103<= not (WX4594 and I14095);
	I14104<= not (WX4594 and I14103);
	I14105<= not (I14095 and I14103);
	I14110<= not (I14112 and I14113);
	I14111<= not (WX4658 and WX4722);
	I14112<= not (WX4658 and I14111);
	I14113<= not (WX4722 and I14111);
	I14118<= not (I14094 and I14110);
	I14119<= not (I14094 and I14118);
	I14120<= not (I14110 and I14118);
	I14125<= not (I14135 and I14136);
	I14126<= not (I14128 and I14129);
	I14127<= not (WX4880 and WX4532);
	I14128<= not (WX4880 and I14127);
	I14129<= not (WX4532 and I14127);
	I14134<= not (WX4596 and I14126);
	I14135<= not (WX4596 and I14134);
	I14136<= not (I14126 and I14134);
	I14141<= not (I14143 and I14144);
	I14142<= not (WX4660 and WX4724);
	I14143<= not (WX4660 and I14142);
	I14144<= not (WX4724 and I14142);
	I14149<= not (I14125 and I14141);
	I14150<= not (I14125 and I14149);
	I14151<= not (I14141 and I14149);
	I14156<= not (I14166 and I14167);
	I14157<= not (I14159 and I14160);
	I14158<= not (WX4880 and WX4534);
	I14159<= not (WX4880 and I14158);
	I14160<= not (WX4534 and I14158);
	I14165<= not (WX4598 and I14157);
	I14166<= not (WX4598 and I14165);
	I14167<= not (I14157 and I14165);
	I14172<= not (I14174 and I14175);
	I14173<= not (WX4662 and WX4726);
	I14174<= not (WX4662 and I14173);
	I14175<= not (WX4726 and I14173);
	I14180<= not (I14156 and I14172);
	I14181<= not (I14156 and I14180);
	I14182<= not (I14172 and I14180);
	I14187<= not (I14197 and I14198);
	I14188<= not (I14190 and I14191);
	I14189<= not (WX4880 and WX4536);
	I14190<= not (WX4880 and I14189);
	I14191<= not (WX4536 and I14189);
	I14196<= not (WX4600 and I14188);
	I14197<= not (WX4600 and I14196);
	I14198<= not (I14188 and I14196);
	I14203<= not (I14205 and I14206);
	I14204<= not (WX4664 and WX4728);
	I14205<= not (WX4664 and I14204);
	I14206<= not (WX4728 and I14204);
	I14211<= not (I14187 and I14203);
	I14212<= not (I14187 and I14211);
	I14213<= not (I14203 and I14211);
	I14218<= not (I14228 and I14229);
	I14219<= not (I14221 and I14222);
	I14220<= not (WX4880 and WX4538);
	I14221<= not (WX4880 and I14220);
	I14222<= not (WX4538 and I14220);
	I14227<= not (WX4602 and I14219);
	I14228<= not (WX4602 and I14227);
	I14229<= not (I14219 and I14227);
	I14234<= not (I14236 and I14237);
	I14235<= not (WX4666 and WX4730);
	I14236<= not (WX4666 and I14235);
	I14237<= not (WX4730 and I14235);
	I14242<= not (I14218 and I14234);
	I14243<= not (I14218 and I14242);
	I14244<= not (I14234 and I14242);
	I14249<= not (I14259 and I14260);
	I14250<= not (I14252 and I14253);
	I14251<= not (WX4880 and WX4540);
	I14252<= not (WX4880 and I14251);
	I14253<= not (WX4540 and I14251);
	I14258<= not (WX4604 and I14250);
	I14259<= not (WX4604 and I14258);
	I14260<= not (I14250 and I14258);
	I14265<= not (I14267 and I14268);
	I14266<= not (WX4668 and WX4732);
	I14267<= not (WX4668 and I14266);
	I14268<= not (WX4732 and I14266);
	I14273<= not (I14249 and I14265);
	I14274<= not (I14249 and I14273);
	I14275<= not (I14265 and I14273);
	I14280<= not (I14290 and I14291);
	I14281<= not (I14283 and I14284);
	I14282<= not (WX4880 and WX4542);
	I14283<= not (WX4880 and I14282);
	I14284<= not (WX4542 and I14282);
	I14289<= not (WX4606 and I14281);
	I14290<= not (WX4606 and I14289);
	I14291<= not (I14281 and I14289);
	I14296<= not (I14298 and I14299);
	I14297<= not (WX4670 and WX4734);
	I14298<= not (WX4670 and I14297);
	I14299<= not (WX4734 and I14297);
	I14304<= not (I14280 and I14296);
	I14305<= not (I14280 and I14304);
	I14306<= not (I14296 and I14304);
	I14311<= not (I14321 and I14322);
	I14312<= not (I14314 and I14315);
	I14313<= not (WX4880 and WX4544);
	I14314<= not (WX4880 and I14313);
	I14315<= not (WX4544 and I14313);
	I14320<= not (WX4608 and I14312);
	I14321<= not (WX4608 and I14320);
	I14322<= not (I14312 and I14320);
	I14327<= not (I14329 and I14330);
	I14328<= not (WX4672 and WX4736);
	I14329<= not (WX4672 and I14328);
	I14330<= not (WX4736 and I14328);
	I14335<= not (I14311 and I14327);
	I14336<= not (I14311 and I14335);
	I14337<= not (I14327 and I14335);
	I14342<= not (I14352 and I14353);
	I14343<= not (I14345 and I14346);
	I14344<= not (WX4880 and WX4546);
	I14345<= not (WX4880 and I14344);
	I14346<= not (WX4546 and I14344);
	I14351<= not (WX4610 and I14343);
	I14352<= not (WX4610 and I14351);
	I14353<= not (I14343 and I14351);
	I14358<= not (I14360 and I14361);
	I14359<= not (WX4674 and WX4738);
	I14360<= not (WX4674 and I14359);
	I14361<= not (WX4738 and I14359);
	I14366<= not (I14342 and I14358);
	I14367<= not (I14342 and I14366);
	I14368<= not (I14358 and I14366);
	I14373<= not (I14383 and I14384);
	I14374<= not (I14376 and I14377);
	I14375<= not (WX4880 and WX4548);
	I14376<= not (WX4880 and I14375);
	I14377<= not (WX4548 and I14375);
	I14382<= not (WX4612 and I14374);
	I14383<= not (WX4612 and I14382);
	I14384<= not (I14374 and I14382);
	I14389<= not (I14391 and I14392);
	I14390<= not (WX4676 and WX4740);
	I14391<= not (WX4676 and I14390);
	I14392<= not (WX4740 and I14390);
	I14397<= not (I14373 and I14389);
	I14398<= not (I14373 and I14397);
	I14399<= not (I14389 and I14397);
	I14404<= not (I14414 and I14415);
	I14405<= not (I14407 and I14408);
	I14406<= not (WX4880 and WX4550);
	I14407<= not (WX4880 and I14406);
	I14408<= not (WX4550 and I14406);
	I14413<= not (WX4614 and I14405);
	I14414<= not (WX4614 and I14413);
	I14415<= not (I14405 and I14413);
	I14420<= not (I14422 and I14423);
	I14421<= not (WX4678 and WX4742);
	I14422<= not (WX4678 and I14421);
	I14423<= not (WX4742 and I14421);
	I14428<= not (I14404 and I14420);
	I14429<= not (I14404 and I14428);
	I14430<= not (I14420 and I14428);
	I14435<= not (I14445 and I14446);
	I14436<= not (I14438 and I14439);
	I14437<= not (WX4880 and WX4552);
	I14438<= not (WX4880 and I14437);
	I14439<= not (WX4552 and I14437);
	I14444<= not (WX4616 and I14436);
	I14445<= not (WX4616 and I14444);
	I14446<= not (I14436 and I14444);
	I14451<= not (I14453 and I14454);
	I14452<= not (WX4680 and WX4744);
	I14453<= not (WX4680 and I14452);
	I14454<= not (WX4744 and I14452);
	I14459<= not (I14435 and I14451);
	I14460<= not (I14435 and I14459);
	I14461<= not (I14451 and I14459);
	I14466<= not (I14476 and I14477);
	I14467<= not (I14469 and I14470);
	I14468<= not (WX4880 and WX4554);
	I14469<= not (WX4880 and I14468);
	I14470<= not (WX4554 and I14468);
	I14475<= not (WX4618 and I14467);
	I14476<= not (WX4618 and I14475);
	I14477<= not (I14467 and I14475);
	I14482<= not (I14484 and I14485);
	I14483<= not (WX4682 and WX4746);
	I14484<= not (WX4682 and I14483);
	I14485<= not (WX4746 and I14483);
	I14490<= not (I14466 and I14482);
	I14491<= not (I14466 and I14490);
	I14492<= not (I14482 and I14490);
	I14497<= not (I14507 and I14508);
	I14498<= not (I14500 and I14501);
	I14499<= not (WX4881 and WX4556);
	I14500<= not (WX4881 and I14499);
	I14501<= not (WX4556 and I14499);
	I14506<= not (WX4620 and I14498);
	I14507<= not (WX4620 and I14506);
	I14508<= not (I14498 and I14506);
	I14513<= not (I14515 and I14516);
	I14514<= not (WX4684 and WX4748);
	I14515<= not (WX4684 and I14514);
	I14516<= not (WX4748 and I14514);
	I14521<= not (I14497 and I14513);
	I14522<= not (I14497 and I14521);
	I14523<= not (I14513 and I14521);
	I14528<= not (I14538 and I14539);
	I14529<= not (I14531 and I14532);
	I14530<= not (WX4881 and WX4558);
	I14531<= not (WX4881 and I14530);
	I14532<= not (WX4558 and I14530);
	I14537<= not (WX4622 and I14529);
	I14538<= not (WX4622 and I14537);
	I14539<= not (I14529 and I14537);
	I14544<= not (I14546 and I14547);
	I14545<= not (WX4686 and WX4750);
	I14546<= not (WX4686 and I14545);
	I14547<= not (WX4750 and I14545);
	I14552<= not (I14528 and I14544);
	I14553<= not (I14528 and I14552);
	I14554<= not (I14544 and I14552);
	I14559<= not (I14569 and I14570);
	I14560<= not (I14562 and I14563);
	I14561<= not (WX4881 and WX4560);
	I14562<= not (WX4881 and I14561);
	I14563<= not (WX4560 and I14561);
	I14568<= not (WX4624 and I14560);
	I14569<= not (WX4624 and I14568);
	I14570<= not (I14560 and I14568);
	I14575<= not (I14577 and I14578);
	I14576<= not (WX4688 and WX4752);
	I14577<= not (WX4688 and I14576);
	I14578<= not (WX4752 and I14576);
	I14583<= not (I14559 and I14575);
	I14584<= not (I14559 and I14583);
	I14585<= not (I14575 and I14583);
	I14590<= not (I14600 and I14601);
	I14591<= not (I14593 and I14594);
	I14592<= not (WX4881 and WX4562);
	I14593<= not (WX4881 and I14592);
	I14594<= not (WX4562 and I14592);
	I14599<= not (WX4626 and I14591);
	I14600<= not (WX4626 and I14599);
	I14601<= not (I14591 and I14599);
	I14606<= not (I14608 and I14609);
	I14607<= not (WX4690 and WX4754);
	I14608<= not (WX4690 and I14607);
	I14609<= not (WX4754 and I14607);
	I14614<= not (I14590 and I14606);
	I14615<= not (I14590 and I14614);
	I14616<= not (I14606 and I14614);
	I14621<= not (I14631 and I14632);
	I14622<= not (I14624 and I14625);
	I14623<= not (WX4881 and WX4564);
	I14624<= not (WX4881 and I14623);
	I14625<= not (WX4564 and I14623);
	I14630<= not (WX4628 and I14622);
	I14631<= not (WX4628 and I14630);
	I14632<= not (I14622 and I14630);
	I14637<= not (I14639 and I14640);
	I14638<= not (WX4692 and WX4756);
	I14639<= not (WX4692 and I14638);
	I14640<= not (WX4756 and I14638);
	I14645<= not (I14621 and I14637);
	I14646<= not (I14621 and I14645);
	I14647<= not (I14637 and I14645);
	I14652<= not (I14662 and I14663);
	I14653<= not (I14655 and I14656);
	I14654<= not (WX4881 and WX4566);
	I14655<= not (WX4881 and I14654);
	I14656<= not (WX4566 and I14654);
	I14661<= not (WX4630 and I14653);
	I14662<= not (WX4630 and I14661);
	I14663<= not (I14653 and I14661);
	I14668<= not (I14670 and I14671);
	I14669<= not (WX4694 and WX4758);
	I14670<= not (WX4694 and I14669);
	I14671<= not (WX4758 and I14669);
	I14676<= not (I14652 and I14668);
	I14677<= not (I14652 and I14676);
	I14678<= not (I14668 and I14676);
	I14683<= not (I14693 and I14694);
	I14684<= not (I14686 and I14687);
	I14685<= not (WX4881 and WX4568);
	I14686<= not (WX4881 and I14685);
	I14687<= not (WX4568 and I14685);
	I14692<= not (WX4632 and I14684);
	I14693<= not (WX4632 and I14692);
	I14694<= not (I14684 and I14692);
	I14699<= not (I14701 and I14702);
	I14700<= not (WX4696 and WX4760);
	I14701<= not (WX4696 and I14700);
	I14702<= not (WX4760 and I14700);
	I14707<= not (I14683 and I14699);
	I14708<= not (I14683 and I14707);
	I14709<= not (I14699 and I14707);
	I14714<= not (I14724 and I14725);
	I14715<= not (I14717 and I14718);
	I14716<= not (WX4881 and WX4570);
	I14717<= not (WX4881 and I14716);
	I14718<= not (WX4570 and I14716);
	I14723<= not (WX4634 and I14715);
	I14724<= not (WX4634 and I14723);
	I14725<= not (I14715 and I14723);
	I14730<= not (I14732 and I14733);
	I14731<= not (WX4698 and WX4762);
	I14732<= not (WX4698 and I14731);
	I14733<= not (WX4762 and I14731);
	I14738<= not (I14714 and I14730);
	I14739<= not (I14714 and I14738);
	I14740<= not (I14730 and I14738);
	I14745<= not (I14755 and I14756);
	I14746<= not (I14748 and I14749);
	I14747<= not (WX4881 and WX4572);
	I14748<= not (WX4881 and I14747);
	I14749<= not (WX4572 and I14747);
	I14754<= not (WX4636 and I14746);
	I14755<= not (WX4636 and I14754);
	I14756<= not (I14746 and I14754);
	I14761<= not (I14763 and I14764);
	I14762<= not (WX4700 and WX4764);
	I14763<= not (WX4700 and I14762);
	I14764<= not (WX4764 and I14762);
	I14769<= not (I14745 and I14761);
	I14770<= not (I14745 and I14769);
	I14771<= not (I14761 and I14769);
	I14776<= not (I14786 and I14787);
	I14777<= not (I14779 and I14780);
	I14778<= not (WX4881 and WX4574);
	I14779<= not (WX4881 and I14778);
	I14780<= not (WX4574 and I14778);
	I14785<= not (WX4638 and I14777);
	I14786<= not (WX4638 and I14785);
	I14787<= not (I14777 and I14785);
	I14792<= not (I14794 and I14795);
	I14793<= not (WX4702 and WX4766);
	I14794<= not (WX4702 and I14793);
	I14795<= not (WX4766 and I14793);
	I14800<= not (I14776 and I14792);
	I14801<= not (I14776 and I14800);
	I14802<= not (I14792 and I14800);
	I14807<= not (I14817 and I14818);
	I14808<= not (I14810 and I14811);
	I14809<= not (WX4881 and WX4576);
	I14810<= not (WX4881 and I14809);
	I14811<= not (WX4576 and I14809);
	I14816<= not (WX4640 and I14808);
	I14817<= not (WX4640 and I14816);
	I14818<= not (I14808 and I14816);
	I14823<= not (I14825 and I14826);
	I14824<= not (WX4704 and WX4768);
	I14825<= not (WX4704 and I14824);
	I14826<= not (WX4768 and I14824);
	I14831<= not (I14807 and I14823);
	I14832<= not (I14807 and I14831);
	I14833<= not (I14823 and I14831);
	I14838<= not (I14848 and I14849);
	I14839<= not (I14841 and I14842);
	I14840<= not (WX4881 and WX4578);
	I14841<= not (WX4881 and I14840);
	I14842<= not (WX4578 and I14840);
	I14847<= not (WX4642 and I14839);
	I14848<= not (WX4642 and I14847);
	I14849<= not (I14839 and I14847);
	I14854<= not (I14856 and I14857);
	I14855<= not (WX4706 and WX4770);
	I14856<= not (WX4706 and I14855);
	I14857<= not (WX4770 and I14855);
	I14862<= not (I14838 and I14854);
	I14863<= not (I14838 and I14862);
	I14864<= not (I14854 and I14862);
	I14869<= not (I14879 and I14880);
	I14870<= not (I14872 and I14873);
	I14871<= not (WX4881 and WX4580);
	I14872<= not (WX4881 and I14871);
	I14873<= not (WX4580 and I14871);
	I14878<= not (WX4644 and I14870);
	I14879<= not (WX4644 and I14878);
	I14880<= not (I14870 and I14878);
	I14885<= not (I14887 and I14888);
	I14886<= not (WX4708 and WX4772);
	I14887<= not (WX4708 and I14886);
	I14888<= not (WX4772 and I14886);
	I14893<= not (I14869 and I14885);
	I14894<= not (I14869 and I14893);
	I14895<= not (I14885 and I14893);
	I14900<= not (I14910 and I14911);
	I14901<= not (I14903 and I14904);
	I14902<= not (WX4881 and WX4582);
	I14903<= not (WX4881 and I14902);
	I14904<= not (WX4582 and I14902);
	I14909<= not (WX4646 and I14901);
	I14910<= not (WX4646 and I14909);
	I14911<= not (I14901 and I14909);
	I14916<= not (I14918 and I14919);
	I14917<= not (WX4710 and WX4774);
	I14918<= not (WX4710 and I14917);
	I14919<= not (WX4774 and I14917);
	I14924<= not (I14900 and I14916);
	I14925<= not (I14900 and I14924);
	I14926<= not (I14916 and I14924);
	I14931<= not (I14941 and I14942);
	I14932<= not (I14934 and I14935);
	I14933<= not (WX4881 and WX4584);
	I14934<= not (WX4881 and I14933);
	I14935<= not (WX4584 and I14933);
	I14940<= not (WX4648 and I14932);
	I14941<= not (WX4648 and I14940);
	I14942<= not (I14932 and I14940);
	I14947<= not (I14949 and I14950);
	I14948<= not (WX4712 and WX4776);
	I14949<= not (WX4712 and I14948);
	I14950<= not (WX4776 and I14948);
	I14955<= not (I14931 and I14947);
	I14956<= not (I14931 and I14955);
	I14957<= not (I14947 and I14955);
	I14962<= not (I14972 and I14973);
	I14963<= not (I14965 and I14966);
	I14964<= not (WX4881 and WX4586);
	I14965<= not (WX4881 and I14964);
	I14966<= not (WX4586 and I14964);
	I14971<= not (WX4650 and I14963);
	I14972<= not (WX4650 and I14971);
	I14973<= not (I14963 and I14971);
	I14978<= not (I14980 and I14981);
	I14979<= not (WX4714 and WX4778);
	I14980<= not (WX4714 and I14979);
	I14981<= not (WX4778 and I14979);
	I14986<= not (I14962 and I14978);
	I14987<= not (I14962 and I14986);
	I14988<= not (I14978 and I14986);
	I15067<= not (WX4459 and WX4364);
	I15068<= not (WX4459 and I15067);
	I15069<= not (WX4364 and I15067);
	I15080<= not (WX4460 and WX4366);
	I15081<= not (WX4460 and I15080);
	I15082<= not (WX4366 and I15080);
	I15093<= not (WX4461 and WX4368);
	I15094<= not (WX4461 and I15093);
	I15095<= not (WX4368 and I15093);
	I15106<= not (WX4462 and WX4370);
	I15107<= not (WX4462 and I15106);
	I15108<= not (WX4370 and I15106);
	I15119<= not (WX4463 and WX4372);
	I15120<= not (WX4463 and I15119);
	I15121<= not (WX4372 and I15119);
	I15132<= not (WX4464 and WX4374);
	I15133<= not (WX4464 and I15132);
	I15134<= not (WX4374 and I15132);
	I15145<= not (WX4465 and WX4376);
	I15146<= not (WX4465 and I15145);
	I15147<= not (WX4376 and I15145);
	I15158<= not (WX4466 and WX4378);
	I15159<= not (WX4466 and I15158);
	I15160<= not (WX4378 and I15158);
	I15171<= not (WX4467 and WX4380);
	I15172<= not (WX4467 and I15171);
	I15173<= not (WX4380 and I15171);
	I15184<= not (WX4468 and WX4382);
	I15185<= not (WX4468 and I15184);
	I15186<= not (WX4382 and I15184);
	I15197<= not (WX4469 and WX4384);
	I15198<= not (WX4469 and I15197);
	I15199<= not (WX4384 and I15197);
	I15210<= not (WX4470 and WX4386);
	I15211<= not (WX4470 and I15210);
	I15212<= not (WX4386 and I15210);
	I15223<= not (WX4471 and WX4388);
	I15224<= not (WX4471 and I15223);
	I15225<= not (WX4388 and I15223);
	I15236<= not (WX4472 and WX4390);
	I15237<= not (WX4472 and I15236);
	I15238<= not (WX4390 and I15236);
	I15249<= not (WX4473 and WX4392);
	I15250<= not (WX4473 and I15249);
	I15251<= not (WX4392 and I15249);
	I15262<= not (WX4474 and WX4394);
	I15263<= not (WX4474 and I15262);
	I15264<= not (WX4394 and I15262);
	I15275<= not (WX4475 and WX4396);
	I15276<= not (WX4475 and I15275);
	I15277<= not (WX4396 and I15275);
	I15288<= not (WX4476 and WX4398);
	I15289<= not (WX4476 and I15288);
	I15290<= not (WX4398 and I15288);
	I15301<= not (WX4477 and WX4400);
	I15302<= not (WX4477 and I15301);
	I15303<= not (WX4400 and I15301);
	I15314<= not (WX4478 and WX4402);
	I15315<= not (WX4478 and I15314);
	I15316<= not (WX4402 and I15314);
	I15327<= not (WX4479 and WX4404);
	I15328<= not (WX4479 and I15327);
	I15329<= not (WX4404 and I15327);
	I15340<= not (WX4480 and WX4406);
	I15341<= not (WX4480 and I15340);
	I15342<= not (WX4406 and I15340);
	I15353<= not (WX4481 and WX4408);
	I15354<= not (WX4481 and I15353);
	I15355<= not (WX4408 and I15353);
	I15366<= not (WX4482 and WX4410);
	I15367<= not (WX4482 and I15366);
	I15368<= not (WX4410 and I15366);
	I15379<= not (WX4483 and WX4412);
	I15380<= not (WX4483 and I15379);
	I15381<= not (WX4412 and I15379);
	I15392<= not (WX4484 and WX4414);
	I15393<= not (WX4484 and I15392);
	I15394<= not (WX4414 and I15392);
	I15405<= not (WX4485 and WX4416);
	I15406<= not (WX4485 and I15405);
	I15407<= not (WX4416 and I15405);
	I15418<= not (WX4486 and WX4418);
	I15419<= not (WX4486 and I15418);
	I15420<= not (WX4418 and I15418);
	I15431<= not (WX4487 and WX4420);
	I15432<= not (WX4487 and I15431);
	I15433<= not (WX4420 and I15431);
	I15444<= not (WX4488 and WX4422);
	I15445<= not (WX4488 and I15444);
	I15446<= not (WX4422 and I15444);
	I15457<= not (WX4489 and WX4424);
	I15458<= not (WX4489 and I15457);
	I15459<= not (WX4424 and I15457);
	I15470<= not (WX4490 and WX4426);
	I15471<= not (WX4490 and I15470);
	I15472<= not (WX4426 and I15470);
	I15484<= not (I15486 and I15487);
	I15485<= not (WX4506 and CRC_OUT_6_31);
	I15486<= not (WX4506 and I15485);
	I15487<= not (CRC_OUT_6_31 and I15485);
	I15492<= not (CRC_OUT_6_15 and I15484);
	I15493<= not (CRC_OUT_6_15 and I15492);
	I15494<= not (I15484 and I15492);
	I15499<= not (I15501 and I15502);
	I15500<= not (WX4511 and CRC_OUT_6_31);
	I15501<= not (WX4511 and I15500);
	I15502<= not (CRC_OUT_6_31 and I15500);
	I15507<= not (CRC_OUT_6_10 and I15499);
	I15508<= not (CRC_OUT_6_10 and I15507);
	I15509<= not (I15499 and I15507);
	I15514<= not (I15516 and I15517);
	I15515<= not (WX4518 and CRC_OUT_6_31);
	I15516<= not (WX4518 and I15515);
	I15517<= not (CRC_OUT_6_31 and I15515);
	I15522<= not (CRC_OUT_6_3 and I15514);
	I15523<= not (CRC_OUT_6_3 and I15522);
	I15524<= not (I15514 and I15522);
	I15529<= not (WX4522 and CRC_OUT_6_31);
	I15530<= not (WX4522 and I15529);
	I15531<= not (CRC_OUT_6_31 and I15529);
	I15536<= not (WX4491 and CRC_OUT_6_30);
	I15537<= not (WX4491 and I15536);
	I15538<= not (CRC_OUT_6_30 and I15536);
	I15543<= not (WX4492 and CRC_OUT_6_29);
	I15544<= not (WX4492 and I15543);
	I15545<= not (CRC_OUT_6_29 and I15543);
	I15550<= not (WX4493 and CRC_OUT_6_28);
	I15551<= not (WX4493 and I15550);
	I15552<= not (CRC_OUT_6_28 and I15550);
	I15557<= not (WX4494 and CRC_OUT_6_27);
	I15558<= not (WX4494 and I15557);
	I15559<= not (CRC_OUT_6_27 and I15557);
	I15564<= not (WX4495 and CRC_OUT_6_26);
	I15565<= not (WX4495 and I15564);
	I15566<= not (CRC_OUT_6_26 and I15564);
	I15571<= not (WX4496 and CRC_OUT_6_25);
	I15572<= not (WX4496 and I15571);
	I15573<= not (CRC_OUT_6_25 and I15571);
	I15578<= not (WX4497 and CRC_OUT_6_24);
	I15579<= not (WX4497 and I15578);
	I15580<= not (CRC_OUT_6_24 and I15578);
	I15585<= not (WX4498 and CRC_OUT_6_23);
	I15586<= not (WX4498 and I15585);
	I15587<= not (CRC_OUT_6_23 and I15585);
	I15592<= not (WX4499 and CRC_OUT_6_22);
	I15593<= not (WX4499 and I15592);
	I15594<= not (CRC_OUT_6_22 and I15592);
	I15599<= not (WX4500 and CRC_OUT_6_21);
	I15600<= not (WX4500 and I15599);
	I15601<= not (CRC_OUT_6_21 and I15599);
	I15606<= not (WX4501 and CRC_OUT_6_20);
	I15607<= not (WX4501 and I15606);
	I15608<= not (CRC_OUT_6_20 and I15606);
	I15613<= not (WX4502 and CRC_OUT_6_19);
	I15614<= not (WX4502 and I15613);
	I15615<= not (CRC_OUT_6_19 and I15613);
	I15620<= not (WX4503 and CRC_OUT_6_18);
	I15621<= not (WX4503 and I15620);
	I15622<= not (CRC_OUT_6_18 and I15620);
	I15627<= not (WX4504 and CRC_OUT_6_17);
	I15628<= not (WX4504 and I15627);
	I15629<= not (CRC_OUT_6_17 and I15627);
	I15634<= not (WX4505 and CRC_OUT_6_16);
	I15635<= not (WX4505 and I15634);
	I15636<= not (CRC_OUT_6_16 and I15634);
	I15641<= not (WX4507 and CRC_OUT_6_14);
	I15642<= not (WX4507 and I15641);
	I15643<= not (CRC_OUT_6_14 and I15641);
	I15648<= not (WX4508 and CRC_OUT_6_13);
	I15649<= not (WX4508 and I15648);
	I15650<= not (CRC_OUT_6_13 and I15648);
	I15655<= not (WX4509 and CRC_OUT_6_12);
	I15656<= not (WX4509 and I15655);
	I15657<= not (CRC_OUT_6_12 and I15655);
	I15662<= not (WX4510 and CRC_OUT_6_11);
	I15663<= not (WX4510 and I15662);
	I15664<= not (CRC_OUT_6_11 and I15662);
	I15669<= not (WX4512 and CRC_OUT_6_9);
	I15670<= not (WX4512 and I15669);
	I15671<= not (CRC_OUT_6_9 and I15669);
	I15676<= not (WX4513 and CRC_OUT_6_8);
	I15677<= not (WX4513 and I15676);
	I15678<= not (CRC_OUT_6_8 and I15676);
	I15683<= not (WX4514 and CRC_OUT_6_7);
	I15684<= not (WX4514 and I15683);
	I15685<= not (CRC_OUT_6_7 and I15683);
	I15690<= not (WX4515 and CRC_OUT_6_6);
	I15691<= not (WX4515 and I15690);
	I15692<= not (CRC_OUT_6_6 and I15690);
	I15697<= not (WX4516 and CRC_OUT_6_5);
	I15698<= not (WX4516 and I15697);
	I15699<= not (CRC_OUT_6_5 and I15697);
	I15704<= not (WX4517 and CRC_OUT_6_4);
	I15705<= not (WX4517 and I15704);
	I15706<= not (CRC_OUT_6_4 and I15704);
	I15711<= not (WX4519 and CRC_OUT_6_2);
	I15712<= not (WX4519 and I15711);
	I15713<= not (CRC_OUT_6_2 and I15711);
	I15718<= not (WX4520 and CRC_OUT_6_1);
	I15719<= not (WX4520 and I15718);
	I15720<= not (CRC_OUT_6_1 and I15718);
	I15725<= not (WX4521 and CRC_OUT_6_0);
	I15726<= not (WX4521 and I15725);
	I15727<= not (CRC_OUT_6_0 and I15725);
	I18006<= not (I18016 and I18017);
	I18007<= not (I18009 and I18010);
	I18008<= not (WX6173 and WX5817);
	I18009<= not (WX6173 and I18008);
	I18010<= not (WX5817 and I18008);
	I18015<= not (WX5881 and I18007);
	I18016<= not (WX5881 and I18015);
	I18017<= not (I18007 and I18015);
	I18022<= not (I18024 and I18025);
	I18023<= not (WX5945 and WX6009);
	I18024<= not (WX5945 and I18023);
	I18025<= not (WX6009 and I18023);
	I18030<= not (I18006 and I18022);
	I18031<= not (I18006 and I18030);
	I18032<= not (I18022 and I18030);
	I18037<= not (I18047 and I18048);
	I18038<= not (I18040 and I18041);
	I18039<= not (WX6173 and WX5819);
	I18040<= not (WX6173 and I18039);
	I18041<= not (WX5819 and I18039);
	I18046<= not (WX5883 and I18038);
	I18047<= not (WX5883 and I18046);
	I18048<= not (I18038 and I18046);
	I18053<= not (I18055 and I18056);
	I18054<= not (WX5947 and WX6011);
	I18055<= not (WX5947 and I18054);
	I18056<= not (WX6011 and I18054);
	I18061<= not (I18037 and I18053);
	I18062<= not (I18037 and I18061);
	I18063<= not (I18053 and I18061);
	I18068<= not (I18078 and I18079);
	I18069<= not (I18071 and I18072);
	I18070<= not (WX6173 and WX5821);
	I18071<= not (WX6173 and I18070);
	I18072<= not (WX5821 and I18070);
	I18077<= not (WX5885 and I18069);
	I18078<= not (WX5885 and I18077);
	I18079<= not (I18069 and I18077);
	I18084<= not (I18086 and I18087);
	I18085<= not (WX5949 and WX6013);
	I18086<= not (WX5949 and I18085);
	I18087<= not (WX6013 and I18085);
	I18092<= not (I18068 and I18084);
	I18093<= not (I18068 and I18092);
	I18094<= not (I18084 and I18092);
	I18099<= not (I18109 and I18110);
	I18100<= not (I18102 and I18103);
	I18101<= not (WX6173 and WX5823);
	I18102<= not (WX6173 and I18101);
	I18103<= not (WX5823 and I18101);
	I18108<= not (WX5887 and I18100);
	I18109<= not (WX5887 and I18108);
	I18110<= not (I18100 and I18108);
	I18115<= not (I18117 and I18118);
	I18116<= not (WX5951 and WX6015);
	I18117<= not (WX5951 and I18116);
	I18118<= not (WX6015 and I18116);
	I18123<= not (I18099 and I18115);
	I18124<= not (I18099 and I18123);
	I18125<= not (I18115 and I18123);
	I18130<= not (I18140 and I18141);
	I18131<= not (I18133 and I18134);
	I18132<= not (WX6173 and WX5825);
	I18133<= not (WX6173 and I18132);
	I18134<= not (WX5825 and I18132);
	I18139<= not (WX5889 and I18131);
	I18140<= not (WX5889 and I18139);
	I18141<= not (I18131 and I18139);
	I18146<= not (I18148 and I18149);
	I18147<= not (WX5953 and WX6017);
	I18148<= not (WX5953 and I18147);
	I18149<= not (WX6017 and I18147);
	I18154<= not (I18130 and I18146);
	I18155<= not (I18130 and I18154);
	I18156<= not (I18146 and I18154);
	I18161<= not (I18171 and I18172);
	I18162<= not (I18164 and I18165);
	I18163<= not (WX6173 and WX5827);
	I18164<= not (WX6173 and I18163);
	I18165<= not (WX5827 and I18163);
	I18170<= not (WX5891 and I18162);
	I18171<= not (WX5891 and I18170);
	I18172<= not (I18162 and I18170);
	I18177<= not (I18179 and I18180);
	I18178<= not (WX5955 and WX6019);
	I18179<= not (WX5955 and I18178);
	I18180<= not (WX6019 and I18178);
	I18185<= not (I18161 and I18177);
	I18186<= not (I18161 and I18185);
	I18187<= not (I18177 and I18185);
	I18192<= not (I18202 and I18203);
	I18193<= not (I18195 and I18196);
	I18194<= not (WX6173 and WX5829);
	I18195<= not (WX6173 and I18194);
	I18196<= not (WX5829 and I18194);
	I18201<= not (WX5893 and I18193);
	I18202<= not (WX5893 and I18201);
	I18203<= not (I18193 and I18201);
	I18208<= not (I18210 and I18211);
	I18209<= not (WX5957 and WX6021);
	I18210<= not (WX5957 and I18209);
	I18211<= not (WX6021 and I18209);
	I18216<= not (I18192 and I18208);
	I18217<= not (I18192 and I18216);
	I18218<= not (I18208 and I18216);
	I18223<= not (I18233 and I18234);
	I18224<= not (I18226 and I18227);
	I18225<= not (WX6173 and WX5831);
	I18226<= not (WX6173 and I18225);
	I18227<= not (WX5831 and I18225);
	I18232<= not (WX5895 and I18224);
	I18233<= not (WX5895 and I18232);
	I18234<= not (I18224 and I18232);
	I18239<= not (I18241 and I18242);
	I18240<= not (WX5959 and WX6023);
	I18241<= not (WX5959 and I18240);
	I18242<= not (WX6023 and I18240);
	I18247<= not (I18223 and I18239);
	I18248<= not (I18223 and I18247);
	I18249<= not (I18239 and I18247);
	I18254<= not (I18264 and I18265);
	I18255<= not (I18257 and I18258);
	I18256<= not (WX6173 and WX5833);
	I18257<= not (WX6173 and I18256);
	I18258<= not (WX5833 and I18256);
	I18263<= not (WX5897 and I18255);
	I18264<= not (WX5897 and I18263);
	I18265<= not (I18255 and I18263);
	I18270<= not (I18272 and I18273);
	I18271<= not (WX5961 and WX6025);
	I18272<= not (WX5961 and I18271);
	I18273<= not (WX6025 and I18271);
	I18278<= not (I18254 and I18270);
	I18279<= not (I18254 and I18278);
	I18280<= not (I18270 and I18278);
	I18285<= not (I18295 and I18296);
	I18286<= not (I18288 and I18289);
	I18287<= not (WX6173 and WX5835);
	I18288<= not (WX6173 and I18287);
	I18289<= not (WX5835 and I18287);
	I18294<= not (WX5899 and I18286);
	I18295<= not (WX5899 and I18294);
	I18296<= not (I18286 and I18294);
	I18301<= not (I18303 and I18304);
	I18302<= not (WX5963 and WX6027);
	I18303<= not (WX5963 and I18302);
	I18304<= not (WX6027 and I18302);
	I18309<= not (I18285 and I18301);
	I18310<= not (I18285 and I18309);
	I18311<= not (I18301 and I18309);
	I18316<= not (I18326 and I18327);
	I18317<= not (I18319 and I18320);
	I18318<= not (WX6173 and WX5837);
	I18319<= not (WX6173 and I18318);
	I18320<= not (WX5837 and I18318);
	I18325<= not (WX5901 and I18317);
	I18326<= not (WX5901 and I18325);
	I18327<= not (I18317 and I18325);
	I18332<= not (I18334 and I18335);
	I18333<= not (WX5965 and WX6029);
	I18334<= not (WX5965 and I18333);
	I18335<= not (WX6029 and I18333);
	I18340<= not (I18316 and I18332);
	I18341<= not (I18316 and I18340);
	I18342<= not (I18332 and I18340);
	I18347<= not (I18357 and I18358);
	I18348<= not (I18350 and I18351);
	I18349<= not (WX6173 and WX5839);
	I18350<= not (WX6173 and I18349);
	I18351<= not (WX5839 and I18349);
	I18356<= not (WX5903 and I18348);
	I18357<= not (WX5903 and I18356);
	I18358<= not (I18348 and I18356);
	I18363<= not (I18365 and I18366);
	I18364<= not (WX5967 and WX6031);
	I18365<= not (WX5967 and I18364);
	I18366<= not (WX6031 and I18364);
	I18371<= not (I18347 and I18363);
	I18372<= not (I18347 and I18371);
	I18373<= not (I18363 and I18371);
	I18378<= not (I18388 and I18389);
	I18379<= not (I18381 and I18382);
	I18380<= not (WX6173 and WX5841);
	I18381<= not (WX6173 and I18380);
	I18382<= not (WX5841 and I18380);
	I18387<= not (WX5905 and I18379);
	I18388<= not (WX5905 and I18387);
	I18389<= not (I18379 and I18387);
	I18394<= not (I18396 and I18397);
	I18395<= not (WX5969 and WX6033);
	I18396<= not (WX5969 and I18395);
	I18397<= not (WX6033 and I18395);
	I18402<= not (I18378 and I18394);
	I18403<= not (I18378 and I18402);
	I18404<= not (I18394 and I18402);
	I18409<= not (I18419 and I18420);
	I18410<= not (I18412 and I18413);
	I18411<= not (WX6173 and WX5843);
	I18412<= not (WX6173 and I18411);
	I18413<= not (WX5843 and I18411);
	I18418<= not (WX5907 and I18410);
	I18419<= not (WX5907 and I18418);
	I18420<= not (I18410 and I18418);
	I18425<= not (I18427 and I18428);
	I18426<= not (WX5971 and WX6035);
	I18427<= not (WX5971 and I18426);
	I18428<= not (WX6035 and I18426);
	I18433<= not (I18409 and I18425);
	I18434<= not (I18409 and I18433);
	I18435<= not (I18425 and I18433);
	I18440<= not (I18450 and I18451);
	I18441<= not (I18443 and I18444);
	I18442<= not (WX6173 and WX5845);
	I18443<= not (WX6173 and I18442);
	I18444<= not (WX5845 and I18442);
	I18449<= not (WX5909 and I18441);
	I18450<= not (WX5909 and I18449);
	I18451<= not (I18441 and I18449);
	I18456<= not (I18458 and I18459);
	I18457<= not (WX5973 and WX6037);
	I18458<= not (WX5973 and I18457);
	I18459<= not (WX6037 and I18457);
	I18464<= not (I18440 and I18456);
	I18465<= not (I18440 and I18464);
	I18466<= not (I18456 and I18464);
	I18471<= not (I18481 and I18482);
	I18472<= not (I18474 and I18475);
	I18473<= not (WX6173 and WX5847);
	I18474<= not (WX6173 and I18473);
	I18475<= not (WX5847 and I18473);
	I18480<= not (WX5911 and I18472);
	I18481<= not (WX5911 and I18480);
	I18482<= not (I18472 and I18480);
	I18487<= not (I18489 and I18490);
	I18488<= not (WX5975 and WX6039);
	I18489<= not (WX5975 and I18488);
	I18490<= not (WX6039 and I18488);
	I18495<= not (I18471 and I18487);
	I18496<= not (I18471 and I18495);
	I18497<= not (I18487 and I18495);
	I18502<= not (I18512 and I18513);
	I18503<= not (I18505 and I18506);
	I18504<= not (WX6174 and WX5849);
	I18505<= not (WX6174 and I18504);
	I18506<= not (WX5849 and I18504);
	I18511<= not (WX5913 and I18503);
	I18512<= not (WX5913 and I18511);
	I18513<= not (I18503 and I18511);
	I18518<= not (I18520 and I18521);
	I18519<= not (WX5977 and WX6041);
	I18520<= not (WX5977 and I18519);
	I18521<= not (WX6041 and I18519);
	I18526<= not (I18502 and I18518);
	I18527<= not (I18502 and I18526);
	I18528<= not (I18518 and I18526);
	I18533<= not (I18543 and I18544);
	I18534<= not (I18536 and I18537);
	I18535<= not (WX6174 and WX5851);
	I18536<= not (WX6174 and I18535);
	I18537<= not (WX5851 and I18535);
	I18542<= not (WX5915 and I18534);
	I18543<= not (WX5915 and I18542);
	I18544<= not (I18534 and I18542);
	I18549<= not (I18551 and I18552);
	I18550<= not (WX5979 and WX6043);
	I18551<= not (WX5979 and I18550);
	I18552<= not (WX6043 and I18550);
	I18557<= not (I18533 and I18549);
	I18558<= not (I18533 and I18557);
	I18559<= not (I18549 and I18557);
	I18564<= not (I18574 and I18575);
	I18565<= not (I18567 and I18568);
	I18566<= not (WX6174 and WX5853);
	I18567<= not (WX6174 and I18566);
	I18568<= not (WX5853 and I18566);
	I18573<= not (WX5917 and I18565);
	I18574<= not (WX5917 and I18573);
	I18575<= not (I18565 and I18573);
	I18580<= not (I18582 and I18583);
	I18581<= not (WX5981 and WX6045);
	I18582<= not (WX5981 and I18581);
	I18583<= not (WX6045 and I18581);
	I18588<= not (I18564 and I18580);
	I18589<= not (I18564 and I18588);
	I18590<= not (I18580 and I18588);
	I18595<= not (I18605 and I18606);
	I18596<= not (I18598 and I18599);
	I18597<= not (WX6174 and WX5855);
	I18598<= not (WX6174 and I18597);
	I18599<= not (WX5855 and I18597);
	I18604<= not (WX5919 and I18596);
	I18605<= not (WX5919 and I18604);
	I18606<= not (I18596 and I18604);
	I18611<= not (I18613 and I18614);
	I18612<= not (WX5983 and WX6047);
	I18613<= not (WX5983 and I18612);
	I18614<= not (WX6047 and I18612);
	I18619<= not (I18595 and I18611);
	I18620<= not (I18595 and I18619);
	I18621<= not (I18611 and I18619);
	I18626<= not (I18636 and I18637);
	I18627<= not (I18629 and I18630);
	I18628<= not (WX6174 and WX5857);
	I18629<= not (WX6174 and I18628);
	I18630<= not (WX5857 and I18628);
	I18635<= not (WX5921 and I18627);
	I18636<= not (WX5921 and I18635);
	I18637<= not (I18627 and I18635);
	I18642<= not (I18644 and I18645);
	I18643<= not (WX5985 and WX6049);
	I18644<= not (WX5985 and I18643);
	I18645<= not (WX6049 and I18643);
	I18650<= not (I18626 and I18642);
	I18651<= not (I18626 and I18650);
	I18652<= not (I18642 and I18650);
	I18657<= not (I18667 and I18668);
	I18658<= not (I18660 and I18661);
	I18659<= not (WX6174 and WX5859);
	I18660<= not (WX6174 and I18659);
	I18661<= not (WX5859 and I18659);
	I18666<= not (WX5923 and I18658);
	I18667<= not (WX5923 and I18666);
	I18668<= not (I18658 and I18666);
	I18673<= not (I18675 and I18676);
	I18674<= not (WX5987 and WX6051);
	I18675<= not (WX5987 and I18674);
	I18676<= not (WX6051 and I18674);
	I18681<= not (I18657 and I18673);
	I18682<= not (I18657 and I18681);
	I18683<= not (I18673 and I18681);
	I18688<= not (I18698 and I18699);
	I18689<= not (I18691 and I18692);
	I18690<= not (WX6174 and WX5861);
	I18691<= not (WX6174 and I18690);
	I18692<= not (WX5861 and I18690);
	I18697<= not (WX5925 and I18689);
	I18698<= not (WX5925 and I18697);
	I18699<= not (I18689 and I18697);
	I18704<= not (I18706 and I18707);
	I18705<= not (WX5989 and WX6053);
	I18706<= not (WX5989 and I18705);
	I18707<= not (WX6053 and I18705);
	I18712<= not (I18688 and I18704);
	I18713<= not (I18688 and I18712);
	I18714<= not (I18704 and I18712);
	I18719<= not (I18729 and I18730);
	I18720<= not (I18722 and I18723);
	I18721<= not (WX6174 and WX5863);
	I18722<= not (WX6174 and I18721);
	I18723<= not (WX5863 and I18721);
	I18728<= not (WX5927 and I18720);
	I18729<= not (WX5927 and I18728);
	I18730<= not (I18720 and I18728);
	I18735<= not (I18737 and I18738);
	I18736<= not (WX5991 and WX6055);
	I18737<= not (WX5991 and I18736);
	I18738<= not (WX6055 and I18736);
	I18743<= not (I18719 and I18735);
	I18744<= not (I18719 and I18743);
	I18745<= not (I18735 and I18743);
	I18750<= not (I18760 and I18761);
	I18751<= not (I18753 and I18754);
	I18752<= not (WX6174 and WX5865);
	I18753<= not (WX6174 and I18752);
	I18754<= not (WX5865 and I18752);
	I18759<= not (WX5929 and I18751);
	I18760<= not (WX5929 and I18759);
	I18761<= not (I18751 and I18759);
	I18766<= not (I18768 and I18769);
	I18767<= not (WX5993 and WX6057);
	I18768<= not (WX5993 and I18767);
	I18769<= not (WX6057 and I18767);
	I18774<= not (I18750 and I18766);
	I18775<= not (I18750 and I18774);
	I18776<= not (I18766 and I18774);
	I18781<= not (I18791 and I18792);
	I18782<= not (I18784 and I18785);
	I18783<= not (WX6174 and WX5867);
	I18784<= not (WX6174 and I18783);
	I18785<= not (WX5867 and I18783);
	I18790<= not (WX5931 and I18782);
	I18791<= not (WX5931 and I18790);
	I18792<= not (I18782 and I18790);
	I18797<= not (I18799 and I18800);
	I18798<= not (WX5995 and WX6059);
	I18799<= not (WX5995 and I18798);
	I18800<= not (WX6059 and I18798);
	I18805<= not (I18781 and I18797);
	I18806<= not (I18781 and I18805);
	I18807<= not (I18797 and I18805);
	I18812<= not (I18822 and I18823);
	I18813<= not (I18815 and I18816);
	I18814<= not (WX6174 and WX5869);
	I18815<= not (WX6174 and I18814);
	I18816<= not (WX5869 and I18814);
	I18821<= not (WX5933 and I18813);
	I18822<= not (WX5933 and I18821);
	I18823<= not (I18813 and I18821);
	I18828<= not (I18830 and I18831);
	I18829<= not (WX5997 and WX6061);
	I18830<= not (WX5997 and I18829);
	I18831<= not (WX6061 and I18829);
	I18836<= not (I18812 and I18828);
	I18837<= not (I18812 and I18836);
	I18838<= not (I18828 and I18836);
	I18843<= not (I18853 and I18854);
	I18844<= not (I18846 and I18847);
	I18845<= not (WX6174 and WX5871);
	I18846<= not (WX6174 and I18845);
	I18847<= not (WX5871 and I18845);
	I18852<= not (WX5935 and I18844);
	I18853<= not (WX5935 and I18852);
	I18854<= not (I18844 and I18852);
	I18859<= not (I18861 and I18862);
	I18860<= not (WX5999 and WX6063);
	I18861<= not (WX5999 and I18860);
	I18862<= not (WX6063 and I18860);
	I18867<= not (I18843 and I18859);
	I18868<= not (I18843 and I18867);
	I18869<= not (I18859 and I18867);
	I18874<= not (I18884 and I18885);
	I18875<= not (I18877 and I18878);
	I18876<= not (WX6174 and WX5873);
	I18877<= not (WX6174 and I18876);
	I18878<= not (WX5873 and I18876);
	I18883<= not (WX5937 and I18875);
	I18884<= not (WX5937 and I18883);
	I18885<= not (I18875 and I18883);
	I18890<= not (I18892 and I18893);
	I18891<= not (WX6001 and WX6065);
	I18892<= not (WX6001 and I18891);
	I18893<= not (WX6065 and I18891);
	I18898<= not (I18874 and I18890);
	I18899<= not (I18874 and I18898);
	I18900<= not (I18890 and I18898);
	I18905<= not (I18915 and I18916);
	I18906<= not (I18908 and I18909);
	I18907<= not (WX6174 and WX5875);
	I18908<= not (WX6174 and I18907);
	I18909<= not (WX5875 and I18907);
	I18914<= not (WX5939 and I18906);
	I18915<= not (WX5939 and I18914);
	I18916<= not (I18906 and I18914);
	I18921<= not (I18923 and I18924);
	I18922<= not (WX6003 and WX6067);
	I18923<= not (WX6003 and I18922);
	I18924<= not (WX6067 and I18922);
	I18929<= not (I18905 and I18921);
	I18930<= not (I18905 and I18929);
	I18931<= not (I18921 and I18929);
	I18936<= not (I18946 and I18947);
	I18937<= not (I18939 and I18940);
	I18938<= not (WX6174 and WX5877);
	I18939<= not (WX6174 and I18938);
	I18940<= not (WX5877 and I18938);
	I18945<= not (WX5941 and I18937);
	I18946<= not (WX5941 and I18945);
	I18947<= not (I18937 and I18945);
	I18952<= not (I18954 and I18955);
	I18953<= not (WX6005 and WX6069);
	I18954<= not (WX6005 and I18953);
	I18955<= not (WX6069 and I18953);
	I18960<= not (I18936 and I18952);
	I18961<= not (I18936 and I18960);
	I18962<= not (I18952 and I18960);
	I18967<= not (I18977 and I18978);
	I18968<= not (I18970 and I18971);
	I18969<= not (WX6174 and WX5879);
	I18970<= not (WX6174 and I18969);
	I18971<= not (WX5879 and I18969);
	I18976<= not (WX5943 and I18968);
	I18977<= not (WX5943 and I18976);
	I18978<= not (I18968 and I18976);
	I18983<= not (I18985 and I18986);
	I18984<= not (WX6007 and WX6071);
	I18985<= not (WX6007 and I18984);
	I18986<= not (WX6071 and I18984);
	I18991<= not (I18967 and I18983);
	I18992<= not (I18967 and I18991);
	I18993<= not (I18983 and I18991);
	I19072<= not (WX5752 and WX5657);
	I19073<= not (WX5752 and I19072);
	I19074<= not (WX5657 and I19072);
	I19085<= not (WX5753 and WX5659);
	I19086<= not (WX5753 and I19085);
	I19087<= not (WX5659 and I19085);
	I19098<= not (WX5754 and WX5661);
	I19099<= not (WX5754 and I19098);
	I19100<= not (WX5661 and I19098);
	I19111<= not (WX5755 and WX5663);
	I19112<= not (WX5755 and I19111);
	I19113<= not (WX5663 and I19111);
	I19124<= not (WX5756 and WX5665);
	I19125<= not (WX5756 and I19124);
	I19126<= not (WX5665 and I19124);
	I19137<= not (WX5757 and WX5667);
	I19138<= not (WX5757 and I19137);
	I19139<= not (WX5667 and I19137);
	I19150<= not (WX5758 and WX5669);
	I19151<= not (WX5758 and I19150);
	I19152<= not (WX5669 and I19150);
	I19163<= not (WX5759 and WX5671);
	I19164<= not (WX5759 and I19163);
	I19165<= not (WX5671 and I19163);
	I19176<= not (WX5760 and WX5673);
	I19177<= not (WX5760 and I19176);
	I19178<= not (WX5673 and I19176);
	I19189<= not (WX5761 and WX5675);
	I19190<= not (WX5761 and I19189);
	I19191<= not (WX5675 and I19189);
	I19202<= not (WX5762 and WX5677);
	I19203<= not (WX5762 and I19202);
	I19204<= not (WX5677 and I19202);
	I19215<= not (WX5763 and WX5679);
	I19216<= not (WX5763 and I19215);
	I19217<= not (WX5679 and I19215);
	I19228<= not (WX5764 and WX5681);
	I19229<= not (WX5764 and I19228);
	I19230<= not (WX5681 and I19228);
	I19241<= not (WX5765 and WX5683);
	I19242<= not (WX5765 and I19241);
	I19243<= not (WX5683 and I19241);
	I19254<= not (WX5766 and WX5685);
	I19255<= not (WX5766 and I19254);
	I19256<= not (WX5685 and I19254);
	I19267<= not (WX5767 and WX5687);
	I19268<= not (WX5767 and I19267);
	I19269<= not (WX5687 and I19267);
	I19280<= not (WX5768 and WX5689);
	I19281<= not (WX5768 and I19280);
	I19282<= not (WX5689 and I19280);
	I19293<= not (WX5769 and WX5691);
	I19294<= not (WX5769 and I19293);
	I19295<= not (WX5691 and I19293);
	I19306<= not (WX5770 and WX5693);
	I19307<= not (WX5770 and I19306);
	I19308<= not (WX5693 and I19306);
	I19319<= not (WX5771 and WX5695);
	I19320<= not (WX5771 and I19319);
	I19321<= not (WX5695 and I19319);
	I19332<= not (WX5772 and WX5697);
	I19333<= not (WX5772 and I19332);
	I19334<= not (WX5697 and I19332);
	I19345<= not (WX5773 and WX5699);
	I19346<= not (WX5773 and I19345);
	I19347<= not (WX5699 and I19345);
	I19358<= not (WX5774 and WX5701);
	I19359<= not (WX5774 and I19358);
	I19360<= not (WX5701 and I19358);
	I19371<= not (WX5775 and WX5703);
	I19372<= not (WX5775 and I19371);
	I19373<= not (WX5703 and I19371);
	I19384<= not (WX5776 and WX5705);
	I19385<= not (WX5776 and I19384);
	I19386<= not (WX5705 and I19384);
	I19397<= not (WX5777 and WX5707);
	I19398<= not (WX5777 and I19397);
	I19399<= not (WX5707 and I19397);
	I19410<= not (WX5778 and WX5709);
	I19411<= not (WX5778 and I19410);
	I19412<= not (WX5709 and I19410);
	I19423<= not (WX5779 and WX5711);
	I19424<= not (WX5779 and I19423);
	I19425<= not (WX5711 and I19423);
	I19436<= not (WX5780 and WX5713);
	I19437<= not (WX5780 and I19436);
	I19438<= not (WX5713 and I19436);
	I19449<= not (WX5781 and WX5715);
	I19450<= not (WX5781 and I19449);
	I19451<= not (WX5715 and I19449);
	I19462<= not (WX5782 and WX5717);
	I19463<= not (WX5782 and I19462);
	I19464<= not (WX5717 and I19462);
	I19475<= not (WX5783 and WX5719);
	I19476<= not (WX5783 and I19475);
	I19477<= not (WX5719 and I19475);
	I19489<= not (I19491 and I19492);
	I19490<= not (WX5799 and CRC_OUT_5_31);
	I19491<= not (WX5799 and I19490);
	I19492<= not (CRC_OUT_5_31 and I19490);
	I19497<= not (CRC_OUT_5_15 and I19489);
	I19498<= not (CRC_OUT_5_15 and I19497);
	I19499<= not (I19489 and I19497);
	I19504<= not (I19506 and I19507);
	I19505<= not (WX5804 and CRC_OUT_5_31);
	I19506<= not (WX5804 and I19505);
	I19507<= not (CRC_OUT_5_31 and I19505);
	I19512<= not (CRC_OUT_5_10 and I19504);
	I19513<= not (CRC_OUT_5_10 and I19512);
	I19514<= not (I19504 and I19512);
	I19519<= not (I19521 and I19522);
	I19520<= not (WX5811 and CRC_OUT_5_31);
	I19521<= not (WX5811 and I19520);
	I19522<= not (CRC_OUT_5_31 and I19520);
	I19527<= not (CRC_OUT_5_3 and I19519);
	I19528<= not (CRC_OUT_5_3 and I19527);
	I19529<= not (I19519 and I19527);
	I19534<= not (WX5815 and CRC_OUT_5_31);
	I19535<= not (WX5815 and I19534);
	I19536<= not (CRC_OUT_5_31 and I19534);
	I19541<= not (WX5784 and CRC_OUT_5_30);
	I19542<= not (WX5784 and I19541);
	I19543<= not (CRC_OUT_5_30 and I19541);
	I19548<= not (WX5785 and CRC_OUT_5_29);
	I19549<= not (WX5785 and I19548);
	I19550<= not (CRC_OUT_5_29 and I19548);
	I19555<= not (WX5786 and CRC_OUT_5_28);
	I19556<= not (WX5786 and I19555);
	I19557<= not (CRC_OUT_5_28 and I19555);
	I19562<= not (WX5787 and CRC_OUT_5_27);
	I19563<= not (WX5787 and I19562);
	I19564<= not (CRC_OUT_5_27 and I19562);
	I19569<= not (WX5788 and CRC_OUT_5_26);
	I19570<= not (WX5788 and I19569);
	I19571<= not (CRC_OUT_5_26 and I19569);
	I19576<= not (WX5789 and CRC_OUT_5_25);
	I19577<= not (WX5789 and I19576);
	I19578<= not (CRC_OUT_5_25 and I19576);
	I19583<= not (WX5790 and CRC_OUT_5_24);
	I19584<= not (WX5790 and I19583);
	I19585<= not (CRC_OUT_5_24 and I19583);
	I19590<= not (WX5791 and CRC_OUT_5_23);
	I19591<= not (WX5791 and I19590);
	I19592<= not (CRC_OUT_5_23 and I19590);
	I19597<= not (WX5792 and CRC_OUT_5_22);
	I19598<= not (WX5792 and I19597);
	I19599<= not (CRC_OUT_5_22 and I19597);
	I19604<= not (WX5793 and CRC_OUT_5_21);
	I19605<= not (WX5793 and I19604);
	I19606<= not (CRC_OUT_5_21 and I19604);
	I19611<= not (WX5794 and CRC_OUT_5_20);
	I19612<= not (WX5794 and I19611);
	I19613<= not (CRC_OUT_5_20 and I19611);
	I19618<= not (WX5795 and CRC_OUT_5_19);
	I19619<= not (WX5795 and I19618);
	I19620<= not (CRC_OUT_5_19 and I19618);
	I19625<= not (WX5796 and CRC_OUT_5_18);
	I19626<= not (WX5796 and I19625);
	I19627<= not (CRC_OUT_5_18 and I19625);
	I19632<= not (WX5797 and CRC_OUT_5_17);
	I19633<= not (WX5797 and I19632);
	I19634<= not (CRC_OUT_5_17 and I19632);
	I19639<= not (WX5798 and CRC_OUT_5_16);
	I19640<= not (WX5798 and I19639);
	I19641<= not (CRC_OUT_5_16 and I19639);
	I19646<= not (WX5800 and CRC_OUT_5_14);
	I19647<= not (WX5800 and I19646);
	I19648<= not (CRC_OUT_5_14 and I19646);
	I19653<= not (WX5801 and CRC_OUT_5_13);
	I19654<= not (WX5801 and I19653);
	I19655<= not (CRC_OUT_5_13 and I19653);
	I19660<= not (WX5802 and CRC_OUT_5_12);
	I19661<= not (WX5802 and I19660);
	I19662<= not (CRC_OUT_5_12 and I19660);
	I19667<= not (WX5803 and CRC_OUT_5_11);
	I19668<= not (WX5803 and I19667);
	I19669<= not (CRC_OUT_5_11 and I19667);
	I19674<= not (WX5805 and CRC_OUT_5_9);
	I19675<= not (WX5805 and I19674);
	I19676<= not (CRC_OUT_5_9 and I19674);
	I19681<= not (WX5806 and CRC_OUT_5_8);
	I19682<= not (WX5806 and I19681);
	I19683<= not (CRC_OUT_5_8 and I19681);
	I19688<= not (WX5807 and CRC_OUT_5_7);
	I19689<= not (WX5807 and I19688);
	I19690<= not (CRC_OUT_5_7 and I19688);
	I19695<= not (WX5808 and CRC_OUT_5_6);
	I19696<= not (WX5808 and I19695);
	I19697<= not (CRC_OUT_5_6 and I19695);
	I19702<= not (WX5809 and CRC_OUT_5_5);
	I19703<= not (WX5809 and I19702);
	I19704<= not (CRC_OUT_5_5 and I19702);
	I19709<= not (WX5810 and CRC_OUT_5_4);
	I19710<= not (WX5810 and I19709);
	I19711<= not (CRC_OUT_5_4 and I19709);
	I19716<= not (WX5812 and CRC_OUT_5_2);
	I19717<= not (WX5812 and I19716);
	I19718<= not (CRC_OUT_5_2 and I19716);
	I19723<= not (WX5813 and CRC_OUT_5_1);
	I19724<= not (WX5813 and I19723);
	I19725<= not (CRC_OUT_5_1 and I19723);
	I19730<= not (WX5814 and CRC_OUT_5_0);
	I19731<= not (WX5814 and I19730);
	I19732<= not (CRC_OUT_5_0 and I19730);
	I22011<= not (I22021 and I22022);
	I22012<= not (I22014 and I22015);
	I22013<= not (WX7466 and WX7110);
	I22014<= not (WX7466 and I22013);
	I22015<= not (WX7110 and I22013);
	I22020<= not (WX7174 and I22012);
	I22021<= not (WX7174 and I22020);
	I22022<= not (I22012 and I22020);
	I22027<= not (I22029 and I22030);
	I22028<= not (WX7238 and WX7302);
	I22029<= not (WX7238 and I22028);
	I22030<= not (WX7302 and I22028);
	I22035<= not (I22011 and I22027);
	I22036<= not (I22011 and I22035);
	I22037<= not (I22027 and I22035);
	I22042<= not (I22052 and I22053);
	I22043<= not (I22045 and I22046);
	I22044<= not (WX7466 and WX7112);
	I22045<= not (WX7466 and I22044);
	I22046<= not (WX7112 and I22044);
	I22051<= not (WX7176 and I22043);
	I22052<= not (WX7176 and I22051);
	I22053<= not (I22043 and I22051);
	I22058<= not (I22060 and I22061);
	I22059<= not (WX7240 and WX7304);
	I22060<= not (WX7240 and I22059);
	I22061<= not (WX7304 and I22059);
	I22066<= not (I22042 and I22058);
	I22067<= not (I22042 and I22066);
	I22068<= not (I22058 and I22066);
	I22073<= not (I22083 and I22084);
	I22074<= not (I22076 and I22077);
	I22075<= not (WX7466 and WX7114);
	I22076<= not (WX7466 and I22075);
	I22077<= not (WX7114 and I22075);
	I22082<= not (WX7178 and I22074);
	I22083<= not (WX7178 and I22082);
	I22084<= not (I22074 and I22082);
	I22089<= not (I22091 and I22092);
	I22090<= not (WX7242 and WX7306);
	I22091<= not (WX7242 and I22090);
	I22092<= not (WX7306 and I22090);
	I22097<= not (I22073 and I22089);
	I22098<= not (I22073 and I22097);
	I22099<= not (I22089 and I22097);
	I22104<= not (I22114 and I22115);
	I22105<= not (I22107 and I22108);
	I22106<= not (WX7466 and WX7116);
	I22107<= not (WX7466 and I22106);
	I22108<= not (WX7116 and I22106);
	I22113<= not (WX7180 and I22105);
	I22114<= not (WX7180 and I22113);
	I22115<= not (I22105 and I22113);
	I22120<= not (I22122 and I22123);
	I22121<= not (WX7244 and WX7308);
	I22122<= not (WX7244 and I22121);
	I22123<= not (WX7308 and I22121);
	I22128<= not (I22104 and I22120);
	I22129<= not (I22104 and I22128);
	I22130<= not (I22120 and I22128);
	I22135<= not (I22145 and I22146);
	I22136<= not (I22138 and I22139);
	I22137<= not (WX7466 and WX7118);
	I22138<= not (WX7466 and I22137);
	I22139<= not (WX7118 and I22137);
	I22144<= not (WX7182 and I22136);
	I22145<= not (WX7182 and I22144);
	I22146<= not (I22136 and I22144);
	I22151<= not (I22153 and I22154);
	I22152<= not (WX7246 and WX7310);
	I22153<= not (WX7246 and I22152);
	I22154<= not (WX7310 and I22152);
	I22159<= not (I22135 and I22151);
	I22160<= not (I22135 and I22159);
	I22161<= not (I22151 and I22159);
	I22166<= not (I22176 and I22177);
	I22167<= not (I22169 and I22170);
	I22168<= not (WX7466 and WX7120);
	I22169<= not (WX7466 and I22168);
	I22170<= not (WX7120 and I22168);
	I22175<= not (WX7184 and I22167);
	I22176<= not (WX7184 and I22175);
	I22177<= not (I22167 and I22175);
	I22182<= not (I22184 and I22185);
	I22183<= not (WX7248 and WX7312);
	I22184<= not (WX7248 and I22183);
	I22185<= not (WX7312 and I22183);
	I22190<= not (I22166 and I22182);
	I22191<= not (I22166 and I22190);
	I22192<= not (I22182 and I22190);
	I22197<= not (I22207 and I22208);
	I22198<= not (I22200 and I22201);
	I22199<= not (WX7466 and WX7122);
	I22200<= not (WX7466 and I22199);
	I22201<= not (WX7122 and I22199);
	I22206<= not (WX7186 and I22198);
	I22207<= not (WX7186 and I22206);
	I22208<= not (I22198 and I22206);
	I22213<= not (I22215 and I22216);
	I22214<= not (WX7250 and WX7314);
	I22215<= not (WX7250 and I22214);
	I22216<= not (WX7314 and I22214);
	I22221<= not (I22197 and I22213);
	I22222<= not (I22197 and I22221);
	I22223<= not (I22213 and I22221);
	I22228<= not (I22238 and I22239);
	I22229<= not (I22231 and I22232);
	I22230<= not (WX7466 and WX7124);
	I22231<= not (WX7466 and I22230);
	I22232<= not (WX7124 and I22230);
	I22237<= not (WX7188 and I22229);
	I22238<= not (WX7188 and I22237);
	I22239<= not (I22229 and I22237);
	I22244<= not (I22246 and I22247);
	I22245<= not (WX7252 and WX7316);
	I22246<= not (WX7252 and I22245);
	I22247<= not (WX7316 and I22245);
	I22252<= not (I22228 and I22244);
	I22253<= not (I22228 and I22252);
	I22254<= not (I22244 and I22252);
	I22259<= not (I22269 and I22270);
	I22260<= not (I22262 and I22263);
	I22261<= not (WX7466 and WX7126);
	I22262<= not (WX7466 and I22261);
	I22263<= not (WX7126 and I22261);
	I22268<= not (WX7190 and I22260);
	I22269<= not (WX7190 and I22268);
	I22270<= not (I22260 and I22268);
	I22275<= not (I22277 and I22278);
	I22276<= not (WX7254 and WX7318);
	I22277<= not (WX7254 and I22276);
	I22278<= not (WX7318 and I22276);
	I22283<= not (I22259 and I22275);
	I22284<= not (I22259 and I22283);
	I22285<= not (I22275 and I22283);
	I22290<= not (I22300 and I22301);
	I22291<= not (I22293 and I22294);
	I22292<= not (WX7466 and WX7128);
	I22293<= not (WX7466 and I22292);
	I22294<= not (WX7128 and I22292);
	I22299<= not (WX7192 and I22291);
	I22300<= not (WX7192 and I22299);
	I22301<= not (I22291 and I22299);
	I22306<= not (I22308 and I22309);
	I22307<= not (WX7256 and WX7320);
	I22308<= not (WX7256 and I22307);
	I22309<= not (WX7320 and I22307);
	I22314<= not (I22290 and I22306);
	I22315<= not (I22290 and I22314);
	I22316<= not (I22306 and I22314);
	I22321<= not (I22331 and I22332);
	I22322<= not (I22324 and I22325);
	I22323<= not (WX7466 and WX7130);
	I22324<= not (WX7466 and I22323);
	I22325<= not (WX7130 and I22323);
	I22330<= not (WX7194 and I22322);
	I22331<= not (WX7194 and I22330);
	I22332<= not (I22322 and I22330);
	I22337<= not (I22339 and I22340);
	I22338<= not (WX7258 and WX7322);
	I22339<= not (WX7258 and I22338);
	I22340<= not (WX7322 and I22338);
	I22345<= not (I22321 and I22337);
	I22346<= not (I22321 and I22345);
	I22347<= not (I22337 and I22345);
	I22352<= not (I22362 and I22363);
	I22353<= not (I22355 and I22356);
	I22354<= not (WX7466 and WX7132);
	I22355<= not (WX7466 and I22354);
	I22356<= not (WX7132 and I22354);
	I22361<= not (WX7196 and I22353);
	I22362<= not (WX7196 and I22361);
	I22363<= not (I22353 and I22361);
	I22368<= not (I22370 and I22371);
	I22369<= not (WX7260 and WX7324);
	I22370<= not (WX7260 and I22369);
	I22371<= not (WX7324 and I22369);
	I22376<= not (I22352 and I22368);
	I22377<= not (I22352 and I22376);
	I22378<= not (I22368 and I22376);
	I22383<= not (I22393 and I22394);
	I22384<= not (I22386 and I22387);
	I22385<= not (WX7466 and WX7134);
	I22386<= not (WX7466 and I22385);
	I22387<= not (WX7134 and I22385);
	I22392<= not (WX7198 and I22384);
	I22393<= not (WX7198 and I22392);
	I22394<= not (I22384 and I22392);
	I22399<= not (I22401 and I22402);
	I22400<= not (WX7262 and WX7326);
	I22401<= not (WX7262 and I22400);
	I22402<= not (WX7326 and I22400);
	I22407<= not (I22383 and I22399);
	I22408<= not (I22383 and I22407);
	I22409<= not (I22399 and I22407);
	I22414<= not (I22424 and I22425);
	I22415<= not (I22417 and I22418);
	I22416<= not (WX7466 and WX7136);
	I22417<= not (WX7466 and I22416);
	I22418<= not (WX7136 and I22416);
	I22423<= not (WX7200 and I22415);
	I22424<= not (WX7200 and I22423);
	I22425<= not (I22415 and I22423);
	I22430<= not (I22432 and I22433);
	I22431<= not (WX7264 and WX7328);
	I22432<= not (WX7264 and I22431);
	I22433<= not (WX7328 and I22431);
	I22438<= not (I22414 and I22430);
	I22439<= not (I22414 and I22438);
	I22440<= not (I22430 and I22438);
	I22445<= not (I22455 and I22456);
	I22446<= not (I22448 and I22449);
	I22447<= not (WX7466 and WX7138);
	I22448<= not (WX7466 and I22447);
	I22449<= not (WX7138 and I22447);
	I22454<= not (WX7202 and I22446);
	I22455<= not (WX7202 and I22454);
	I22456<= not (I22446 and I22454);
	I22461<= not (I22463 and I22464);
	I22462<= not (WX7266 and WX7330);
	I22463<= not (WX7266 and I22462);
	I22464<= not (WX7330 and I22462);
	I22469<= not (I22445 and I22461);
	I22470<= not (I22445 and I22469);
	I22471<= not (I22461 and I22469);
	I22476<= not (I22486 and I22487);
	I22477<= not (I22479 and I22480);
	I22478<= not (WX7466 and WX7140);
	I22479<= not (WX7466 and I22478);
	I22480<= not (WX7140 and I22478);
	I22485<= not (WX7204 and I22477);
	I22486<= not (WX7204 and I22485);
	I22487<= not (I22477 and I22485);
	I22492<= not (I22494 and I22495);
	I22493<= not (WX7268 and WX7332);
	I22494<= not (WX7268 and I22493);
	I22495<= not (WX7332 and I22493);
	I22500<= not (I22476 and I22492);
	I22501<= not (I22476 and I22500);
	I22502<= not (I22492 and I22500);
	I22507<= not (I22517 and I22518);
	I22508<= not (I22510 and I22511);
	I22509<= not (WX7467 and WX7142);
	I22510<= not (WX7467 and I22509);
	I22511<= not (WX7142 and I22509);
	I22516<= not (WX7206 and I22508);
	I22517<= not (WX7206 and I22516);
	I22518<= not (I22508 and I22516);
	I22523<= not (I22525 and I22526);
	I22524<= not (WX7270 and WX7334);
	I22525<= not (WX7270 and I22524);
	I22526<= not (WX7334 and I22524);
	I22531<= not (I22507 and I22523);
	I22532<= not (I22507 and I22531);
	I22533<= not (I22523 and I22531);
	I22538<= not (I22548 and I22549);
	I22539<= not (I22541 and I22542);
	I22540<= not (WX7467 and WX7144);
	I22541<= not (WX7467 and I22540);
	I22542<= not (WX7144 and I22540);
	I22547<= not (WX7208 and I22539);
	I22548<= not (WX7208 and I22547);
	I22549<= not (I22539 and I22547);
	I22554<= not (I22556 and I22557);
	I22555<= not (WX7272 and WX7336);
	I22556<= not (WX7272 and I22555);
	I22557<= not (WX7336 and I22555);
	I22562<= not (I22538 and I22554);
	I22563<= not (I22538 and I22562);
	I22564<= not (I22554 and I22562);
	I22569<= not (I22579 and I22580);
	I22570<= not (I22572 and I22573);
	I22571<= not (WX7467 and WX7146);
	I22572<= not (WX7467 and I22571);
	I22573<= not (WX7146 and I22571);
	I22578<= not (WX7210 and I22570);
	I22579<= not (WX7210 and I22578);
	I22580<= not (I22570 and I22578);
	I22585<= not (I22587 and I22588);
	I22586<= not (WX7274 and WX7338);
	I22587<= not (WX7274 and I22586);
	I22588<= not (WX7338 and I22586);
	I22593<= not (I22569 and I22585);
	I22594<= not (I22569 and I22593);
	I22595<= not (I22585 and I22593);
	I22600<= not (I22610 and I22611);
	I22601<= not (I22603 and I22604);
	I22602<= not (WX7467 and WX7148);
	I22603<= not (WX7467 and I22602);
	I22604<= not (WX7148 and I22602);
	I22609<= not (WX7212 and I22601);
	I22610<= not (WX7212 and I22609);
	I22611<= not (I22601 and I22609);
	I22616<= not (I22618 and I22619);
	I22617<= not (WX7276 and WX7340);
	I22618<= not (WX7276 and I22617);
	I22619<= not (WX7340 and I22617);
	I22624<= not (I22600 and I22616);
	I22625<= not (I22600 and I22624);
	I22626<= not (I22616 and I22624);
	I22631<= not (I22641 and I22642);
	I22632<= not (I22634 and I22635);
	I22633<= not (WX7467 and WX7150);
	I22634<= not (WX7467 and I22633);
	I22635<= not (WX7150 and I22633);
	I22640<= not (WX7214 and I22632);
	I22641<= not (WX7214 and I22640);
	I22642<= not (I22632 and I22640);
	I22647<= not (I22649 and I22650);
	I22648<= not (WX7278 and WX7342);
	I22649<= not (WX7278 and I22648);
	I22650<= not (WX7342 and I22648);
	I22655<= not (I22631 and I22647);
	I22656<= not (I22631 and I22655);
	I22657<= not (I22647 and I22655);
	I22662<= not (I22672 and I22673);
	I22663<= not (I22665 and I22666);
	I22664<= not (WX7467 and WX7152);
	I22665<= not (WX7467 and I22664);
	I22666<= not (WX7152 and I22664);
	I22671<= not (WX7216 and I22663);
	I22672<= not (WX7216 and I22671);
	I22673<= not (I22663 and I22671);
	I22678<= not (I22680 and I22681);
	I22679<= not (WX7280 and WX7344);
	I22680<= not (WX7280 and I22679);
	I22681<= not (WX7344 and I22679);
	I22686<= not (I22662 and I22678);
	I22687<= not (I22662 and I22686);
	I22688<= not (I22678 and I22686);
	I22693<= not (I22703 and I22704);
	I22694<= not (I22696 and I22697);
	I22695<= not (WX7467 and WX7154);
	I22696<= not (WX7467 and I22695);
	I22697<= not (WX7154 and I22695);
	I22702<= not (WX7218 and I22694);
	I22703<= not (WX7218 and I22702);
	I22704<= not (I22694 and I22702);
	I22709<= not (I22711 and I22712);
	I22710<= not (WX7282 and WX7346);
	I22711<= not (WX7282 and I22710);
	I22712<= not (WX7346 and I22710);
	I22717<= not (I22693 and I22709);
	I22718<= not (I22693 and I22717);
	I22719<= not (I22709 and I22717);
	I22724<= not (I22734 and I22735);
	I22725<= not (I22727 and I22728);
	I22726<= not (WX7467 and WX7156);
	I22727<= not (WX7467 and I22726);
	I22728<= not (WX7156 and I22726);
	I22733<= not (WX7220 and I22725);
	I22734<= not (WX7220 and I22733);
	I22735<= not (I22725 and I22733);
	I22740<= not (I22742 and I22743);
	I22741<= not (WX7284 and WX7348);
	I22742<= not (WX7284 and I22741);
	I22743<= not (WX7348 and I22741);
	I22748<= not (I22724 and I22740);
	I22749<= not (I22724 and I22748);
	I22750<= not (I22740 and I22748);
	I22755<= not (I22765 and I22766);
	I22756<= not (I22758 and I22759);
	I22757<= not (WX7467 and WX7158);
	I22758<= not (WX7467 and I22757);
	I22759<= not (WX7158 and I22757);
	I22764<= not (WX7222 and I22756);
	I22765<= not (WX7222 and I22764);
	I22766<= not (I22756 and I22764);
	I22771<= not (I22773 and I22774);
	I22772<= not (WX7286 and WX7350);
	I22773<= not (WX7286 and I22772);
	I22774<= not (WX7350 and I22772);
	I22779<= not (I22755 and I22771);
	I22780<= not (I22755 and I22779);
	I22781<= not (I22771 and I22779);
	I22786<= not (I22796 and I22797);
	I22787<= not (I22789 and I22790);
	I22788<= not (WX7467 and WX7160);
	I22789<= not (WX7467 and I22788);
	I22790<= not (WX7160 and I22788);
	I22795<= not (WX7224 and I22787);
	I22796<= not (WX7224 and I22795);
	I22797<= not (I22787 and I22795);
	I22802<= not (I22804 and I22805);
	I22803<= not (WX7288 and WX7352);
	I22804<= not (WX7288 and I22803);
	I22805<= not (WX7352 and I22803);
	I22810<= not (I22786 and I22802);
	I22811<= not (I22786 and I22810);
	I22812<= not (I22802 and I22810);
	I22817<= not (I22827 and I22828);
	I22818<= not (I22820 and I22821);
	I22819<= not (WX7467 and WX7162);
	I22820<= not (WX7467 and I22819);
	I22821<= not (WX7162 and I22819);
	I22826<= not (WX7226 and I22818);
	I22827<= not (WX7226 and I22826);
	I22828<= not (I22818 and I22826);
	I22833<= not (I22835 and I22836);
	I22834<= not (WX7290 and WX7354);
	I22835<= not (WX7290 and I22834);
	I22836<= not (WX7354 and I22834);
	I22841<= not (I22817 and I22833);
	I22842<= not (I22817 and I22841);
	I22843<= not (I22833 and I22841);
	I22848<= not (I22858 and I22859);
	I22849<= not (I22851 and I22852);
	I22850<= not (WX7467 and WX7164);
	I22851<= not (WX7467 and I22850);
	I22852<= not (WX7164 and I22850);
	I22857<= not (WX7228 and I22849);
	I22858<= not (WX7228 and I22857);
	I22859<= not (I22849 and I22857);
	I22864<= not (I22866 and I22867);
	I22865<= not (WX7292 and WX7356);
	I22866<= not (WX7292 and I22865);
	I22867<= not (WX7356 and I22865);
	I22872<= not (I22848 and I22864);
	I22873<= not (I22848 and I22872);
	I22874<= not (I22864 and I22872);
	I22879<= not (I22889 and I22890);
	I22880<= not (I22882 and I22883);
	I22881<= not (WX7467 and WX7166);
	I22882<= not (WX7467 and I22881);
	I22883<= not (WX7166 and I22881);
	I22888<= not (WX7230 and I22880);
	I22889<= not (WX7230 and I22888);
	I22890<= not (I22880 and I22888);
	I22895<= not (I22897 and I22898);
	I22896<= not (WX7294 and WX7358);
	I22897<= not (WX7294 and I22896);
	I22898<= not (WX7358 and I22896);
	I22903<= not (I22879 and I22895);
	I22904<= not (I22879 and I22903);
	I22905<= not (I22895 and I22903);
	I22910<= not (I22920 and I22921);
	I22911<= not (I22913 and I22914);
	I22912<= not (WX7467 and WX7168);
	I22913<= not (WX7467 and I22912);
	I22914<= not (WX7168 and I22912);
	I22919<= not (WX7232 and I22911);
	I22920<= not (WX7232 and I22919);
	I22921<= not (I22911 and I22919);
	I22926<= not (I22928 and I22929);
	I22927<= not (WX7296 and WX7360);
	I22928<= not (WX7296 and I22927);
	I22929<= not (WX7360 and I22927);
	I22934<= not (I22910 and I22926);
	I22935<= not (I22910 and I22934);
	I22936<= not (I22926 and I22934);
	I22941<= not (I22951 and I22952);
	I22942<= not (I22944 and I22945);
	I22943<= not (WX7467 and WX7170);
	I22944<= not (WX7467 and I22943);
	I22945<= not (WX7170 and I22943);
	I22950<= not (WX7234 and I22942);
	I22951<= not (WX7234 and I22950);
	I22952<= not (I22942 and I22950);
	I22957<= not (I22959 and I22960);
	I22958<= not (WX7298 and WX7362);
	I22959<= not (WX7298 and I22958);
	I22960<= not (WX7362 and I22958);
	I22965<= not (I22941 and I22957);
	I22966<= not (I22941 and I22965);
	I22967<= not (I22957 and I22965);
	I22972<= not (I22982 and I22983);
	I22973<= not (I22975 and I22976);
	I22974<= not (WX7467 and WX7172);
	I22975<= not (WX7467 and I22974);
	I22976<= not (WX7172 and I22974);
	I22981<= not (WX7236 and I22973);
	I22982<= not (WX7236 and I22981);
	I22983<= not (I22973 and I22981);
	I22988<= not (I22990 and I22991);
	I22989<= not (WX7300 and WX7364);
	I22990<= not (WX7300 and I22989);
	I22991<= not (WX7364 and I22989);
	I22996<= not (I22972 and I22988);
	I22997<= not (I22972 and I22996);
	I22998<= not (I22988 and I22996);
	I23077<= not (WX7045 and WX6950);
	I23078<= not (WX7045 and I23077);
	I23079<= not (WX6950 and I23077);
	I23090<= not (WX7046 and WX6952);
	I23091<= not (WX7046 and I23090);
	I23092<= not (WX6952 and I23090);
	I23103<= not (WX7047 and WX6954);
	I23104<= not (WX7047 and I23103);
	I23105<= not (WX6954 and I23103);
	I23116<= not (WX7048 and WX6956);
	I23117<= not (WX7048 and I23116);
	I23118<= not (WX6956 and I23116);
	I23129<= not (WX7049 and WX6958);
	I23130<= not (WX7049 and I23129);
	I23131<= not (WX6958 and I23129);
	I23142<= not (WX7050 and WX6960);
	I23143<= not (WX7050 and I23142);
	I23144<= not (WX6960 and I23142);
	I23155<= not (WX7051 and WX6962);
	I23156<= not (WX7051 and I23155);
	I23157<= not (WX6962 and I23155);
	I23168<= not (WX7052 and WX6964);
	I23169<= not (WX7052 and I23168);
	I23170<= not (WX6964 and I23168);
	I23181<= not (WX7053 and WX6966);
	I23182<= not (WX7053 and I23181);
	I23183<= not (WX6966 and I23181);
	I23194<= not (WX7054 and WX6968);
	I23195<= not (WX7054 and I23194);
	I23196<= not (WX6968 and I23194);
	I23207<= not (WX7055 and WX6970);
	I23208<= not (WX7055 and I23207);
	I23209<= not (WX6970 and I23207);
	I23220<= not (WX7056 and WX6972);
	I23221<= not (WX7056 and I23220);
	I23222<= not (WX6972 and I23220);
	I23233<= not (WX7057 and WX6974);
	I23234<= not (WX7057 and I23233);
	I23235<= not (WX6974 and I23233);
	I23246<= not (WX7058 and WX6976);
	I23247<= not (WX7058 and I23246);
	I23248<= not (WX6976 and I23246);
	I23259<= not (WX7059 and WX6978);
	I23260<= not (WX7059 and I23259);
	I23261<= not (WX6978 and I23259);
	I23272<= not (WX7060 and WX6980);
	I23273<= not (WX7060 and I23272);
	I23274<= not (WX6980 and I23272);
	I23285<= not (WX7061 and WX6982);
	I23286<= not (WX7061 and I23285);
	I23287<= not (WX6982 and I23285);
	I23298<= not (WX7062 and WX6984);
	I23299<= not (WX7062 and I23298);
	I23300<= not (WX6984 and I23298);
	I23311<= not (WX7063 and WX6986);
	I23312<= not (WX7063 and I23311);
	I23313<= not (WX6986 and I23311);
	I23324<= not (WX7064 and WX6988);
	I23325<= not (WX7064 and I23324);
	I23326<= not (WX6988 and I23324);
	I23337<= not (WX7065 and WX6990);
	I23338<= not (WX7065 and I23337);
	I23339<= not (WX6990 and I23337);
	I23350<= not (WX7066 and WX6992);
	I23351<= not (WX7066 and I23350);
	I23352<= not (WX6992 and I23350);
	I23363<= not (WX7067 and WX6994);
	I23364<= not (WX7067 and I23363);
	I23365<= not (WX6994 and I23363);
	I23376<= not (WX7068 and WX6996);
	I23377<= not (WX7068 and I23376);
	I23378<= not (WX6996 and I23376);
	I23389<= not (WX7069 and WX6998);
	I23390<= not (WX7069 and I23389);
	I23391<= not (WX6998 and I23389);
	I23402<= not (WX7070 and WX7000);
	I23403<= not (WX7070 and I23402);
	I23404<= not (WX7000 and I23402);
	I23415<= not (WX7071 and WX7002);
	I23416<= not (WX7071 and I23415);
	I23417<= not (WX7002 and I23415);
	I23428<= not (WX7072 and WX7004);
	I23429<= not (WX7072 and I23428);
	I23430<= not (WX7004 and I23428);
	I23441<= not (WX7073 and WX7006);
	I23442<= not (WX7073 and I23441);
	I23443<= not (WX7006 and I23441);
	I23454<= not (WX7074 and WX7008);
	I23455<= not (WX7074 and I23454);
	I23456<= not (WX7008 and I23454);
	I23467<= not (WX7075 and WX7010);
	I23468<= not (WX7075 and I23467);
	I23469<= not (WX7010 and I23467);
	I23480<= not (WX7076 and WX7012);
	I23481<= not (WX7076 and I23480);
	I23482<= not (WX7012 and I23480);
	I23494<= not (I23496 and I23497);
	I23495<= not (WX7092 and CRC_OUT_4_31);
	I23496<= not (WX7092 and I23495);
	I23497<= not (CRC_OUT_4_31 and I23495);
	I23502<= not (CRC_OUT_4_15 and I23494);
	I23503<= not (CRC_OUT_4_15 and I23502);
	I23504<= not (I23494 and I23502);
	I23509<= not (I23511 and I23512);
	I23510<= not (WX7097 and CRC_OUT_4_31);
	I23511<= not (WX7097 and I23510);
	I23512<= not (CRC_OUT_4_31 and I23510);
	I23517<= not (CRC_OUT_4_10 and I23509);
	I23518<= not (CRC_OUT_4_10 and I23517);
	I23519<= not (I23509 and I23517);
	I23524<= not (I23526 and I23527);
	I23525<= not (WX7104 and CRC_OUT_4_31);
	I23526<= not (WX7104 and I23525);
	I23527<= not (CRC_OUT_4_31 and I23525);
	I23532<= not (CRC_OUT_4_3 and I23524);
	I23533<= not (CRC_OUT_4_3 and I23532);
	I23534<= not (I23524 and I23532);
	I23539<= not (WX7108 and CRC_OUT_4_31);
	I23540<= not (WX7108 and I23539);
	I23541<= not (CRC_OUT_4_31 and I23539);
	I23546<= not (WX7077 and CRC_OUT_4_30);
	I23547<= not (WX7077 and I23546);
	I23548<= not (CRC_OUT_4_30 and I23546);
	I23553<= not (WX7078 and CRC_OUT_4_29);
	I23554<= not (WX7078 and I23553);
	I23555<= not (CRC_OUT_4_29 and I23553);
	I23560<= not (WX7079 and CRC_OUT_4_28);
	I23561<= not (WX7079 and I23560);
	I23562<= not (CRC_OUT_4_28 and I23560);
	I23567<= not (WX7080 and CRC_OUT_4_27);
	I23568<= not (WX7080 and I23567);
	I23569<= not (CRC_OUT_4_27 and I23567);
	I23574<= not (WX7081 and CRC_OUT_4_26);
	I23575<= not (WX7081 and I23574);
	I23576<= not (CRC_OUT_4_26 and I23574);
	I23581<= not (WX7082 and CRC_OUT_4_25);
	I23582<= not (WX7082 and I23581);
	I23583<= not (CRC_OUT_4_25 and I23581);
	I23588<= not (WX7083 and CRC_OUT_4_24);
	I23589<= not (WX7083 and I23588);
	I23590<= not (CRC_OUT_4_24 and I23588);
	I23595<= not (WX7084 and CRC_OUT_4_23);
	I23596<= not (WX7084 and I23595);
	I23597<= not (CRC_OUT_4_23 and I23595);
	I23602<= not (WX7085 and CRC_OUT_4_22);
	I23603<= not (WX7085 and I23602);
	I23604<= not (CRC_OUT_4_22 and I23602);
	I23609<= not (WX7086 and CRC_OUT_4_21);
	I23610<= not (WX7086 and I23609);
	I23611<= not (CRC_OUT_4_21 and I23609);
	I23616<= not (WX7087 and CRC_OUT_4_20);
	I23617<= not (WX7087 and I23616);
	I23618<= not (CRC_OUT_4_20 and I23616);
	I23623<= not (WX7088 and CRC_OUT_4_19);
	I23624<= not (WX7088 and I23623);
	I23625<= not (CRC_OUT_4_19 and I23623);
	I23630<= not (WX7089 and CRC_OUT_4_18);
	I23631<= not (WX7089 and I23630);
	I23632<= not (CRC_OUT_4_18 and I23630);
	I23637<= not (WX7090 and CRC_OUT_4_17);
	I23638<= not (WX7090 and I23637);
	I23639<= not (CRC_OUT_4_17 and I23637);
	I23644<= not (WX7091 and CRC_OUT_4_16);
	I23645<= not (WX7091 and I23644);
	I23646<= not (CRC_OUT_4_16 and I23644);
	I23651<= not (WX7093 and CRC_OUT_4_14);
	I23652<= not (WX7093 and I23651);
	I23653<= not (CRC_OUT_4_14 and I23651);
	I23658<= not (WX7094 and CRC_OUT_4_13);
	I23659<= not (WX7094 and I23658);
	I23660<= not (CRC_OUT_4_13 and I23658);
	I23665<= not (WX7095 and CRC_OUT_4_12);
	I23666<= not (WX7095 and I23665);
	I23667<= not (CRC_OUT_4_12 and I23665);
	I23672<= not (WX7096 and CRC_OUT_4_11);
	I23673<= not (WX7096 and I23672);
	I23674<= not (CRC_OUT_4_11 and I23672);
	I23679<= not (WX7098 and CRC_OUT_4_9);
	I23680<= not (WX7098 and I23679);
	I23681<= not (CRC_OUT_4_9 and I23679);
	I23686<= not (WX7099 and CRC_OUT_4_8);
	I23687<= not (WX7099 and I23686);
	I23688<= not (CRC_OUT_4_8 and I23686);
	I23693<= not (WX7100 and CRC_OUT_4_7);
	I23694<= not (WX7100 and I23693);
	I23695<= not (CRC_OUT_4_7 and I23693);
	I23700<= not (WX7101 and CRC_OUT_4_6);
	I23701<= not (WX7101 and I23700);
	I23702<= not (CRC_OUT_4_6 and I23700);
	I23707<= not (WX7102 and CRC_OUT_4_5);
	I23708<= not (WX7102 and I23707);
	I23709<= not (CRC_OUT_4_5 and I23707);
	I23714<= not (WX7103 and CRC_OUT_4_4);
	I23715<= not (WX7103 and I23714);
	I23716<= not (CRC_OUT_4_4 and I23714);
	I23721<= not (WX7105 and CRC_OUT_4_2);
	I23722<= not (WX7105 and I23721);
	I23723<= not (CRC_OUT_4_2 and I23721);
	I23728<= not (WX7106 and CRC_OUT_4_1);
	I23729<= not (WX7106 and I23728);
	I23730<= not (CRC_OUT_4_1 and I23728);
	I23735<= not (WX7107 and CRC_OUT_4_0);
	I23736<= not (WX7107 and I23735);
	I23737<= not (CRC_OUT_4_0 and I23735);
	I26016<= not (I26026 and I26027);
	I26017<= not (I26019 and I26020);
	I26018<= not (WX8759 and WX8403);
	I26019<= not (WX8759 and I26018);
	I26020<= not (WX8403 and I26018);
	I26025<= not (WX8467 and I26017);
	I26026<= not (WX8467 and I26025);
	I26027<= not (I26017 and I26025);
	I26032<= not (I26034 and I26035);
	I26033<= not (WX8531 and WX8595);
	I26034<= not (WX8531 and I26033);
	I26035<= not (WX8595 and I26033);
	I26040<= not (I26016 and I26032);
	I26041<= not (I26016 and I26040);
	I26042<= not (I26032 and I26040);
	I26047<= not (I26057 and I26058);
	I26048<= not (I26050 and I26051);
	I26049<= not (WX8759 and WX8405);
	I26050<= not (WX8759 and I26049);
	I26051<= not (WX8405 and I26049);
	I26056<= not (WX8469 and I26048);
	I26057<= not (WX8469 and I26056);
	I26058<= not (I26048 and I26056);
	I26063<= not (I26065 and I26066);
	I26064<= not (WX8533 and WX8597);
	I26065<= not (WX8533 and I26064);
	I26066<= not (WX8597 and I26064);
	I26071<= not (I26047 and I26063);
	I26072<= not (I26047 and I26071);
	I26073<= not (I26063 and I26071);
	I26078<= not (I26088 and I26089);
	I26079<= not (I26081 and I26082);
	I26080<= not (WX8759 and WX8407);
	I26081<= not (WX8759 and I26080);
	I26082<= not (WX8407 and I26080);
	I26087<= not (WX8471 and I26079);
	I26088<= not (WX8471 and I26087);
	I26089<= not (I26079 and I26087);
	I26094<= not (I26096 and I26097);
	I26095<= not (WX8535 and WX8599);
	I26096<= not (WX8535 and I26095);
	I26097<= not (WX8599 and I26095);
	I26102<= not (I26078 and I26094);
	I26103<= not (I26078 and I26102);
	I26104<= not (I26094 and I26102);
	I26109<= not (I26119 and I26120);
	I26110<= not (I26112 and I26113);
	I26111<= not (WX8759 and WX8409);
	I26112<= not (WX8759 and I26111);
	I26113<= not (WX8409 and I26111);
	I26118<= not (WX8473 and I26110);
	I26119<= not (WX8473 and I26118);
	I26120<= not (I26110 and I26118);
	I26125<= not (I26127 and I26128);
	I26126<= not (WX8537 and WX8601);
	I26127<= not (WX8537 and I26126);
	I26128<= not (WX8601 and I26126);
	I26133<= not (I26109 and I26125);
	I26134<= not (I26109 and I26133);
	I26135<= not (I26125 and I26133);
	I26140<= not (I26150 and I26151);
	I26141<= not (I26143 and I26144);
	I26142<= not (WX8759 and WX8411);
	I26143<= not (WX8759 and I26142);
	I26144<= not (WX8411 and I26142);
	I26149<= not (WX8475 and I26141);
	I26150<= not (WX8475 and I26149);
	I26151<= not (I26141 and I26149);
	I26156<= not (I26158 and I26159);
	I26157<= not (WX8539 and WX8603);
	I26158<= not (WX8539 and I26157);
	I26159<= not (WX8603 and I26157);
	I26164<= not (I26140 and I26156);
	I26165<= not (I26140 and I26164);
	I26166<= not (I26156 and I26164);
	I26171<= not (I26181 and I26182);
	I26172<= not (I26174 and I26175);
	I26173<= not (WX8759 and WX8413);
	I26174<= not (WX8759 and I26173);
	I26175<= not (WX8413 and I26173);
	I26180<= not (WX8477 and I26172);
	I26181<= not (WX8477 and I26180);
	I26182<= not (I26172 and I26180);
	I26187<= not (I26189 and I26190);
	I26188<= not (WX8541 and WX8605);
	I26189<= not (WX8541 and I26188);
	I26190<= not (WX8605 and I26188);
	I26195<= not (I26171 and I26187);
	I26196<= not (I26171 and I26195);
	I26197<= not (I26187 and I26195);
	I26202<= not (I26212 and I26213);
	I26203<= not (I26205 and I26206);
	I26204<= not (WX8759 and WX8415);
	I26205<= not (WX8759 and I26204);
	I26206<= not (WX8415 and I26204);
	I26211<= not (WX8479 and I26203);
	I26212<= not (WX8479 and I26211);
	I26213<= not (I26203 and I26211);
	I26218<= not (I26220 and I26221);
	I26219<= not (WX8543 and WX8607);
	I26220<= not (WX8543 and I26219);
	I26221<= not (WX8607 and I26219);
	I26226<= not (I26202 and I26218);
	I26227<= not (I26202 and I26226);
	I26228<= not (I26218 and I26226);
	I26233<= not (I26243 and I26244);
	I26234<= not (I26236 and I26237);
	I26235<= not (WX8759 and WX8417);
	I26236<= not (WX8759 and I26235);
	I26237<= not (WX8417 and I26235);
	I26242<= not (WX8481 and I26234);
	I26243<= not (WX8481 and I26242);
	I26244<= not (I26234 and I26242);
	I26249<= not (I26251 and I26252);
	I26250<= not (WX8545 and WX8609);
	I26251<= not (WX8545 and I26250);
	I26252<= not (WX8609 and I26250);
	I26257<= not (I26233 and I26249);
	I26258<= not (I26233 and I26257);
	I26259<= not (I26249 and I26257);
	I26264<= not (I26274 and I26275);
	I26265<= not (I26267 and I26268);
	I26266<= not (WX8759 and WX8419);
	I26267<= not (WX8759 and I26266);
	I26268<= not (WX8419 and I26266);
	I26273<= not (WX8483 and I26265);
	I26274<= not (WX8483 and I26273);
	I26275<= not (I26265 and I26273);
	I26280<= not (I26282 and I26283);
	I26281<= not (WX8547 and WX8611);
	I26282<= not (WX8547 and I26281);
	I26283<= not (WX8611 and I26281);
	I26288<= not (I26264 and I26280);
	I26289<= not (I26264 and I26288);
	I26290<= not (I26280 and I26288);
	I26295<= not (I26305 and I26306);
	I26296<= not (I26298 and I26299);
	I26297<= not (WX8759 and WX8421);
	I26298<= not (WX8759 and I26297);
	I26299<= not (WX8421 and I26297);
	I26304<= not (WX8485 and I26296);
	I26305<= not (WX8485 and I26304);
	I26306<= not (I26296 and I26304);
	I26311<= not (I26313 and I26314);
	I26312<= not (WX8549 and WX8613);
	I26313<= not (WX8549 and I26312);
	I26314<= not (WX8613 and I26312);
	I26319<= not (I26295 and I26311);
	I26320<= not (I26295 and I26319);
	I26321<= not (I26311 and I26319);
	I26326<= not (I26336 and I26337);
	I26327<= not (I26329 and I26330);
	I26328<= not (WX8759 and WX8423);
	I26329<= not (WX8759 and I26328);
	I26330<= not (WX8423 and I26328);
	I26335<= not (WX8487 and I26327);
	I26336<= not (WX8487 and I26335);
	I26337<= not (I26327 and I26335);
	I26342<= not (I26344 and I26345);
	I26343<= not (WX8551 and WX8615);
	I26344<= not (WX8551 and I26343);
	I26345<= not (WX8615 and I26343);
	I26350<= not (I26326 and I26342);
	I26351<= not (I26326 and I26350);
	I26352<= not (I26342 and I26350);
	I26357<= not (I26367 and I26368);
	I26358<= not (I26360 and I26361);
	I26359<= not (WX8759 and WX8425);
	I26360<= not (WX8759 and I26359);
	I26361<= not (WX8425 and I26359);
	I26366<= not (WX8489 and I26358);
	I26367<= not (WX8489 and I26366);
	I26368<= not (I26358 and I26366);
	I26373<= not (I26375 and I26376);
	I26374<= not (WX8553 and WX8617);
	I26375<= not (WX8553 and I26374);
	I26376<= not (WX8617 and I26374);
	I26381<= not (I26357 and I26373);
	I26382<= not (I26357 and I26381);
	I26383<= not (I26373 and I26381);
	I26388<= not (I26398 and I26399);
	I26389<= not (I26391 and I26392);
	I26390<= not (WX8759 and WX8427);
	I26391<= not (WX8759 and I26390);
	I26392<= not (WX8427 and I26390);
	I26397<= not (WX8491 and I26389);
	I26398<= not (WX8491 and I26397);
	I26399<= not (I26389 and I26397);
	I26404<= not (I26406 and I26407);
	I26405<= not (WX8555 and WX8619);
	I26406<= not (WX8555 and I26405);
	I26407<= not (WX8619 and I26405);
	I26412<= not (I26388 and I26404);
	I26413<= not (I26388 and I26412);
	I26414<= not (I26404 and I26412);
	I26419<= not (I26429 and I26430);
	I26420<= not (I26422 and I26423);
	I26421<= not (WX8759 and WX8429);
	I26422<= not (WX8759 and I26421);
	I26423<= not (WX8429 and I26421);
	I26428<= not (WX8493 and I26420);
	I26429<= not (WX8493 and I26428);
	I26430<= not (I26420 and I26428);
	I26435<= not (I26437 and I26438);
	I26436<= not (WX8557 and WX8621);
	I26437<= not (WX8557 and I26436);
	I26438<= not (WX8621 and I26436);
	I26443<= not (I26419 and I26435);
	I26444<= not (I26419 and I26443);
	I26445<= not (I26435 and I26443);
	I26450<= not (I26460 and I26461);
	I26451<= not (I26453 and I26454);
	I26452<= not (WX8759 and WX8431);
	I26453<= not (WX8759 and I26452);
	I26454<= not (WX8431 and I26452);
	I26459<= not (WX8495 and I26451);
	I26460<= not (WX8495 and I26459);
	I26461<= not (I26451 and I26459);
	I26466<= not (I26468 and I26469);
	I26467<= not (WX8559 and WX8623);
	I26468<= not (WX8559 and I26467);
	I26469<= not (WX8623 and I26467);
	I26474<= not (I26450 and I26466);
	I26475<= not (I26450 and I26474);
	I26476<= not (I26466 and I26474);
	I26481<= not (I26491 and I26492);
	I26482<= not (I26484 and I26485);
	I26483<= not (WX8759 and WX8433);
	I26484<= not (WX8759 and I26483);
	I26485<= not (WX8433 and I26483);
	I26490<= not (WX8497 and I26482);
	I26491<= not (WX8497 and I26490);
	I26492<= not (I26482 and I26490);
	I26497<= not (I26499 and I26500);
	I26498<= not (WX8561 and WX8625);
	I26499<= not (WX8561 and I26498);
	I26500<= not (WX8625 and I26498);
	I26505<= not (I26481 and I26497);
	I26506<= not (I26481 and I26505);
	I26507<= not (I26497 and I26505);
	I26512<= not (I26522 and I26523);
	I26513<= not (I26515 and I26516);
	I26514<= not (WX8760 and WX8435);
	I26515<= not (WX8760 and I26514);
	I26516<= not (WX8435 and I26514);
	I26521<= not (WX8499 and I26513);
	I26522<= not (WX8499 and I26521);
	I26523<= not (I26513 and I26521);
	I26528<= not (I26530 and I26531);
	I26529<= not (WX8563 and WX8627);
	I26530<= not (WX8563 and I26529);
	I26531<= not (WX8627 and I26529);
	I26536<= not (I26512 and I26528);
	I26537<= not (I26512 and I26536);
	I26538<= not (I26528 and I26536);
	I26543<= not (I26553 and I26554);
	I26544<= not (I26546 and I26547);
	I26545<= not (WX8760 and WX8437);
	I26546<= not (WX8760 and I26545);
	I26547<= not (WX8437 and I26545);
	I26552<= not (WX8501 and I26544);
	I26553<= not (WX8501 and I26552);
	I26554<= not (I26544 and I26552);
	I26559<= not (I26561 and I26562);
	I26560<= not (WX8565 and WX8629);
	I26561<= not (WX8565 and I26560);
	I26562<= not (WX8629 and I26560);
	I26567<= not (I26543 and I26559);
	I26568<= not (I26543 and I26567);
	I26569<= not (I26559 and I26567);
	I26574<= not (I26584 and I26585);
	I26575<= not (I26577 and I26578);
	I26576<= not (WX8760 and WX8439);
	I26577<= not (WX8760 and I26576);
	I26578<= not (WX8439 and I26576);
	I26583<= not (WX8503 and I26575);
	I26584<= not (WX8503 and I26583);
	I26585<= not (I26575 and I26583);
	I26590<= not (I26592 and I26593);
	I26591<= not (WX8567 and WX8631);
	I26592<= not (WX8567 and I26591);
	I26593<= not (WX8631 and I26591);
	I26598<= not (I26574 and I26590);
	I26599<= not (I26574 and I26598);
	I26600<= not (I26590 and I26598);
	I26605<= not (I26615 and I26616);
	I26606<= not (I26608 and I26609);
	I26607<= not (WX8760 and WX8441);
	I26608<= not (WX8760 and I26607);
	I26609<= not (WX8441 and I26607);
	I26614<= not (WX8505 and I26606);
	I26615<= not (WX8505 and I26614);
	I26616<= not (I26606 and I26614);
	I26621<= not (I26623 and I26624);
	I26622<= not (WX8569 and WX8633);
	I26623<= not (WX8569 and I26622);
	I26624<= not (WX8633 and I26622);
	I26629<= not (I26605 and I26621);
	I26630<= not (I26605 and I26629);
	I26631<= not (I26621 and I26629);
	I26636<= not (I26646 and I26647);
	I26637<= not (I26639 and I26640);
	I26638<= not (WX8760 and WX8443);
	I26639<= not (WX8760 and I26638);
	I26640<= not (WX8443 and I26638);
	I26645<= not (WX8507 and I26637);
	I26646<= not (WX8507 and I26645);
	I26647<= not (I26637 and I26645);
	I26652<= not (I26654 and I26655);
	I26653<= not (WX8571 and WX8635);
	I26654<= not (WX8571 and I26653);
	I26655<= not (WX8635 and I26653);
	I26660<= not (I26636 and I26652);
	I26661<= not (I26636 and I26660);
	I26662<= not (I26652 and I26660);
	I26667<= not (I26677 and I26678);
	I26668<= not (I26670 and I26671);
	I26669<= not (WX8760 and WX8445);
	I26670<= not (WX8760 and I26669);
	I26671<= not (WX8445 and I26669);
	I26676<= not (WX8509 and I26668);
	I26677<= not (WX8509 and I26676);
	I26678<= not (I26668 and I26676);
	I26683<= not (I26685 and I26686);
	I26684<= not (WX8573 and WX8637);
	I26685<= not (WX8573 and I26684);
	I26686<= not (WX8637 and I26684);
	I26691<= not (I26667 and I26683);
	I26692<= not (I26667 and I26691);
	I26693<= not (I26683 and I26691);
	I26698<= not (I26708 and I26709);
	I26699<= not (I26701 and I26702);
	I26700<= not (WX8760 and WX8447);
	I26701<= not (WX8760 and I26700);
	I26702<= not (WX8447 and I26700);
	I26707<= not (WX8511 and I26699);
	I26708<= not (WX8511 and I26707);
	I26709<= not (I26699 and I26707);
	I26714<= not (I26716 and I26717);
	I26715<= not (WX8575 and WX8639);
	I26716<= not (WX8575 and I26715);
	I26717<= not (WX8639 and I26715);
	I26722<= not (I26698 and I26714);
	I26723<= not (I26698 and I26722);
	I26724<= not (I26714 and I26722);
	I26729<= not (I26739 and I26740);
	I26730<= not (I26732 and I26733);
	I26731<= not (WX8760 and WX8449);
	I26732<= not (WX8760 and I26731);
	I26733<= not (WX8449 and I26731);
	I26738<= not (WX8513 and I26730);
	I26739<= not (WX8513 and I26738);
	I26740<= not (I26730 and I26738);
	I26745<= not (I26747 and I26748);
	I26746<= not (WX8577 and WX8641);
	I26747<= not (WX8577 and I26746);
	I26748<= not (WX8641 and I26746);
	I26753<= not (I26729 and I26745);
	I26754<= not (I26729 and I26753);
	I26755<= not (I26745 and I26753);
	I26760<= not (I26770 and I26771);
	I26761<= not (I26763 and I26764);
	I26762<= not (WX8760 and WX8451);
	I26763<= not (WX8760 and I26762);
	I26764<= not (WX8451 and I26762);
	I26769<= not (WX8515 and I26761);
	I26770<= not (WX8515 and I26769);
	I26771<= not (I26761 and I26769);
	I26776<= not (I26778 and I26779);
	I26777<= not (WX8579 and WX8643);
	I26778<= not (WX8579 and I26777);
	I26779<= not (WX8643 and I26777);
	I26784<= not (I26760 and I26776);
	I26785<= not (I26760 and I26784);
	I26786<= not (I26776 and I26784);
	I26791<= not (I26801 and I26802);
	I26792<= not (I26794 and I26795);
	I26793<= not (WX8760 and WX8453);
	I26794<= not (WX8760 and I26793);
	I26795<= not (WX8453 and I26793);
	I26800<= not (WX8517 and I26792);
	I26801<= not (WX8517 and I26800);
	I26802<= not (I26792 and I26800);
	I26807<= not (I26809 and I26810);
	I26808<= not (WX8581 and WX8645);
	I26809<= not (WX8581 and I26808);
	I26810<= not (WX8645 and I26808);
	I26815<= not (I26791 and I26807);
	I26816<= not (I26791 and I26815);
	I26817<= not (I26807 and I26815);
	I26822<= not (I26832 and I26833);
	I26823<= not (I26825 and I26826);
	I26824<= not (WX8760 and WX8455);
	I26825<= not (WX8760 and I26824);
	I26826<= not (WX8455 and I26824);
	I26831<= not (WX8519 and I26823);
	I26832<= not (WX8519 and I26831);
	I26833<= not (I26823 and I26831);
	I26838<= not (I26840 and I26841);
	I26839<= not (WX8583 and WX8647);
	I26840<= not (WX8583 and I26839);
	I26841<= not (WX8647 and I26839);
	I26846<= not (I26822 and I26838);
	I26847<= not (I26822 and I26846);
	I26848<= not (I26838 and I26846);
	I26853<= not (I26863 and I26864);
	I26854<= not (I26856 and I26857);
	I26855<= not (WX8760 and WX8457);
	I26856<= not (WX8760 and I26855);
	I26857<= not (WX8457 and I26855);
	I26862<= not (WX8521 and I26854);
	I26863<= not (WX8521 and I26862);
	I26864<= not (I26854 and I26862);
	I26869<= not (I26871 and I26872);
	I26870<= not (WX8585 and WX8649);
	I26871<= not (WX8585 and I26870);
	I26872<= not (WX8649 and I26870);
	I26877<= not (I26853 and I26869);
	I26878<= not (I26853 and I26877);
	I26879<= not (I26869 and I26877);
	I26884<= not (I26894 and I26895);
	I26885<= not (I26887 and I26888);
	I26886<= not (WX8760 and WX8459);
	I26887<= not (WX8760 and I26886);
	I26888<= not (WX8459 and I26886);
	I26893<= not (WX8523 and I26885);
	I26894<= not (WX8523 and I26893);
	I26895<= not (I26885 and I26893);
	I26900<= not (I26902 and I26903);
	I26901<= not (WX8587 and WX8651);
	I26902<= not (WX8587 and I26901);
	I26903<= not (WX8651 and I26901);
	I26908<= not (I26884 and I26900);
	I26909<= not (I26884 and I26908);
	I26910<= not (I26900 and I26908);
	I26915<= not (I26925 and I26926);
	I26916<= not (I26918 and I26919);
	I26917<= not (WX8760 and WX8461);
	I26918<= not (WX8760 and I26917);
	I26919<= not (WX8461 and I26917);
	I26924<= not (WX8525 and I26916);
	I26925<= not (WX8525 and I26924);
	I26926<= not (I26916 and I26924);
	I26931<= not (I26933 and I26934);
	I26932<= not (WX8589 and WX8653);
	I26933<= not (WX8589 and I26932);
	I26934<= not (WX8653 and I26932);
	I26939<= not (I26915 and I26931);
	I26940<= not (I26915 and I26939);
	I26941<= not (I26931 and I26939);
	I26946<= not (I26956 and I26957);
	I26947<= not (I26949 and I26950);
	I26948<= not (WX8760 and WX8463);
	I26949<= not (WX8760 and I26948);
	I26950<= not (WX8463 and I26948);
	I26955<= not (WX8527 and I26947);
	I26956<= not (WX8527 and I26955);
	I26957<= not (I26947 and I26955);
	I26962<= not (I26964 and I26965);
	I26963<= not (WX8591 and WX8655);
	I26964<= not (WX8591 and I26963);
	I26965<= not (WX8655 and I26963);
	I26970<= not (I26946 and I26962);
	I26971<= not (I26946 and I26970);
	I26972<= not (I26962 and I26970);
	I26977<= not (I26987 and I26988);
	I26978<= not (I26980 and I26981);
	I26979<= not (WX8760 and WX8465);
	I26980<= not (WX8760 and I26979);
	I26981<= not (WX8465 and I26979);
	I26986<= not (WX8529 and I26978);
	I26987<= not (WX8529 and I26986);
	I26988<= not (I26978 and I26986);
	I26993<= not (I26995 and I26996);
	I26994<= not (WX8593 and WX8657);
	I26995<= not (WX8593 and I26994);
	I26996<= not (WX8657 and I26994);
	I27001<= not (I26977 and I26993);
	I27002<= not (I26977 and I27001);
	I27003<= not (I26993 and I27001);
	I27082<= not (WX8338 and WX8243);
	I27083<= not (WX8338 and I27082);
	I27084<= not (WX8243 and I27082);
	I27095<= not (WX8339 and WX8245);
	I27096<= not (WX8339 and I27095);
	I27097<= not (WX8245 and I27095);
	I27108<= not (WX8340 and WX8247);
	I27109<= not (WX8340 and I27108);
	I27110<= not (WX8247 and I27108);
	I27121<= not (WX8341 and WX8249);
	I27122<= not (WX8341 and I27121);
	I27123<= not (WX8249 and I27121);
	I27134<= not (WX8342 and WX8251);
	I27135<= not (WX8342 and I27134);
	I27136<= not (WX8251 and I27134);
	I27147<= not (WX8343 and WX8253);
	I27148<= not (WX8343 and I27147);
	I27149<= not (WX8253 and I27147);
	I27160<= not (WX8344 and WX8255);
	I27161<= not (WX8344 and I27160);
	I27162<= not (WX8255 and I27160);
	I27173<= not (WX8345 and WX8257);
	I27174<= not (WX8345 and I27173);
	I27175<= not (WX8257 and I27173);
	I27186<= not (WX8346 and WX8259);
	I27187<= not (WX8346 and I27186);
	I27188<= not (WX8259 and I27186);
	I27199<= not (WX8347 and WX8261);
	I27200<= not (WX8347 and I27199);
	I27201<= not (WX8261 and I27199);
	I27212<= not (WX8348 and WX8263);
	I27213<= not (WX8348 and I27212);
	I27214<= not (WX8263 and I27212);
	I27225<= not (WX8349 and WX8265);
	I27226<= not (WX8349 and I27225);
	I27227<= not (WX8265 and I27225);
	I27238<= not (WX8350 and WX8267);
	I27239<= not (WX8350 and I27238);
	I27240<= not (WX8267 and I27238);
	I27251<= not (WX8351 and WX8269);
	I27252<= not (WX8351 and I27251);
	I27253<= not (WX8269 and I27251);
	I27264<= not (WX8352 and WX8271);
	I27265<= not (WX8352 and I27264);
	I27266<= not (WX8271 and I27264);
	I27277<= not (WX8353 and WX8273);
	I27278<= not (WX8353 and I27277);
	I27279<= not (WX8273 and I27277);
	I27290<= not (WX8354 and WX8275);
	I27291<= not (WX8354 and I27290);
	I27292<= not (WX8275 and I27290);
	I27303<= not (WX8355 and WX8277);
	I27304<= not (WX8355 and I27303);
	I27305<= not (WX8277 and I27303);
	I27316<= not (WX8356 and WX8279);
	I27317<= not (WX8356 and I27316);
	I27318<= not (WX8279 and I27316);
	I27329<= not (WX8357 and WX8281);
	I27330<= not (WX8357 and I27329);
	I27331<= not (WX8281 and I27329);
	I27342<= not (WX8358 and WX8283);
	I27343<= not (WX8358 and I27342);
	I27344<= not (WX8283 and I27342);
	I27355<= not (WX8359 and WX8285);
	I27356<= not (WX8359 and I27355);
	I27357<= not (WX8285 and I27355);
	I27368<= not (WX8360 and WX8287);
	I27369<= not (WX8360 and I27368);
	I27370<= not (WX8287 and I27368);
	I27381<= not (WX8361 and WX8289);
	I27382<= not (WX8361 and I27381);
	I27383<= not (WX8289 and I27381);
	I27394<= not (WX8362 and WX8291);
	I27395<= not (WX8362 and I27394);
	I27396<= not (WX8291 and I27394);
	I27407<= not (WX8363 and WX8293);
	I27408<= not (WX8363 and I27407);
	I27409<= not (WX8293 and I27407);
	I27420<= not (WX8364 and WX8295);
	I27421<= not (WX8364 and I27420);
	I27422<= not (WX8295 and I27420);
	I27433<= not (WX8365 and WX8297);
	I27434<= not (WX8365 and I27433);
	I27435<= not (WX8297 and I27433);
	I27446<= not (WX8366 and WX8299);
	I27447<= not (WX8366 and I27446);
	I27448<= not (WX8299 and I27446);
	I27459<= not (WX8367 and WX8301);
	I27460<= not (WX8367 and I27459);
	I27461<= not (WX8301 and I27459);
	I27472<= not (WX8368 and WX8303);
	I27473<= not (WX8368 and I27472);
	I27474<= not (WX8303 and I27472);
	I27485<= not (WX8369 and WX8305);
	I27486<= not (WX8369 and I27485);
	I27487<= not (WX8305 and I27485);
	I27499<= not (I27501 and I27502);
	I27500<= not (WX8385 and CRC_OUT_3_31);
	I27501<= not (WX8385 and I27500);
	I27502<= not (CRC_OUT_3_31 and I27500);
	I27507<= not (CRC_OUT_3_15 and I27499);
	I27508<= not (CRC_OUT_3_15 and I27507);
	I27509<= not (I27499 and I27507);
	I27514<= not (I27516 and I27517);
	I27515<= not (WX8390 and CRC_OUT_3_31);
	I27516<= not (WX8390 and I27515);
	I27517<= not (CRC_OUT_3_31 and I27515);
	I27522<= not (CRC_OUT_3_10 and I27514);
	I27523<= not (CRC_OUT_3_10 and I27522);
	I27524<= not (I27514 and I27522);
	I27529<= not (I27531 and I27532);
	I27530<= not (WX8397 and CRC_OUT_3_31);
	I27531<= not (WX8397 and I27530);
	I27532<= not (CRC_OUT_3_31 and I27530);
	I27537<= not (CRC_OUT_3_3 and I27529);
	I27538<= not (CRC_OUT_3_3 and I27537);
	I27539<= not (I27529 and I27537);
	I27544<= not (WX8401 and CRC_OUT_3_31);
	I27545<= not (WX8401 and I27544);
	I27546<= not (CRC_OUT_3_31 and I27544);
	I27551<= not (WX8370 and CRC_OUT_3_30);
	I27552<= not (WX8370 and I27551);
	I27553<= not (CRC_OUT_3_30 and I27551);
	I27558<= not (WX8371 and CRC_OUT_3_29);
	I27559<= not (WX8371 and I27558);
	I27560<= not (CRC_OUT_3_29 and I27558);
	I27565<= not (WX8372 and CRC_OUT_3_28);
	I27566<= not (WX8372 and I27565);
	I27567<= not (CRC_OUT_3_28 and I27565);
	I27572<= not (WX8373 and CRC_OUT_3_27);
	I27573<= not (WX8373 and I27572);
	I27574<= not (CRC_OUT_3_27 and I27572);
	I27579<= not (WX8374 and CRC_OUT_3_26);
	I27580<= not (WX8374 and I27579);
	I27581<= not (CRC_OUT_3_26 and I27579);
	I27586<= not (WX8375 and CRC_OUT_3_25);
	I27587<= not (WX8375 and I27586);
	I27588<= not (CRC_OUT_3_25 and I27586);
	I27593<= not (WX8376 and CRC_OUT_3_24);
	I27594<= not (WX8376 and I27593);
	I27595<= not (CRC_OUT_3_24 and I27593);
	I27600<= not (WX8377 and CRC_OUT_3_23);
	I27601<= not (WX8377 and I27600);
	I27602<= not (CRC_OUT_3_23 and I27600);
	I27607<= not (WX8378 and CRC_OUT_3_22);
	I27608<= not (WX8378 and I27607);
	I27609<= not (CRC_OUT_3_22 and I27607);
	I27614<= not (WX8379 and CRC_OUT_3_21);
	I27615<= not (WX8379 and I27614);
	I27616<= not (CRC_OUT_3_21 and I27614);
	I27621<= not (WX8380 and CRC_OUT_3_20);
	I27622<= not (WX8380 and I27621);
	I27623<= not (CRC_OUT_3_20 and I27621);
	I27628<= not (WX8381 and CRC_OUT_3_19);
	I27629<= not (WX8381 and I27628);
	I27630<= not (CRC_OUT_3_19 and I27628);
	I27635<= not (WX8382 and CRC_OUT_3_18);
	I27636<= not (WX8382 and I27635);
	I27637<= not (CRC_OUT_3_18 and I27635);
	I27642<= not (WX8383 and CRC_OUT_3_17);
	I27643<= not (WX8383 and I27642);
	I27644<= not (CRC_OUT_3_17 and I27642);
	I27649<= not (WX8384 and CRC_OUT_3_16);
	I27650<= not (WX8384 and I27649);
	I27651<= not (CRC_OUT_3_16 and I27649);
	I27656<= not (WX8386 and CRC_OUT_3_14);
	I27657<= not (WX8386 and I27656);
	I27658<= not (CRC_OUT_3_14 and I27656);
	I27663<= not (WX8387 and CRC_OUT_3_13);
	I27664<= not (WX8387 and I27663);
	I27665<= not (CRC_OUT_3_13 and I27663);
	I27670<= not (WX8388 and CRC_OUT_3_12);
	I27671<= not (WX8388 and I27670);
	I27672<= not (CRC_OUT_3_12 and I27670);
	I27677<= not (WX8389 and CRC_OUT_3_11);
	I27678<= not (WX8389 and I27677);
	I27679<= not (CRC_OUT_3_11 and I27677);
	I27684<= not (WX8391 and CRC_OUT_3_9);
	I27685<= not (WX8391 and I27684);
	I27686<= not (CRC_OUT_3_9 and I27684);
	I27691<= not (WX8392 and CRC_OUT_3_8);
	I27692<= not (WX8392 and I27691);
	I27693<= not (CRC_OUT_3_8 and I27691);
	I27698<= not (WX8393 and CRC_OUT_3_7);
	I27699<= not (WX8393 and I27698);
	I27700<= not (CRC_OUT_3_7 and I27698);
	I27705<= not (WX8394 and CRC_OUT_3_6);
	I27706<= not (WX8394 and I27705);
	I27707<= not (CRC_OUT_3_6 and I27705);
	I27712<= not (WX8395 and CRC_OUT_3_5);
	I27713<= not (WX8395 and I27712);
	I27714<= not (CRC_OUT_3_5 and I27712);
	I27719<= not (WX8396 and CRC_OUT_3_4);
	I27720<= not (WX8396 and I27719);
	I27721<= not (CRC_OUT_3_4 and I27719);
	I27726<= not (WX8398 and CRC_OUT_3_2);
	I27727<= not (WX8398 and I27726);
	I27728<= not (CRC_OUT_3_2 and I27726);
	I27733<= not (WX8399 and CRC_OUT_3_1);
	I27734<= not (WX8399 and I27733);
	I27735<= not (CRC_OUT_3_1 and I27733);
	I27740<= not (WX8400 and CRC_OUT_3_0);
	I27741<= not (WX8400 and I27740);
	I27742<= not (CRC_OUT_3_0 and I27740);
	I30021<= not (I30031 and I30032);
	I30022<= not (I30024 and I30025);
	I30023<= not (WX10052 and WX9696);
	I30024<= not (WX10052 and I30023);
	I30025<= not (WX9696 and I30023);
	I30030<= not (WX9760 and I30022);
	I30031<= not (WX9760 and I30030);
	I30032<= not (I30022 and I30030);
	I30037<= not (I30039 and I30040);
	I30038<= not (WX9824 and WX9888);
	I30039<= not (WX9824 and I30038);
	I30040<= not (WX9888 and I30038);
	I30045<= not (I30021 and I30037);
	I30046<= not (I30021 and I30045);
	I30047<= not (I30037 and I30045);
	I30052<= not (I30062 and I30063);
	I30053<= not (I30055 and I30056);
	I30054<= not (WX10052 and WX9698);
	I30055<= not (WX10052 and I30054);
	I30056<= not (WX9698 and I30054);
	I30061<= not (WX9762 and I30053);
	I30062<= not (WX9762 and I30061);
	I30063<= not (I30053 and I30061);
	I30068<= not (I30070 and I30071);
	I30069<= not (WX9826 and WX9890);
	I30070<= not (WX9826 and I30069);
	I30071<= not (WX9890 and I30069);
	I30076<= not (I30052 and I30068);
	I30077<= not (I30052 and I30076);
	I30078<= not (I30068 and I30076);
	I30083<= not (I30093 and I30094);
	I30084<= not (I30086 and I30087);
	I30085<= not (WX10052 and WX9700);
	I30086<= not (WX10052 and I30085);
	I30087<= not (WX9700 and I30085);
	I30092<= not (WX9764 and I30084);
	I30093<= not (WX9764 and I30092);
	I30094<= not (I30084 and I30092);
	I30099<= not (I30101 and I30102);
	I30100<= not (WX9828 and WX9892);
	I30101<= not (WX9828 and I30100);
	I30102<= not (WX9892 and I30100);
	I30107<= not (I30083 and I30099);
	I30108<= not (I30083 and I30107);
	I30109<= not (I30099 and I30107);
	I30114<= not (I30124 and I30125);
	I30115<= not (I30117 and I30118);
	I30116<= not (WX10052 and WX9702);
	I30117<= not (WX10052 and I30116);
	I30118<= not (WX9702 and I30116);
	I30123<= not (WX9766 and I30115);
	I30124<= not (WX9766 and I30123);
	I30125<= not (I30115 and I30123);
	I30130<= not (I30132 and I30133);
	I30131<= not (WX9830 and WX9894);
	I30132<= not (WX9830 and I30131);
	I30133<= not (WX9894 and I30131);
	I30138<= not (I30114 and I30130);
	I30139<= not (I30114 and I30138);
	I30140<= not (I30130 and I30138);
	I30145<= not (I30155 and I30156);
	I30146<= not (I30148 and I30149);
	I30147<= not (WX10052 and WX9704);
	I30148<= not (WX10052 and I30147);
	I30149<= not (WX9704 and I30147);
	I30154<= not (WX9768 and I30146);
	I30155<= not (WX9768 and I30154);
	I30156<= not (I30146 and I30154);
	I30161<= not (I30163 and I30164);
	I30162<= not (WX9832 and WX9896);
	I30163<= not (WX9832 and I30162);
	I30164<= not (WX9896 and I30162);
	I30169<= not (I30145 and I30161);
	I30170<= not (I30145 and I30169);
	I30171<= not (I30161 and I30169);
	I30176<= not (I30186 and I30187);
	I30177<= not (I30179 and I30180);
	I30178<= not (WX10052 and WX9706);
	I30179<= not (WX10052 and I30178);
	I30180<= not (WX9706 and I30178);
	I30185<= not (WX9770 and I30177);
	I30186<= not (WX9770 and I30185);
	I30187<= not (I30177 and I30185);
	I30192<= not (I30194 and I30195);
	I30193<= not (WX9834 and WX9898);
	I30194<= not (WX9834 and I30193);
	I30195<= not (WX9898 and I30193);
	I30200<= not (I30176 and I30192);
	I30201<= not (I30176 and I30200);
	I30202<= not (I30192 and I30200);
	I30207<= not (I30217 and I30218);
	I30208<= not (I30210 and I30211);
	I30209<= not (WX10052 and WX9708);
	I30210<= not (WX10052 and I30209);
	I30211<= not (WX9708 and I30209);
	I30216<= not (WX9772 and I30208);
	I30217<= not (WX9772 and I30216);
	I30218<= not (I30208 and I30216);
	I30223<= not (I30225 and I30226);
	I30224<= not (WX9836 and WX9900);
	I30225<= not (WX9836 and I30224);
	I30226<= not (WX9900 and I30224);
	I30231<= not (I30207 and I30223);
	I30232<= not (I30207 and I30231);
	I30233<= not (I30223 and I30231);
	I30238<= not (I30248 and I30249);
	I30239<= not (I30241 and I30242);
	I30240<= not (WX10052 and WX9710);
	I30241<= not (WX10052 and I30240);
	I30242<= not (WX9710 and I30240);
	I30247<= not (WX9774 and I30239);
	I30248<= not (WX9774 and I30247);
	I30249<= not (I30239 and I30247);
	I30254<= not (I30256 and I30257);
	I30255<= not (WX9838 and WX9902);
	I30256<= not (WX9838 and I30255);
	I30257<= not (WX9902 and I30255);
	I30262<= not (I30238 and I30254);
	I30263<= not (I30238 and I30262);
	I30264<= not (I30254 and I30262);
	I30269<= not (I30279 and I30280);
	I30270<= not (I30272 and I30273);
	I30271<= not (WX10052 and WX9712);
	I30272<= not (WX10052 and I30271);
	I30273<= not (WX9712 and I30271);
	I30278<= not (WX9776 and I30270);
	I30279<= not (WX9776 and I30278);
	I30280<= not (I30270 and I30278);
	I30285<= not (I30287 and I30288);
	I30286<= not (WX9840 and WX9904);
	I30287<= not (WX9840 and I30286);
	I30288<= not (WX9904 and I30286);
	I30293<= not (I30269 and I30285);
	I30294<= not (I30269 and I30293);
	I30295<= not (I30285 and I30293);
	I30300<= not (I30310 and I30311);
	I30301<= not (I30303 and I30304);
	I30302<= not (WX10052 and WX9714);
	I30303<= not (WX10052 and I30302);
	I30304<= not (WX9714 and I30302);
	I30309<= not (WX9778 and I30301);
	I30310<= not (WX9778 and I30309);
	I30311<= not (I30301 and I30309);
	I30316<= not (I30318 and I30319);
	I30317<= not (WX9842 and WX9906);
	I30318<= not (WX9842 and I30317);
	I30319<= not (WX9906 and I30317);
	I30324<= not (I30300 and I30316);
	I30325<= not (I30300 and I30324);
	I30326<= not (I30316 and I30324);
	I30331<= not (I30341 and I30342);
	I30332<= not (I30334 and I30335);
	I30333<= not (WX10052 and WX9716);
	I30334<= not (WX10052 and I30333);
	I30335<= not (WX9716 and I30333);
	I30340<= not (WX9780 and I30332);
	I30341<= not (WX9780 and I30340);
	I30342<= not (I30332 and I30340);
	I30347<= not (I30349 and I30350);
	I30348<= not (WX9844 and WX9908);
	I30349<= not (WX9844 and I30348);
	I30350<= not (WX9908 and I30348);
	I30355<= not (I30331 and I30347);
	I30356<= not (I30331 and I30355);
	I30357<= not (I30347 and I30355);
	I30362<= not (I30372 and I30373);
	I30363<= not (I30365 and I30366);
	I30364<= not (WX10052 and WX9718);
	I30365<= not (WX10052 and I30364);
	I30366<= not (WX9718 and I30364);
	I30371<= not (WX9782 and I30363);
	I30372<= not (WX9782 and I30371);
	I30373<= not (I30363 and I30371);
	I30378<= not (I30380 and I30381);
	I30379<= not (WX9846 and WX9910);
	I30380<= not (WX9846 and I30379);
	I30381<= not (WX9910 and I30379);
	I30386<= not (I30362 and I30378);
	I30387<= not (I30362 and I30386);
	I30388<= not (I30378 and I30386);
	I30393<= not (I30403 and I30404);
	I30394<= not (I30396 and I30397);
	I30395<= not (WX10052 and WX9720);
	I30396<= not (WX10052 and I30395);
	I30397<= not (WX9720 and I30395);
	I30402<= not (WX9784 and I30394);
	I30403<= not (WX9784 and I30402);
	I30404<= not (I30394 and I30402);
	I30409<= not (I30411 and I30412);
	I30410<= not (WX9848 and WX9912);
	I30411<= not (WX9848 and I30410);
	I30412<= not (WX9912 and I30410);
	I30417<= not (I30393 and I30409);
	I30418<= not (I30393 and I30417);
	I30419<= not (I30409 and I30417);
	I30424<= not (I30434 and I30435);
	I30425<= not (I30427 and I30428);
	I30426<= not (WX10052 and WX9722);
	I30427<= not (WX10052 and I30426);
	I30428<= not (WX9722 and I30426);
	I30433<= not (WX9786 and I30425);
	I30434<= not (WX9786 and I30433);
	I30435<= not (I30425 and I30433);
	I30440<= not (I30442 and I30443);
	I30441<= not (WX9850 and WX9914);
	I30442<= not (WX9850 and I30441);
	I30443<= not (WX9914 and I30441);
	I30448<= not (I30424 and I30440);
	I30449<= not (I30424 and I30448);
	I30450<= not (I30440 and I30448);
	I30455<= not (I30465 and I30466);
	I30456<= not (I30458 and I30459);
	I30457<= not (WX10052 and WX9724);
	I30458<= not (WX10052 and I30457);
	I30459<= not (WX9724 and I30457);
	I30464<= not (WX9788 and I30456);
	I30465<= not (WX9788 and I30464);
	I30466<= not (I30456 and I30464);
	I30471<= not (I30473 and I30474);
	I30472<= not (WX9852 and WX9916);
	I30473<= not (WX9852 and I30472);
	I30474<= not (WX9916 and I30472);
	I30479<= not (I30455 and I30471);
	I30480<= not (I30455 and I30479);
	I30481<= not (I30471 and I30479);
	I30486<= not (I30496 and I30497);
	I30487<= not (I30489 and I30490);
	I30488<= not (WX10052 and WX9726);
	I30489<= not (WX10052 and I30488);
	I30490<= not (WX9726 and I30488);
	I30495<= not (WX9790 and I30487);
	I30496<= not (WX9790 and I30495);
	I30497<= not (I30487 and I30495);
	I30502<= not (I30504 and I30505);
	I30503<= not (WX9854 and WX9918);
	I30504<= not (WX9854 and I30503);
	I30505<= not (WX9918 and I30503);
	I30510<= not (I30486 and I30502);
	I30511<= not (I30486 and I30510);
	I30512<= not (I30502 and I30510);
	I30517<= not (I30527 and I30528);
	I30518<= not (I30520 and I30521);
	I30519<= not (WX10053 and WX9728);
	I30520<= not (WX10053 and I30519);
	I30521<= not (WX9728 and I30519);
	I30526<= not (WX9792 and I30518);
	I30527<= not (WX9792 and I30526);
	I30528<= not (I30518 and I30526);
	I30533<= not (I30535 and I30536);
	I30534<= not (WX9856 and WX9920);
	I30535<= not (WX9856 and I30534);
	I30536<= not (WX9920 and I30534);
	I30541<= not (I30517 and I30533);
	I30542<= not (I30517 and I30541);
	I30543<= not (I30533 and I30541);
	I30548<= not (I30558 and I30559);
	I30549<= not (I30551 and I30552);
	I30550<= not (WX10053 and WX9730);
	I30551<= not (WX10053 and I30550);
	I30552<= not (WX9730 and I30550);
	I30557<= not (WX9794 and I30549);
	I30558<= not (WX9794 and I30557);
	I30559<= not (I30549 and I30557);
	I30564<= not (I30566 and I30567);
	I30565<= not (WX9858 and WX9922);
	I30566<= not (WX9858 and I30565);
	I30567<= not (WX9922 and I30565);
	I30572<= not (I30548 and I30564);
	I30573<= not (I30548 and I30572);
	I30574<= not (I30564 and I30572);
	I30579<= not (I30589 and I30590);
	I30580<= not (I30582 and I30583);
	I30581<= not (WX10053 and WX9732);
	I30582<= not (WX10053 and I30581);
	I30583<= not (WX9732 and I30581);
	I30588<= not (WX9796 and I30580);
	I30589<= not (WX9796 and I30588);
	I30590<= not (I30580 and I30588);
	I30595<= not (I30597 and I30598);
	I30596<= not (WX9860 and WX9924);
	I30597<= not (WX9860 and I30596);
	I30598<= not (WX9924 and I30596);
	I30603<= not (I30579 and I30595);
	I30604<= not (I30579 and I30603);
	I30605<= not (I30595 and I30603);
	I30610<= not (I30620 and I30621);
	I30611<= not (I30613 and I30614);
	I30612<= not (WX10053 and WX9734);
	I30613<= not (WX10053 and I30612);
	I30614<= not (WX9734 and I30612);
	I30619<= not (WX9798 and I30611);
	I30620<= not (WX9798 and I30619);
	I30621<= not (I30611 and I30619);
	I30626<= not (I30628 and I30629);
	I30627<= not (WX9862 and WX9926);
	I30628<= not (WX9862 and I30627);
	I30629<= not (WX9926 and I30627);
	I30634<= not (I30610 and I30626);
	I30635<= not (I30610 and I30634);
	I30636<= not (I30626 and I30634);
	I30641<= not (I30651 and I30652);
	I30642<= not (I30644 and I30645);
	I30643<= not (WX10053 and WX9736);
	I30644<= not (WX10053 and I30643);
	I30645<= not (WX9736 and I30643);
	I30650<= not (WX9800 and I30642);
	I30651<= not (WX9800 and I30650);
	I30652<= not (I30642 and I30650);
	I30657<= not (I30659 and I30660);
	I30658<= not (WX9864 and WX9928);
	I30659<= not (WX9864 and I30658);
	I30660<= not (WX9928 and I30658);
	I30665<= not (I30641 and I30657);
	I30666<= not (I30641 and I30665);
	I30667<= not (I30657 and I30665);
	I30672<= not (I30682 and I30683);
	I30673<= not (I30675 and I30676);
	I30674<= not (WX10053 and WX9738);
	I30675<= not (WX10053 and I30674);
	I30676<= not (WX9738 and I30674);
	I30681<= not (WX9802 and I30673);
	I30682<= not (WX9802 and I30681);
	I30683<= not (I30673 and I30681);
	I30688<= not (I30690 and I30691);
	I30689<= not (WX9866 and WX9930);
	I30690<= not (WX9866 and I30689);
	I30691<= not (WX9930 and I30689);
	I30696<= not (I30672 and I30688);
	I30697<= not (I30672 and I30696);
	I30698<= not (I30688 and I30696);
	I30703<= not (I30713 and I30714);
	I30704<= not (I30706 and I30707);
	I30705<= not (WX10053 and WX9740);
	I30706<= not (WX10053 and I30705);
	I30707<= not (WX9740 and I30705);
	I30712<= not (WX9804 and I30704);
	I30713<= not (WX9804 and I30712);
	I30714<= not (I30704 and I30712);
	I30719<= not (I30721 and I30722);
	I30720<= not (WX9868 and WX9932);
	I30721<= not (WX9868 and I30720);
	I30722<= not (WX9932 and I30720);
	I30727<= not (I30703 and I30719);
	I30728<= not (I30703 and I30727);
	I30729<= not (I30719 and I30727);
	I30734<= not (I30744 and I30745);
	I30735<= not (I30737 and I30738);
	I30736<= not (WX10053 and WX9742);
	I30737<= not (WX10053 and I30736);
	I30738<= not (WX9742 and I30736);
	I30743<= not (WX9806 and I30735);
	I30744<= not (WX9806 and I30743);
	I30745<= not (I30735 and I30743);
	I30750<= not (I30752 and I30753);
	I30751<= not (WX9870 and WX9934);
	I30752<= not (WX9870 and I30751);
	I30753<= not (WX9934 and I30751);
	I30758<= not (I30734 and I30750);
	I30759<= not (I30734 and I30758);
	I30760<= not (I30750 and I30758);
	I30765<= not (I30775 and I30776);
	I30766<= not (I30768 and I30769);
	I30767<= not (WX10053 and WX9744);
	I30768<= not (WX10053 and I30767);
	I30769<= not (WX9744 and I30767);
	I30774<= not (WX9808 and I30766);
	I30775<= not (WX9808 and I30774);
	I30776<= not (I30766 and I30774);
	I30781<= not (I30783 and I30784);
	I30782<= not (WX9872 and WX9936);
	I30783<= not (WX9872 and I30782);
	I30784<= not (WX9936 and I30782);
	I30789<= not (I30765 and I30781);
	I30790<= not (I30765 and I30789);
	I30791<= not (I30781 and I30789);
	I30796<= not (I30806 and I30807);
	I30797<= not (I30799 and I30800);
	I30798<= not (WX10053 and WX9746);
	I30799<= not (WX10053 and I30798);
	I30800<= not (WX9746 and I30798);
	I30805<= not (WX9810 and I30797);
	I30806<= not (WX9810 and I30805);
	I30807<= not (I30797 and I30805);
	I30812<= not (I30814 and I30815);
	I30813<= not (WX9874 and WX9938);
	I30814<= not (WX9874 and I30813);
	I30815<= not (WX9938 and I30813);
	I30820<= not (I30796 and I30812);
	I30821<= not (I30796 and I30820);
	I30822<= not (I30812 and I30820);
	I30827<= not (I30837 and I30838);
	I30828<= not (I30830 and I30831);
	I30829<= not (WX10053 and WX9748);
	I30830<= not (WX10053 and I30829);
	I30831<= not (WX9748 and I30829);
	I30836<= not (WX9812 and I30828);
	I30837<= not (WX9812 and I30836);
	I30838<= not (I30828 and I30836);
	I30843<= not (I30845 and I30846);
	I30844<= not (WX9876 and WX9940);
	I30845<= not (WX9876 and I30844);
	I30846<= not (WX9940 and I30844);
	I30851<= not (I30827 and I30843);
	I30852<= not (I30827 and I30851);
	I30853<= not (I30843 and I30851);
	I30858<= not (I30868 and I30869);
	I30859<= not (I30861 and I30862);
	I30860<= not (WX10053 and WX9750);
	I30861<= not (WX10053 and I30860);
	I30862<= not (WX9750 and I30860);
	I30867<= not (WX9814 and I30859);
	I30868<= not (WX9814 and I30867);
	I30869<= not (I30859 and I30867);
	I30874<= not (I30876 and I30877);
	I30875<= not (WX9878 and WX9942);
	I30876<= not (WX9878 and I30875);
	I30877<= not (WX9942 and I30875);
	I30882<= not (I30858 and I30874);
	I30883<= not (I30858 and I30882);
	I30884<= not (I30874 and I30882);
	I30889<= not (I30899 and I30900);
	I30890<= not (I30892 and I30893);
	I30891<= not (WX10053 and WX9752);
	I30892<= not (WX10053 and I30891);
	I30893<= not (WX9752 and I30891);
	I30898<= not (WX9816 and I30890);
	I30899<= not (WX9816 and I30898);
	I30900<= not (I30890 and I30898);
	I30905<= not (I30907 and I30908);
	I30906<= not (WX9880 and WX9944);
	I30907<= not (WX9880 and I30906);
	I30908<= not (WX9944 and I30906);
	I30913<= not (I30889 and I30905);
	I30914<= not (I30889 and I30913);
	I30915<= not (I30905 and I30913);
	I30920<= not (I30930 and I30931);
	I30921<= not (I30923 and I30924);
	I30922<= not (WX10053 and WX9754);
	I30923<= not (WX10053 and I30922);
	I30924<= not (WX9754 and I30922);
	I30929<= not (WX9818 and I30921);
	I30930<= not (WX9818 and I30929);
	I30931<= not (I30921 and I30929);
	I30936<= not (I30938 and I30939);
	I30937<= not (WX9882 and WX9946);
	I30938<= not (WX9882 and I30937);
	I30939<= not (WX9946 and I30937);
	I30944<= not (I30920 and I30936);
	I30945<= not (I30920 and I30944);
	I30946<= not (I30936 and I30944);
	I30951<= not (I30961 and I30962);
	I30952<= not (I30954 and I30955);
	I30953<= not (WX10053 and WX9756);
	I30954<= not (WX10053 and I30953);
	I30955<= not (WX9756 and I30953);
	I30960<= not (WX9820 and I30952);
	I30961<= not (WX9820 and I30960);
	I30962<= not (I30952 and I30960);
	I30967<= not (I30969 and I30970);
	I30968<= not (WX9884 and WX9948);
	I30969<= not (WX9884 and I30968);
	I30970<= not (WX9948 and I30968);
	I30975<= not (I30951 and I30967);
	I30976<= not (I30951 and I30975);
	I30977<= not (I30967 and I30975);
	I30982<= not (I30992 and I30993);
	I30983<= not (I30985 and I30986);
	I30984<= not (WX10053 and WX9758);
	I30985<= not (WX10053 and I30984);
	I30986<= not (WX9758 and I30984);
	I30991<= not (WX9822 and I30983);
	I30992<= not (WX9822 and I30991);
	I30993<= not (I30983 and I30991);
	I30998<= not (I31000 and I31001);
	I30999<= not (WX9886 and WX9950);
	I31000<= not (WX9886 and I30999);
	I31001<= not (WX9950 and I30999);
	I31006<= not (I30982 and I30998);
	I31007<= not (I30982 and I31006);
	I31008<= not (I30998 and I31006);
	I31087<= not (WX9631 and WX9536);
	I31088<= not (WX9631 and I31087);
	I31089<= not (WX9536 and I31087);
	I31100<= not (WX9632 and WX9538);
	I31101<= not (WX9632 and I31100);
	I31102<= not (WX9538 and I31100);
	I31113<= not (WX9633 and WX9540);
	I31114<= not (WX9633 and I31113);
	I31115<= not (WX9540 and I31113);
	I31126<= not (WX9634 and WX9542);
	I31127<= not (WX9634 and I31126);
	I31128<= not (WX9542 and I31126);
	I31139<= not (WX9635 and WX9544);
	I31140<= not (WX9635 and I31139);
	I31141<= not (WX9544 and I31139);
	I31152<= not (WX9636 and WX9546);
	I31153<= not (WX9636 and I31152);
	I31154<= not (WX9546 and I31152);
	I31165<= not (WX9637 and WX9548);
	I31166<= not (WX9637 and I31165);
	I31167<= not (WX9548 and I31165);
	I31178<= not (WX9638 and WX9550);
	I31179<= not (WX9638 and I31178);
	I31180<= not (WX9550 and I31178);
	I31191<= not (WX9639 and WX9552);
	I31192<= not (WX9639 and I31191);
	I31193<= not (WX9552 and I31191);
	I31204<= not (WX9640 and WX9554);
	I31205<= not (WX9640 and I31204);
	I31206<= not (WX9554 and I31204);
	I31217<= not (WX9641 and WX9556);
	I31218<= not (WX9641 and I31217);
	I31219<= not (WX9556 and I31217);
	I31230<= not (WX9642 and WX9558);
	I31231<= not (WX9642 and I31230);
	I31232<= not (WX9558 and I31230);
	I31243<= not (WX9643 and WX9560);
	I31244<= not (WX9643 and I31243);
	I31245<= not (WX9560 and I31243);
	I31256<= not (WX9644 and WX9562);
	I31257<= not (WX9644 and I31256);
	I31258<= not (WX9562 and I31256);
	I31269<= not (WX9645 and WX9564);
	I31270<= not (WX9645 and I31269);
	I31271<= not (WX9564 and I31269);
	I31282<= not (WX9646 and WX9566);
	I31283<= not (WX9646 and I31282);
	I31284<= not (WX9566 and I31282);
	I31295<= not (WX9647 and WX9568);
	I31296<= not (WX9647 and I31295);
	I31297<= not (WX9568 and I31295);
	I31308<= not (WX9648 and WX9570);
	I31309<= not (WX9648 and I31308);
	I31310<= not (WX9570 and I31308);
	I31321<= not (WX9649 and WX9572);
	I31322<= not (WX9649 and I31321);
	I31323<= not (WX9572 and I31321);
	I31334<= not (WX9650 and WX9574);
	I31335<= not (WX9650 and I31334);
	I31336<= not (WX9574 and I31334);
	I31347<= not (WX9651 and WX9576);
	I31348<= not (WX9651 and I31347);
	I31349<= not (WX9576 and I31347);
	I31360<= not (WX9652 and WX9578);
	I31361<= not (WX9652 and I31360);
	I31362<= not (WX9578 and I31360);
	I31373<= not (WX9653 and WX9580);
	I31374<= not (WX9653 and I31373);
	I31375<= not (WX9580 and I31373);
	I31386<= not (WX9654 and WX9582);
	I31387<= not (WX9654 and I31386);
	I31388<= not (WX9582 and I31386);
	I31399<= not (WX9655 and WX9584);
	I31400<= not (WX9655 and I31399);
	I31401<= not (WX9584 and I31399);
	I31412<= not (WX9656 and WX9586);
	I31413<= not (WX9656 and I31412);
	I31414<= not (WX9586 and I31412);
	I31425<= not (WX9657 and WX9588);
	I31426<= not (WX9657 and I31425);
	I31427<= not (WX9588 and I31425);
	I31438<= not (WX9658 and WX9590);
	I31439<= not (WX9658 and I31438);
	I31440<= not (WX9590 and I31438);
	I31451<= not (WX9659 and WX9592);
	I31452<= not (WX9659 and I31451);
	I31453<= not (WX9592 and I31451);
	I31464<= not (WX9660 and WX9594);
	I31465<= not (WX9660 and I31464);
	I31466<= not (WX9594 and I31464);
	I31477<= not (WX9661 and WX9596);
	I31478<= not (WX9661 and I31477);
	I31479<= not (WX9596 and I31477);
	I31490<= not (WX9662 and WX9598);
	I31491<= not (WX9662 and I31490);
	I31492<= not (WX9598 and I31490);
	I31504<= not (I31506 and I31507);
	I31505<= not (WX9678 and CRC_OUT_2_31);
	I31506<= not (WX9678 and I31505);
	I31507<= not (CRC_OUT_2_31 and I31505);
	I31512<= not (CRC_OUT_2_15 and I31504);
	I31513<= not (CRC_OUT_2_15 and I31512);
	I31514<= not (I31504 and I31512);
	I31519<= not (I31521 and I31522);
	I31520<= not (WX9683 and CRC_OUT_2_31);
	I31521<= not (WX9683 and I31520);
	I31522<= not (CRC_OUT_2_31 and I31520);
	I31527<= not (CRC_OUT_2_10 and I31519);
	I31528<= not (CRC_OUT_2_10 and I31527);
	I31529<= not (I31519 and I31527);
	I31534<= not (I31536 and I31537);
	I31535<= not (WX9690 and CRC_OUT_2_31);
	I31536<= not (WX9690 and I31535);
	I31537<= not (CRC_OUT_2_31 and I31535);
	I31542<= not (CRC_OUT_2_3 and I31534);
	I31543<= not (CRC_OUT_2_3 and I31542);
	I31544<= not (I31534 and I31542);
	I31549<= not (WX9694 and CRC_OUT_2_31);
	I31550<= not (WX9694 and I31549);
	I31551<= not (CRC_OUT_2_31 and I31549);
	I31556<= not (WX9663 and CRC_OUT_2_30);
	I31557<= not (WX9663 and I31556);
	I31558<= not (CRC_OUT_2_30 and I31556);
	I31563<= not (WX9664 and CRC_OUT_2_29);
	I31564<= not (WX9664 and I31563);
	I31565<= not (CRC_OUT_2_29 and I31563);
	I31570<= not (WX9665 and CRC_OUT_2_28);
	I31571<= not (WX9665 and I31570);
	I31572<= not (CRC_OUT_2_28 and I31570);
	I31577<= not (WX9666 and CRC_OUT_2_27);
	I31578<= not (WX9666 and I31577);
	I31579<= not (CRC_OUT_2_27 and I31577);
	I31584<= not (WX9667 and CRC_OUT_2_26);
	I31585<= not (WX9667 and I31584);
	I31586<= not (CRC_OUT_2_26 and I31584);
	I31591<= not (WX9668 and CRC_OUT_2_25);
	I31592<= not (WX9668 and I31591);
	I31593<= not (CRC_OUT_2_25 and I31591);
	I31598<= not (WX9669 and CRC_OUT_2_24);
	I31599<= not (WX9669 and I31598);
	I31600<= not (CRC_OUT_2_24 and I31598);
	I31605<= not (WX9670 and CRC_OUT_2_23);
	I31606<= not (WX9670 and I31605);
	I31607<= not (CRC_OUT_2_23 and I31605);
	I31612<= not (WX9671 and CRC_OUT_2_22);
	I31613<= not (WX9671 and I31612);
	I31614<= not (CRC_OUT_2_22 and I31612);
	I31619<= not (WX9672 and CRC_OUT_2_21);
	I31620<= not (WX9672 and I31619);
	I31621<= not (CRC_OUT_2_21 and I31619);
	I31626<= not (WX9673 and CRC_OUT_2_20);
	I31627<= not (WX9673 and I31626);
	I31628<= not (CRC_OUT_2_20 and I31626);
	I31633<= not (WX9674 and CRC_OUT_2_19);
	I31634<= not (WX9674 and I31633);
	I31635<= not (CRC_OUT_2_19 and I31633);
	I31640<= not (WX9675 and CRC_OUT_2_18);
	I31641<= not (WX9675 and I31640);
	I31642<= not (CRC_OUT_2_18 and I31640);
	I31647<= not (WX9676 and CRC_OUT_2_17);
	I31648<= not (WX9676 and I31647);
	I31649<= not (CRC_OUT_2_17 and I31647);
	I31654<= not (WX9677 and CRC_OUT_2_16);
	I31655<= not (WX9677 and I31654);
	I31656<= not (CRC_OUT_2_16 and I31654);
	I31661<= not (WX9679 and CRC_OUT_2_14);
	I31662<= not (WX9679 and I31661);
	I31663<= not (CRC_OUT_2_14 and I31661);
	I31668<= not (WX9680 and CRC_OUT_2_13);
	I31669<= not (WX9680 and I31668);
	I31670<= not (CRC_OUT_2_13 and I31668);
	I31675<= not (WX9681 and CRC_OUT_2_12);
	I31676<= not (WX9681 and I31675);
	I31677<= not (CRC_OUT_2_12 and I31675);
	I31682<= not (WX9682 and CRC_OUT_2_11);
	I31683<= not (WX9682 and I31682);
	I31684<= not (CRC_OUT_2_11 and I31682);
	I31689<= not (WX9684 and CRC_OUT_2_9);
	I31690<= not (WX9684 and I31689);
	I31691<= not (CRC_OUT_2_9 and I31689);
	I31696<= not (WX9685 and CRC_OUT_2_8);
	I31697<= not (WX9685 and I31696);
	I31698<= not (CRC_OUT_2_8 and I31696);
	I31703<= not (WX9686 and CRC_OUT_2_7);
	I31704<= not (WX9686 and I31703);
	I31705<= not (CRC_OUT_2_7 and I31703);
	I31710<= not (WX9687 and CRC_OUT_2_6);
	I31711<= not (WX9687 and I31710);
	I31712<= not (CRC_OUT_2_6 and I31710);
	I31717<= not (WX9688 and CRC_OUT_2_5);
	I31718<= not (WX9688 and I31717);
	I31719<= not (CRC_OUT_2_5 and I31717);
	I31724<= not (WX9689 and CRC_OUT_2_4);
	I31725<= not (WX9689 and I31724);
	I31726<= not (CRC_OUT_2_4 and I31724);
	I31731<= not (WX9691 and CRC_OUT_2_2);
	I31732<= not (WX9691 and I31731);
	I31733<= not (CRC_OUT_2_2 and I31731);
	I31738<= not (WX9692 and CRC_OUT_2_1);
	I31739<= not (WX9692 and I31738);
	I31740<= not (CRC_OUT_2_1 and I31738);
	I31745<= not (WX9693 and CRC_OUT_2_0);
	I31746<= not (WX9693 and I31745);
	I31747<= not (CRC_OUT_2_0 and I31745);
	I34026<= not (I34036 and I34037);
	I34027<= not (I34029 and I34030);
	I34028<= not (WX11345 and WX10989);
	I34029<= not (WX11345 and I34028);
	I34030<= not (WX10989 and I34028);
	I34035<= not (WX11053 and I34027);
	I34036<= not (WX11053 and I34035);
	I34037<= not (I34027 and I34035);
	I34042<= not (I34044 and I34045);
	I34043<= not (WX11117 and WX11181);
	I34044<= not (WX11117 and I34043);
	I34045<= not (WX11181 and I34043);
	I34050<= not (I34026 and I34042);
	I34051<= not (I34026 and I34050);
	I34052<= not (I34042 and I34050);
	I34057<= not (I34067 and I34068);
	I34058<= not (I34060 and I34061);
	I34059<= not (WX11345 and WX10991);
	I34060<= not (WX11345 and I34059);
	I34061<= not (WX10991 and I34059);
	I34066<= not (WX11055 and I34058);
	I34067<= not (WX11055 and I34066);
	I34068<= not (I34058 and I34066);
	I34073<= not (I34075 and I34076);
	I34074<= not (WX11119 and WX11183);
	I34075<= not (WX11119 and I34074);
	I34076<= not (WX11183 and I34074);
	I34081<= not (I34057 and I34073);
	I34082<= not (I34057 and I34081);
	I34083<= not (I34073 and I34081);
	I34088<= not (I34098 and I34099);
	I34089<= not (I34091 and I34092);
	I34090<= not (WX11345 and WX10993);
	I34091<= not (WX11345 and I34090);
	I34092<= not (WX10993 and I34090);
	I34097<= not (WX11057 and I34089);
	I34098<= not (WX11057 and I34097);
	I34099<= not (I34089 and I34097);
	I34104<= not (I34106 and I34107);
	I34105<= not (WX11121 and WX11185);
	I34106<= not (WX11121 and I34105);
	I34107<= not (WX11185 and I34105);
	I34112<= not (I34088 and I34104);
	I34113<= not (I34088 and I34112);
	I34114<= not (I34104 and I34112);
	I34119<= not (I34129 and I34130);
	I34120<= not (I34122 and I34123);
	I34121<= not (WX11345 and WX10995);
	I34122<= not (WX11345 and I34121);
	I34123<= not (WX10995 and I34121);
	I34128<= not (WX11059 and I34120);
	I34129<= not (WX11059 and I34128);
	I34130<= not (I34120 and I34128);
	I34135<= not (I34137 and I34138);
	I34136<= not (WX11123 and WX11187);
	I34137<= not (WX11123 and I34136);
	I34138<= not (WX11187 and I34136);
	I34143<= not (I34119 and I34135);
	I34144<= not (I34119 and I34143);
	I34145<= not (I34135 and I34143);
	I34150<= not (I34160 and I34161);
	I34151<= not (I34153 and I34154);
	I34152<= not (WX11345 and WX10997);
	I34153<= not (WX11345 and I34152);
	I34154<= not (WX10997 and I34152);
	I34159<= not (WX11061 and I34151);
	I34160<= not (WX11061 and I34159);
	I34161<= not (I34151 and I34159);
	I34166<= not (I34168 and I34169);
	I34167<= not (WX11125 and WX11189);
	I34168<= not (WX11125 and I34167);
	I34169<= not (WX11189 and I34167);
	I34174<= not (I34150 and I34166);
	I34175<= not (I34150 and I34174);
	I34176<= not (I34166 and I34174);
	I34181<= not (I34191 and I34192);
	I34182<= not (I34184 and I34185);
	I34183<= not (WX11345 and WX10999);
	I34184<= not (WX11345 and I34183);
	I34185<= not (WX10999 and I34183);
	I34190<= not (WX11063 and I34182);
	I34191<= not (WX11063 and I34190);
	I34192<= not (I34182 and I34190);
	I34197<= not (I34199 and I34200);
	I34198<= not (WX11127 and WX11191);
	I34199<= not (WX11127 and I34198);
	I34200<= not (WX11191 and I34198);
	I34205<= not (I34181 and I34197);
	I34206<= not (I34181 and I34205);
	I34207<= not (I34197 and I34205);
	I34212<= not (I34222 and I34223);
	I34213<= not (I34215 and I34216);
	I34214<= not (WX11345 and WX11001);
	I34215<= not (WX11345 and I34214);
	I34216<= not (WX11001 and I34214);
	I34221<= not (WX11065 and I34213);
	I34222<= not (WX11065 and I34221);
	I34223<= not (I34213 and I34221);
	I34228<= not (I34230 and I34231);
	I34229<= not (WX11129 and WX11193);
	I34230<= not (WX11129 and I34229);
	I34231<= not (WX11193 and I34229);
	I34236<= not (I34212 and I34228);
	I34237<= not (I34212 and I34236);
	I34238<= not (I34228 and I34236);
	I34243<= not (I34253 and I34254);
	I34244<= not (I34246 and I34247);
	I34245<= not (WX11345 and WX11003);
	I34246<= not (WX11345 and I34245);
	I34247<= not (WX11003 and I34245);
	I34252<= not (WX11067 and I34244);
	I34253<= not (WX11067 and I34252);
	I34254<= not (I34244 and I34252);
	I34259<= not (I34261 and I34262);
	I34260<= not (WX11131 and WX11195);
	I34261<= not (WX11131 and I34260);
	I34262<= not (WX11195 and I34260);
	I34267<= not (I34243 and I34259);
	I34268<= not (I34243 and I34267);
	I34269<= not (I34259 and I34267);
	I34274<= not (I34284 and I34285);
	I34275<= not (I34277 and I34278);
	I34276<= not (WX11345 and WX11005);
	I34277<= not (WX11345 and I34276);
	I34278<= not (WX11005 and I34276);
	I34283<= not (WX11069 and I34275);
	I34284<= not (WX11069 and I34283);
	I34285<= not (I34275 and I34283);
	I34290<= not (I34292 and I34293);
	I34291<= not (WX11133 and WX11197);
	I34292<= not (WX11133 and I34291);
	I34293<= not (WX11197 and I34291);
	I34298<= not (I34274 and I34290);
	I34299<= not (I34274 and I34298);
	I34300<= not (I34290 and I34298);
	I34305<= not (I34315 and I34316);
	I34306<= not (I34308 and I34309);
	I34307<= not (WX11345 and WX11007);
	I34308<= not (WX11345 and I34307);
	I34309<= not (WX11007 and I34307);
	I34314<= not (WX11071 and I34306);
	I34315<= not (WX11071 and I34314);
	I34316<= not (I34306 and I34314);
	I34321<= not (I34323 and I34324);
	I34322<= not (WX11135 and WX11199);
	I34323<= not (WX11135 and I34322);
	I34324<= not (WX11199 and I34322);
	I34329<= not (I34305 and I34321);
	I34330<= not (I34305 and I34329);
	I34331<= not (I34321 and I34329);
	I34336<= not (I34346 and I34347);
	I34337<= not (I34339 and I34340);
	I34338<= not (WX11345 and WX11009);
	I34339<= not (WX11345 and I34338);
	I34340<= not (WX11009 and I34338);
	I34345<= not (WX11073 and I34337);
	I34346<= not (WX11073 and I34345);
	I34347<= not (I34337 and I34345);
	I34352<= not (I34354 and I34355);
	I34353<= not (WX11137 and WX11201);
	I34354<= not (WX11137 and I34353);
	I34355<= not (WX11201 and I34353);
	I34360<= not (I34336 and I34352);
	I34361<= not (I34336 and I34360);
	I34362<= not (I34352 and I34360);
	I34367<= not (I34377 and I34378);
	I34368<= not (I34370 and I34371);
	I34369<= not (WX11345 and WX11011);
	I34370<= not (WX11345 and I34369);
	I34371<= not (WX11011 and I34369);
	I34376<= not (WX11075 and I34368);
	I34377<= not (WX11075 and I34376);
	I34378<= not (I34368 and I34376);
	I34383<= not (I34385 and I34386);
	I34384<= not (WX11139 and WX11203);
	I34385<= not (WX11139 and I34384);
	I34386<= not (WX11203 and I34384);
	I34391<= not (I34367 and I34383);
	I34392<= not (I34367 and I34391);
	I34393<= not (I34383 and I34391);
	I34398<= not (I34408 and I34409);
	I34399<= not (I34401 and I34402);
	I34400<= not (WX11345 and WX11013);
	I34401<= not (WX11345 and I34400);
	I34402<= not (WX11013 and I34400);
	I34407<= not (WX11077 and I34399);
	I34408<= not (WX11077 and I34407);
	I34409<= not (I34399 and I34407);
	I34414<= not (I34416 and I34417);
	I34415<= not (WX11141 and WX11205);
	I34416<= not (WX11141 and I34415);
	I34417<= not (WX11205 and I34415);
	I34422<= not (I34398 and I34414);
	I34423<= not (I34398 and I34422);
	I34424<= not (I34414 and I34422);
	I34429<= not (I34439 and I34440);
	I34430<= not (I34432 and I34433);
	I34431<= not (WX11345 and WX11015);
	I34432<= not (WX11345 and I34431);
	I34433<= not (WX11015 and I34431);
	I34438<= not (WX11079 and I34430);
	I34439<= not (WX11079 and I34438);
	I34440<= not (I34430 and I34438);
	I34445<= not (I34447 and I34448);
	I34446<= not (WX11143 and WX11207);
	I34447<= not (WX11143 and I34446);
	I34448<= not (WX11207 and I34446);
	I34453<= not (I34429 and I34445);
	I34454<= not (I34429 and I34453);
	I34455<= not (I34445 and I34453);
	I34460<= not (I34470 and I34471);
	I34461<= not (I34463 and I34464);
	I34462<= not (WX11345 and WX11017);
	I34463<= not (WX11345 and I34462);
	I34464<= not (WX11017 and I34462);
	I34469<= not (WX11081 and I34461);
	I34470<= not (WX11081 and I34469);
	I34471<= not (I34461 and I34469);
	I34476<= not (I34478 and I34479);
	I34477<= not (WX11145 and WX11209);
	I34478<= not (WX11145 and I34477);
	I34479<= not (WX11209 and I34477);
	I34484<= not (I34460 and I34476);
	I34485<= not (I34460 and I34484);
	I34486<= not (I34476 and I34484);
	I34491<= not (I34501 and I34502);
	I34492<= not (I34494 and I34495);
	I34493<= not (WX11345 and WX11019);
	I34494<= not (WX11345 and I34493);
	I34495<= not (WX11019 and I34493);
	I34500<= not (WX11083 and I34492);
	I34501<= not (WX11083 and I34500);
	I34502<= not (I34492 and I34500);
	I34507<= not (I34509 and I34510);
	I34508<= not (WX11147 and WX11211);
	I34509<= not (WX11147 and I34508);
	I34510<= not (WX11211 and I34508);
	I34515<= not (I34491 and I34507);
	I34516<= not (I34491 and I34515);
	I34517<= not (I34507 and I34515);
	I34522<= not (I34532 and I34533);
	I34523<= not (I34525 and I34526);
	I34524<= not (WX11346 and WX11021);
	I34525<= not (WX11346 and I34524);
	I34526<= not (WX11021 and I34524);
	I34531<= not (WX11085 and I34523);
	I34532<= not (WX11085 and I34531);
	I34533<= not (I34523 and I34531);
	I34538<= not (I34540 and I34541);
	I34539<= not (WX11149 and WX11213);
	I34540<= not (WX11149 and I34539);
	I34541<= not (WX11213 and I34539);
	I34546<= not (I34522 and I34538);
	I34547<= not (I34522 and I34546);
	I34548<= not (I34538 and I34546);
	I34553<= not (I34563 and I34564);
	I34554<= not (I34556 and I34557);
	I34555<= not (WX11346 and WX11023);
	I34556<= not (WX11346 and I34555);
	I34557<= not (WX11023 and I34555);
	I34562<= not (WX11087 and I34554);
	I34563<= not (WX11087 and I34562);
	I34564<= not (I34554 and I34562);
	I34569<= not (I34571 and I34572);
	I34570<= not (WX11151 and WX11215);
	I34571<= not (WX11151 and I34570);
	I34572<= not (WX11215 and I34570);
	I34577<= not (I34553 and I34569);
	I34578<= not (I34553 and I34577);
	I34579<= not (I34569 and I34577);
	I34584<= not (I34594 and I34595);
	I34585<= not (I34587 and I34588);
	I34586<= not (WX11346 and WX11025);
	I34587<= not (WX11346 and I34586);
	I34588<= not (WX11025 and I34586);
	I34593<= not (WX11089 and I34585);
	I34594<= not (WX11089 and I34593);
	I34595<= not (I34585 and I34593);
	I34600<= not (I34602 and I34603);
	I34601<= not (WX11153 and WX11217);
	I34602<= not (WX11153 and I34601);
	I34603<= not (WX11217 and I34601);
	I34608<= not (I34584 and I34600);
	I34609<= not (I34584 and I34608);
	I34610<= not (I34600 and I34608);
	I34615<= not (I34625 and I34626);
	I34616<= not (I34618 and I34619);
	I34617<= not (WX11346 and WX11027);
	I34618<= not (WX11346 and I34617);
	I34619<= not (WX11027 and I34617);
	I34624<= not (WX11091 and I34616);
	I34625<= not (WX11091 and I34624);
	I34626<= not (I34616 and I34624);
	I34631<= not (I34633 and I34634);
	I34632<= not (WX11155 and WX11219);
	I34633<= not (WX11155 and I34632);
	I34634<= not (WX11219 and I34632);
	I34639<= not (I34615 and I34631);
	I34640<= not (I34615 and I34639);
	I34641<= not (I34631 and I34639);
	I34646<= not (I34656 and I34657);
	I34647<= not (I34649 and I34650);
	I34648<= not (WX11346 and WX11029);
	I34649<= not (WX11346 and I34648);
	I34650<= not (WX11029 and I34648);
	I34655<= not (WX11093 and I34647);
	I34656<= not (WX11093 and I34655);
	I34657<= not (I34647 and I34655);
	I34662<= not (I34664 and I34665);
	I34663<= not (WX11157 and WX11221);
	I34664<= not (WX11157 and I34663);
	I34665<= not (WX11221 and I34663);
	I34670<= not (I34646 and I34662);
	I34671<= not (I34646 and I34670);
	I34672<= not (I34662 and I34670);
	I34677<= not (I34687 and I34688);
	I34678<= not (I34680 and I34681);
	I34679<= not (WX11346 and WX11031);
	I34680<= not (WX11346 and I34679);
	I34681<= not (WX11031 and I34679);
	I34686<= not (WX11095 and I34678);
	I34687<= not (WX11095 and I34686);
	I34688<= not (I34678 and I34686);
	I34693<= not (I34695 and I34696);
	I34694<= not (WX11159 and WX11223);
	I34695<= not (WX11159 and I34694);
	I34696<= not (WX11223 and I34694);
	I34701<= not (I34677 and I34693);
	I34702<= not (I34677 and I34701);
	I34703<= not (I34693 and I34701);
	I34708<= not (I34718 and I34719);
	I34709<= not (I34711 and I34712);
	I34710<= not (WX11346 and WX11033);
	I34711<= not (WX11346 and I34710);
	I34712<= not (WX11033 and I34710);
	I34717<= not (WX11097 and I34709);
	I34718<= not (WX11097 and I34717);
	I34719<= not (I34709 and I34717);
	I34724<= not (I34726 and I34727);
	I34725<= not (WX11161 and WX11225);
	I34726<= not (WX11161 and I34725);
	I34727<= not (WX11225 and I34725);
	I34732<= not (I34708 and I34724);
	I34733<= not (I34708 and I34732);
	I34734<= not (I34724 and I34732);
	I34739<= not (I34749 and I34750);
	I34740<= not (I34742 and I34743);
	I34741<= not (WX11346 and WX11035);
	I34742<= not (WX11346 and I34741);
	I34743<= not (WX11035 and I34741);
	I34748<= not (WX11099 and I34740);
	I34749<= not (WX11099 and I34748);
	I34750<= not (I34740 and I34748);
	I34755<= not (I34757 and I34758);
	I34756<= not (WX11163 and WX11227);
	I34757<= not (WX11163 and I34756);
	I34758<= not (WX11227 and I34756);
	I34763<= not (I34739 and I34755);
	I34764<= not (I34739 and I34763);
	I34765<= not (I34755 and I34763);
	I34770<= not (I34780 and I34781);
	I34771<= not (I34773 and I34774);
	I34772<= not (WX11346 and WX11037);
	I34773<= not (WX11346 and I34772);
	I34774<= not (WX11037 and I34772);
	I34779<= not (WX11101 and I34771);
	I34780<= not (WX11101 and I34779);
	I34781<= not (I34771 and I34779);
	I34786<= not (I34788 and I34789);
	I34787<= not (WX11165 and WX11229);
	I34788<= not (WX11165 and I34787);
	I34789<= not (WX11229 and I34787);
	I34794<= not (I34770 and I34786);
	I34795<= not (I34770 and I34794);
	I34796<= not (I34786 and I34794);
	I34801<= not (I34811 and I34812);
	I34802<= not (I34804 and I34805);
	I34803<= not (WX11346 and WX11039);
	I34804<= not (WX11346 and I34803);
	I34805<= not (WX11039 and I34803);
	I34810<= not (WX11103 and I34802);
	I34811<= not (WX11103 and I34810);
	I34812<= not (I34802 and I34810);
	I34817<= not (I34819 and I34820);
	I34818<= not (WX11167 and WX11231);
	I34819<= not (WX11167 and I34818);
	I34820<= not (WX11231 and I34818);
	I34825<= not (I34801 and I34817);
	I34826<= not (I34801 and I34825);
	I34827<= not (I34817 and I34825);
	I34832<= not (I34842 and I34843);
	I34833<= not (I34835 and I34836);
	I34834<= not (WX11346 and WX11041);
	I34835<= not (WX11346 and I34834);
	I34836<= not (WX11041 and I34834);
	I34841<= not (WX11105 and I34833);
	I34842<= not (WX11105 and I34841);
	I34843<= not (I34833 and I34841);
	I34848<= not (I34850 and I34851);
	I34849<= not (WX11169 and WX11233);
	I34850<= not (WX11169 and I34849);
	I34851<= not (WX11233 and I34849);
	I34856<= not (I34832 and I34848);
	I34857<= not (I34832 and I34856);
	I34858<= not (I34848 and I34856);
	I34863<= not (I34873 and I34874);
	I34864<= not (I34866 and I34867);
	I34865<= not (WX11346 and WX11043);
	I34866<= not (WX11346 and I34865);
	I34867<= not (WX11043 and I34865);
	I34872<= not (WX11107 and I34864);
	I34873<= not (WX11107 and I34872);
	I34874<= not (I34864 and I34872);
	I34879<= not (I34881 and I34882);
	I34880<= not (WX11171 and WX11235);
	I34881<= not (WX11171 and I34880);
	I34882<= not (WX11235 and I34880);
	I34887<= not (I34863 and I34879);
	I34888<= not (I34863 and I34887);
	I34889<= not (I34879 and I34887);
	I34894<= not (I34904 and I34905);
	I34895<= not (I34897 and I34898);
	I34896<= not (WX11346 and WX11045);
	I34897<= not (WX11346 and I34896);
	I34898<= not (WX11045 and I34896);
	I34903<= not (WX11109 and I34895);
	I34904<= not (WX11109 and I34903);
	I34905<= not (I34895 and I34903);
	I34910<= not (I34912 and I34913);
	I34911<= not (WX11173 and WX11237);
	I34912<= not (WX11173 and I34911);
	I34913<= not (WX11237 and I34911);
	I34918<= not (I34894 and I34910);
	I34919<= not (I34894 and I34918);
	I34920<= not (I34910 and I34918);
	I34925<= not (I34935 and I34936);
	I34926<= not (I34928 and I34929);
	I34927<= not (WX11346 and WX11047);
	I34928<= not (WX11346 and I34927);
	I34929<= not (WX11047 and I34927);
	I34934<= not (WX11111 and I34926);
	I34935<= not (WX11111 and I34934);
	I34936<= not (I34926 and I34934);
	I34941<= not (I34943 and I34944);
	I34942<= not (WX11175 and WX11239);
	I34943<= not (WX11175 and I34942);
	I34944<= not (WX11239 and I34942);
	I34949<= not (I34925 and I34941);
	I34950<= not (I34925 and I34949);
	I34951<= not (I34941 and I34949);
	I34956<= not (I34966 and I34967);
	I34957<= not (I34959 and I34960);
	I34958<= not (WX11346 and WX11049);
	I34959<= not (WX11346 and I34958);
	I34960<= not (WX11049 and I34958);
	I34965<= not (WX11113 and I34957);
	I34966<= not (WX11113 and I34965);
	I34967<= not (I34957 and I34965);
	I34972<= not (I34974 and I34975);
	I34973<= not (WX11177 and WX11241);
	I34974<= not (WX11177 and I34973);
	I34975<= not (WX11241 and I34973);
	I34980<= not (I34956 and I34972);
	I34981<= not (I34956 and I34980);
	I34982<= not (I34972 and I34980);
	I34987<= not (I34997 and I34998);
	I34988<= not (I34990 and I34991);
	I34989<= not (WX11346 and WX11051);
	I34990<= not (WX11346 and I34989);
	I34991<= not (WX11051 and I34989);
	I34996<= not (WX11115 and I34988);
	I34997<= not (WX11115 and I34996);
	I34998<= not (I34988 and I34996);
	I35003<= not (I35005 and I35006);
	I35004<= not (WX11179 and WX11243);
	I35005<= not (WX11179 and I35004);
	I35006<= not (WX11243 and I35004);
	I35011<= not (I34987 and I35003);
	I35012<= not (I34987 and I35011);
	I35013<= not (I35003 and I35011);
	I35092<= not (WX10924 and WX10829);
	I35093<= not (WX10924 and I35092);
	I35094<= not (WX10829 and I35092);
	I35105<= not (WX10925 and WX10831);
	I35106<= not (WX10925 and I35105);
	I35107<= not (WX10831 and I35105);
	I35118<= not (WX10926 and WX10833);
	I35119<= not (WX10926 and I35118);
	I35120<= not (WX10833 and I35118);
	I35131<= not (WX10927 and WX10835);
	I35132<= not (WX10927 and I35131);
	I35133<= not (WX10835 and I35131);
	I35144<= not (WX10928 and WX10837);
	I35145<= not (WX10928 and I35144);
	I35146<= not (WX10837 and I35144);
	I35157<= not (WX10929 and WX10839);
	I35158<= not (WX10929 and I35157);
	I35159<= not (WX10839 and I35157);
	I35170<= not (WX10930 and WX10841);
	I35171<= not (WX10930 and I35170);
	I35172<= not (WX10841 and I35170);
	I35183<= not (WX10931 and WX10843);
	I35184<= not (WX10931 and I35183);
	I35185<= not (WX10843 and I35183);
	I35196<= not (WX10932 and WX10845);
	I35197<= not (WX10932 and I35196);
	I35198<= not (WX10845 and I35196);
	I35209<= not (WX10933 and WX10847);
	I35210<= not (WX10933 and I35209);
	I35211<= not (WX10847 and I35209);
	I35222<= not (WX10934 and WX10849);
	I35223<= not (WX10934 and I35222);
	I35224<= not (WX10849 and I35222);
	I35235<= not (WX10935 and WX10851);
	I35236<= not (WX10935 and I35235);
	I35237<= not (WX10851 and I35235);
	I35248<= not (WX10936 and WX10853);
	I35249<= not (WX10936 and I35248);
	I35250<= not (WX10853 and I35248);
	I35261<= not (WX10937 and WX10855);
	I35262<= not (WX10937 and I35261);
	I35263<= not (WX10855 and I35261);
	I35274<= not (WX10938 and WX10857);
	I35275<= not (WX10938 and I35274);
	I35276<= not (WX10857 and I35274);
	I35287<= not (WX10939 and WX10859);
	I35288<= not (WX10939 and I35287);
	I35289<= not (WX10859 and I35287);
	I35300<= not (WX10940 and WX10861);
	I35301<= not (WX10940 and I35300);
	I35302<= not (WX10861 and I35300);
	I35313<= not (WX10941 and WX10863);
	I35314<= not (WX10941 and I35313);
	I35315<= not (WX10863 and I35313);
	I35326<= not (WX10942 and WX10865);
	I35327<= not (WX10942 and I35326);
	I35328<= not (WX10865 and I35326);
	I35339<= not (WX10943 and WX10867);
	I35340<= not (WX10943 and I35339);
	I35341<= not (WX10867 and I35339);
	I35352<= not (WX10944 and WX10869);
	I35353<= not (WX10944 and I35352);
	I35354<= not (WX10869 and I35352);
	I35365<= not (WX10945 and WX10871);
	I35366<= not (WX10945 and I35365);
	I35367<= not (WX10871 and I35365);
	I35378<= not (WX10946 and WX10873);
	I35379<= not (WX10946 and I35378);
	I35380<= not (WX10873 and I35378);
	I35391<= not (WX10947 and WX10875);
	I35392<= not (WX10947 and I35391);
	I35393<= not (WX10875 and I35391);
	I35404<= not (WX10948 and WX10877);
	I35405<= not (WX10948 and I35404);
	I35406<= not (WX10877 and I35404);
	I35417<= not (WX10949 and WX10879);
	I35418<= not (WX10949 and I35417);
	I35419<= not (WX10879 and I35417);
	I35430<= not (WX10950 and WX10881);
	I35431<= not (WX10950 and I35430);
	I35432<= not (WX10881 and I35430);
	I35443<= not (WX10951 and WX10883);
	I35444<= not (WX10951 and I35443);
	I35445<= not (WX10883 and I35443);
	I35456<= not (WX10952 and WX10885);
	I35457<= not (WX10952 and I35456);
	I35458<= not (WX10885 and I35456);
	I35469<= not (WX10953 and WX10887);
	I35470<= not (WX10953 and I35469);
	I35471<= not (WX10887 and I35469);
	I35482<= not (WX10954 and WX10889);
	I35483<= not (WX10954 and I35482);
	I35484<= not (WX10889 and I35482);
	I35495<= not (WX10955 and WX10891);
	I35496<= not (WX10955 and I35495);
	I35497<= not (WX10891 and I35495);
	I35509<= not (I35511 and I35512);
	I35510<= not (WX10971 and CRC_OUT_1_31);
	I35511<= not (WX10971 and I35510);
	I35512<= not (CRC_OUT_1_31 and I35510);
	I35517<= not (CRC_OUT_1_15 and I35509);
	I35518<= not (CRC_OUT_1_15 and I35517);
	I35519<= not (I35509 and I35517);
	I35524<= not (I35526 and I35527);
	I35525<= not (WX10976 and CRC_OUT_1_31);
	I35526<= not (WX10976 and I35525);
	I35527<= not (CRC_OUT_1_31 and I35525);
	I35532<= not (CRC_OUT_1_10 and I35524);
	I35533<= not (CRC_OUT_1_10 and I35532);
	I35534<= not (I35524 and I35532);
	I35539<= not (I35541 and I35542);
	I35540<= not (WX10983 and CRC_OUT_1_31);
	I35541<= not (WX10983 and I35540);
	I35542<= not (CRC_OUT_1_31 and I35540);
	I35547<= not (CRC_OUT_1_3 and I35539);
	I35548<= not (CRC_OUT_1_3 and I35547);
	I35549<= not (I35539 and I35547);
	I35554<= not (WX10987 and CRC_OUT_1_31);
	I35555<= not (WX10987 and I35554);
	I35556<= not (CRC_OUT_1_31 and I35554);
	I35561<= not (WX10956 and CRC_OUT_1_30);
	I35562<= not (WX10956 and I35561);
	I35563<= not (CRC_OUT_1_30 and I35561);
	I35568<= not (WX10957 and CRC_OUT_1_29);
	I35569<= not (WX10957 and I35568);
	I35570<= not (CRC_OUT_1_29 and I35568);
	I35575<= not (WX10958 and CRC_OUT_1_28);
	I35576<= not (WX10958 and I35575);
	I35577<= not (CRC_OUT_1_28 and I35575);
	I35582<= not (WX10959 and CRC_OUT_1_27);
	I35583<= not (WX10959 and I35582);
	I35584<= not (CRC_OUT_1_27 and I35582);
	I35589<= not (WX10960 and CRC_OUT_1_26);
	I35590<= not (WX10960 and I35589);
	I35591<= not (CRC_OUT_1_26 and I35589);
	I35596<= not (WX10961 and CRC_OUT_1_25);
	I35597<= not (WX10961 and I35596);
	I35598<= not (CRC_OUT_1_25 and I35596);
	I35603<= not (WX10962 and CRC_OUT_1_24);
	I35604<= not (WX10962 and I35603);
	I35605<= not (CRC_OUT_1_24 and I35603);
	I35610<= not (WX10963 and CRC_OUT_1_23);
	I35611<= not (WX10963 and I35610);
	I35612<= not (CRC_OUT_1_23 and I35610);
	I35617<= not (WX10964 and CRC_OUT_1_22);
	I35618<= not (WX10964 and I35617);
	I35619<= not (CRC_OUT_1_22 and I35617);
	I35624<= not (WX10965 and CRC_OUT_1_21);
	I35625<= not (WX10965 and I35624);
	I35626<= not (CRC_OUT_1_21 and I35624);
	I35631<= not (WX10966 and CRC_OUT_1_20);
	I35632<= not (WX10966 and I35631);
	I35633<= not (CRC_OUT_1_20 and I35631);
	I35638<= not (WX10967 and CRC_OUT_1_19);
	I35639<= not (WX10967 and I35638);
	I35640<= not (CRC_OUT_1_19 and I35638);
	I35645<= not (WX10968 and CRC_OUT_1_18);
	I35646<= not (WX10968 and I35645);
	I35647<= not (CRC_OUT_1_18 and I35645);
	I35652<= not (WX10969 and CRC_OUT_1_17);
	I35653<= not (WX10969 and I35652);
	I35654<= not (CRC_OUT_1_17 and I35652);
	I35659<= not (WX10970 and CRC_OUT_1_16);
	I35660<= not (WX10970 and I35659);
	I35661<= not (CRC_OUT_1_16 and I35659);
	I35666<= not (WX10972 and CRC_OUT_1_14);
	I35667<= not (WX10972 and I35666);
	I35668<= not (CRC_OUT_1_14 and I35666);
	I35673<= not (WX10973 and CRC_OUT_1_13);
	I35674<= not (WX10973 and I35673);
	I35675<= not (CRC_OUT_1_13 and I35673);
	I35680<= not (WX10974 and CRC_OUT_1_12);
	I35681<= not (WX10974 and I35680);
	I35682<= not (CRC_OUT_1_12 and I35680);
	I35687<= not (WX10975 and CRC_OUT_1_11);
	I35688<= not (WX10975 and I35687);
	I35689<= not (CRC_OUT_1_11 and I35687);
	I35694<= not (WX10977 and CRC_OUT_1_9);
	I35695<= not (WX10977 and I35694);
	I35696<= not (CRC_OUT_1_9 and I35694);
	I35701<= not (WX10978 and CRC_OUT_1_8);
	I35702<= not (WX10978 and I35701);
	I35703<= not (CRC_OUT_1_8 and I35701);
	I35708<= not (WX10979 and CRC_OUT_1_7);
	I35709<= not (WX10979 and I35708);
	I35710<= not (CRC_OUT_1_7 and I35708);
	I35715<= not (WX10980 and CRC_OUT_1_6);
	I35716<= not (WX10980 and I35715);
	I35717<= not (CRC_OUT_1_6 and I35715);
	I35722<= not (WX10981 and CRC_OUT_1_5);
	I35723<= not (WX10981 and I35722);
	I35724<= not (CRC_OUT_1_5 and I35722);
	I35729<= not (WX10982 and CRC_OUT_1_4);
	I35730<= not (WX10982 and I35729);
	I35731<= not (CRC_OUT_1_4 and I35729);
	I35736<= not (WX10984 and CRC_OUT_1_2);
	I35737<= not (WX10984 and I35736);
	I35738<= not (CRC_OUT_1_2 and I35736);
	I35743<= not (WX10985 and CRC_OUT_1_1);
	I35744<= not (WX10985 and I35743);
	I35745<= not (CRC_OUT_1_1 and I35743);
	I35750<= not (WX10986 and CRC_OUT_1_0);
	I35751<= not (WX10986 and I35750);
	I35752<= not (CRC_OUT_1_0 and I35750);
	WX900<= not (I2011 and I2012);
	WX901<= not (I2042 and I2043);
	WX902<= not (I2073 and I2074);
	WX903<= not (I2104 and I2105);
	WX904<= not (I2135 and I2136);
	WX905<= not (I2166 and I2167);
	WX906<= not (I2197 and I2198);
	WX907<= not (I2228 and I2229);
	WX908<= not (I2259 and I2260);
	WX909<= not (I2290 and I2291);
	WX910<= not (I2321 and I2322);
	WX911<= not (I2352 and I2353);
	WX912<= not (I2383 and I2384);
	WX913<= not (I2414 and I2415);
	WX914<= not (I2445 and I2446);
	WX915<= not (I2476 and I2477);
	WX916<= not (I2507 and I2508);
	WX917<= not (I2538 and I2539);
	WX918<= not (I2569 and I2570);
	WX919<= not (I2600 and I2601);
	WX920<= not (I2631 and I2632);
	WX921<= not (I2662 and I2663);
	WX922<= not (I2693 and I2694);
	WX923<= not (I2724 and I2725);
	WX924<= not (I2755 and I2756);
	WX925<= not (I2786 and I2787);
	WX926<= not (I2817 and I2818);
	WX927<= not (I2848 and I2849);
	WX928<= not (I2879 and I2880);
	WX929<= not (I2910 and I2911);
	WX930<= not (I2941 and I2942);
	WX931<= not (I2972 and I2973);
	WX1006<= not (I3053 and I3054);
	WX1013<= not (I3066 and I3067);
	WX1020<= not (I3079 and I3080);
	WX1027<= not (I3092 and I3093);
	WX1034<= not (I3105 and I3106);
	WX1041<= not (I3118 and I3119);
	WX1048<= not (I3131 and I3132);
	WX1055<= not (I3144 and I3145);
	WX1062<= not (I3157 and I3158);
	WX1069<= not (I3170 and I3171);
	WX1076<= not (I3183 and I3184);
	WX1083<= not (I3196 and I3197);
	WX1090<= not (I3209 and I3210);
	WX1097<= not (I3222 and I3223);
	WX1104<= not (I3235 and I3236);
	WX1111<= not (I3248 and I3249);
	WX1118<= not (I3261 and I3262);
	WX1125<= not (I3274 and I3275);
	WX1132<= not (I3287 and I3288);
	WX1139<= not (I3300 and I3301);
	WX1146<= not (I3313 and I3314);
	WX1153<= not (I3326 and I3327);
	WX1160<= not (I3339 and I3340);
	WX1167<= not (I3352 and I3353);
	WX1174<= not (I3365 and I3366);
	WX1181<= not (I3378 and I3379);
	WX1188<= not (I3391 and I3392);
	WX1195<= not (I3404 and I3405);
	WX1202<= not (I3417 and I3418);
	WX1209<= not (I3430 and I3431);
	WX1216<= not (I3443 and I3444);
	WX1223<= not (I3456 and I3457);
	WX1231<= not (I3478 and I3479);
	WX1232<= not (I3493 and I3494);
	WX1233<= not (I3508 and I3509);
	WX1234<= not (I3515 and I3516);
	WX1235<= not (I3522 and I3523);
	WX1236<= not (I3529 and I3530);
	WX1237<= not (I3536 and I3537);
	WX1238<= not (I3543 and I3544);
	WX1239<= not (I3550 and I3551);
	WX1240<= not (I3557 and I3558);
	WX1241<= not (I3564 and I3565);
	WX1242<= not (I3571 and I3572);
	WX1243<= not (I3578 and I3579);
	WX1244<= not (I3585 and I3586);
	WX1245<= not (I3592 and I3593);
	WX1246<= not (I3599 and I3600);
	WX1247<= not (I3606 and I3607);
	WX1248<= not (I3613 and I3614);
	WX1249<= not (I3620 and I3621);
	WX1250<= not (I3627 and I3628);
	WX1251<= not (I3634 and I3635);
	WX1252<= not (I3641 and I3642);
	WX1253<= not (I3648 and I3649);
	WX1254<= not (I3655 and I3656);
	WX1255<= not (I3662 and I3663);
	WX1256<= not (I3669 and I3670);
	WX1257<= not (I3676 and I3677);
	WX1258<= not (I3683 and I3684);
	WX1259<= not (I3690 and I3691);
	WX1260<= not (I3697 and I3698);
	WX1261<= not (I3704 and I3705);
	WX1262<= not (I3711 and I3712);
	WX2193<= not (I6016 and I6017);
	WX2194<= not (I6047 and I6048);
	WX2195<= not (I6078 and I6079);
	WX2196<= not (I6109 and I6110);
	WX2197<= not (I6140 and I6141);
	WX2198<= not (I6171 and I6172);
	WX2199<= not (I6202 and I6203);
	WX2200<= not (I6233 and I6234);
	WX2201<= not (I6264 and I6265);
	WX2202<= not (I6295 and I6296);
	WX2203<= not (I6326 and I6327);
	WX2204<= not (I6357 and I6358);
	WX2205<= not (I6388 and I6389);
	WX2206<= not (I6419 and I6420);
	WX2207<= not (I6450 and I6451);
	WX2208<= not (I6481 and I6482);
	WX2209<= not (I6512 and I6513);
	WX2210<= not (I6543 and I6544);
	WX2211<= not (I6574 and I6575);
	WX2212<= not (I6605 and I6606);
	WX2213<= not (I6636 and I6637);
	WX2214<= not (I6667 and I6668);
	WX2215<= not (I6698 and I6699);
	WX2216<= not (I6729 and I6730);
	WX2217<= not (I6760 and I6761);
	WX2218<= not (I6791 and I6792);
	WX2219<= not (I6822 and I6823);
	WX2220<= not (I6853 and I6854);
	WX2221<= not (I6884 and I6885);
	WX2222<= not (I6915 and I6916);
	WX2223<= not (I6946 and I6947);
	WX2224<= not (I6977 and I6978);
	WX2299<= not (I7058 and I7059);
	WX2306<= not (I7071 and I7072);
	WX2313<= not (I7084 and I7085);
	WX2320<= not (I7097 and I7098);
	WX2327<= not (I7110 and I7111);
	WX2334<= not (I7123 and I7124);
	WX2341<= not (I7136 and I7137);
	WX2348<= not (I7149 and I7150);
	WX2355<= not (I7162 and I7163);
	WX2362<= not (I7175 and I7176);
	WX2369<= not (I7188 and I7189);
	WX2376<= not (I7201 and I7202);
	WX2383<= not (I7214 and I7215);
	WX2390<= not (I7227 and I7228);
	WX2397<= not (I7240 and I7241);
	WX2404<= not (I7253 and I7254);
	WX2411<= not (I7266 and I7267);
	WX2418<= not (I7279 and I7280);
	WX2425<= not (I7292 and I7293);
	WX2432<= not (I7305 and I7306);
	WX2439<= not (I7318 and I7319);
	WX2446<= not (I7331 and I7332);
	WX2453<= not (I7344 and I7345);
	WX2460<= not (I7357 and I7358);
	WX2467<= not (I7370 and I7371);
	WX2474<= not (I7383 and I7384);
	WX2481<= not (I7396 and I7397);
	WX2488<= not (I7409 and I7410);
	WX2495<= not (I7422 and I7423);
	WX2502<= not (I7435 and I7436);
	WX2509<= not (I7448 and I7449);
	WX2516<= not (I7461 and I7462);
	WX2524<= not (I7483 and I7484);
	WX2525<= not (I7498 and I7499);
	WX2526<= not (I7513 and I7514);
	WX2527<= not (I7520 and I7521);
	WX2528<= not (I7527 and I7528);
	WX2529<= not (I7534 and I7535);
	WX2530<= not (I7541 and I7542);
	WX2531<= not (I7548 and I7549);
	WX2532<= not (I7555 and I7556);
	WX2533<= not (I7562 and I7563);
	WX2534<= not (I7569 and I7570);
	WX2535<= not (I7576 and I7577);
	WX2536<= not (I7583 and I7584);
	WX2537<= not (I7590 and I7591);
	WX2538<= not (I7597 and I7598);
	WX2539<= not (I7604 and I7605);
	WX2540<= not (I7611 and I7612);
	WX2541<= not (I7618 and I7619);
	WX2542<= not (I7625 and I7626);
	WX2543<= not (I7632 and I7633);
	WX2544<= not (I7639 and I7640);
	WX2545<= not (I7646 and I7647);
	WX2546<= not (I7653 and I7654);
	WX2547<= not (I7660 and I7661);
	WX2548<= not (I7667 and I7668);
	WX2549<= not (I7674 and I7675);
	WX2550<= not (I7681 and I7682);
	WX2551<= not (I7688 and I7689);
	WX2552<= not (I7695 and I7696);
	WX2553<= not (I7702 and I7703);
	WX2554<= not (I7709 and I7710);
	WX2555<= not (I7716 and I7717);
	WX3486<= not (I10021 and I10022);
	WX3487<= not (I10052 and I10053);
	WX3488<= not (I10083 and I10084);
	WX3489<= not (I10114 and I10115);
	WX3490<= not (I10145 and I10146);
	WX3491<= not (I10176 and I10177);
	WX3492<= not (I10207 and I10208);
	WX3493<= not (I10238 and I10239);
	WX3494<= not (I10269 and I10270);
	WX3495<= not (I10300 and I10301);
	WX3496<= not (I10331 and I10332);
	WX3497<= not (I10362 and I10363);
	WX3498<= not (I10393 and I10394);
	WX3499<= not (I10424 and I10425);
	WX3500<= not (I10455 and I10456);
	WX3501<= not (I10486 and I10487);
	WX3502<= not (I10517 and I10518);
	WX3503<= not (I10548 and I10549);
	WX3504<= not (I10579 and I10580);
	WX3505<= not (I10610 and I10611);
	WX3506<= not (I10641 and I10642);
	WX3507<= not (I10672 and I10673);
	WX3508<= not (I10703 and I10704);
	WX3509<= not (I10734 and I10735);
	WX3510<= not (I10765 and I10766);
	WX3511<= not (I10796 and I10797);
	WX3512<= not (I10827 and I10828);
	WX3513<= not (I10858 and I10859);
	WX3514<= not (I10889 and I10890);
	WX3515<= not (I10920 and I10921);
	WX3516<= not (I10951 and I10952);
	WX3517<= not (I10982 and I10983);
	WX3592<= not (I11063 and I11064);
	WX3599<= not (I11076 and I11077);
	WX3606<= not (I11089 and I11090);
	WX3613<= not (I11102 and I11103);
	WX3620<= not (I11115 and I11116);
	WX3627<= not (I11128 and I11129);
	WX3634<= not (I11141 and I11142);
	WX3641<= not (I11154 and I11155);
	WX3648<= not (I11167 and I11168);
	WX3655<= not (I11180 and I11181);
	WX3662<= not (I11193 and I11194);
	WX3669<= not (I11206 and I11207);
	WX3676<= not (I11219 and I11220);
	WX3683<= not (I11232 and I11233);
	WX3690<= not (I11245 and I11246);
	WX3697<= not (I11258 and I11259);
	WX3704<= not (I11271 and I11272);
	WX3711<= not (I11284 and I11285);
	WX3718<= not (I11297 and I11298);
	WX3725<= not (I11310 and I11311);
	WX3732<= not (I11323 and I11324);
	WX3739<= not (I11336 and I11337);
	WX3746<= not (I11349 and I11350);
	WX3753<= not (I11362 and I11363);
	WX3760<= not (I11375 and I11376);
	WX3767<= not (I11388 and I11389);
	WX3774<= not (I11401 and I11402);
	WX3781<= not (I11414 and I11415);
	WX3788<= not (I11427 and I11428);
	WX3795<= not (I11440 and I11441);
	WX3802<= not (I11453 and I11454);
	WX3809<= not (I11466 and I11467);
	WX3817<= not (I11488 and I11489);
	WX3818<= not (I11503 and I11504);
	WX3819<= not (I11518 and I11519);
	WX3820<= not (I11525 and I11526);
	WX3821<= not (I11532 and I11533);
	WX3822<= not (I11539 and I11540);
	WX3823<= not (I11546 and I11547);
	WX3824<= not (I11553 and I11554);
	WX3825<= not (I11560 and I11561);
	WX3826<= not (I11567 and I11568);
	WX3827<= not (I11574 and I11575);
	WX3828<= not (I11581 and I11582);
	WX3829<= not (I11588 and I11589);
	WX3830<= not (I11595 and I11596);
	WX3831<= not (I11602 and I11603);
	WX3832<= not (I11609 and I11610);
	WX3833<= not (I11616 and I11617);
	WX3834<= not (I11623 and I11624);
	WX3835<= not (I11630 and I11631);
	WX3836<= not (I11637 and I11638);
	WX3837<= not (I11644 and I11645);
	WX3838<= not (I11651 and I11652);
	WX3839<= not (I11658 and I11659);
	WX3840<= not (I11665 and I11666);
	WX3841<= not (I11672 and I11673);
	WX3842<= not (I11679 and I11680);
	WX3843<= not (I11686 and I11687);
	WX3844<= not (I11693 and I11694);
	WX3845<= not (I11700 and I11701);
	WX3846<= not (I11707 and I11708);
	WX3847<= not (I11714 and I11715);
	WX3848<= not (I11721 and I11722);
	WX4779<= not (I14026 and I14027);
	WX4780<= not (I14057 and I14058);
	WX4781<= not (I14088 and I14089);
	WX4782<= not (I14119 and I14120);
	WX4783<= not (I14150 and I14151);
	WX4784<= not (I14181 and I14182);
	WX4785<= not (I14212 and I14213);
	WX4786<= not (I14243 and I14244);
	WX4787<= not (I14274 and I14275);
	WX4788<= not (I14305 and I14306);
	WX4789<= not (I14336 and I14337);
	WX4790<= not (I14367 and I14368);
	WX4791<= not (I14398 and I14399);
	WX4792<= not (I14429 and I14430);
	WX4793<= not (I14460 and I14461);
	WX4794<= not (I14491 and I14492);
	WX4795<= not (I14522 and I14523);
	WX4796<= not (I14553 and I14554);
	WX4797<= not (I14584 and I14585);
	WX4798<= not (I14615 and I14616);
	WX4799<= not (I14646 and I14647);
	WX4800<= not (I14677 and I14678);
	WX4801<= not (I14708 and I14709);
	WX4802<= not (I14739 and I14740);
	WX4803<= not (I14770 and I14771);
	WX4804<= not (I14801 and I14802);
	WX4805<= not (I14832 and I14833);
	WX4806<= not (I14863 and I14864);
	WX4807<= not (I14894 and I14895);
	WX4808<= not (I14925 and I14926);
	WX4809<= not (I14956 and I14957);
	WX4810<= not (I14987 and I14988);
	WX4885<= not (I15068 and I15069);
	WX4892<= not (I15081 and I15082);
	WX4899<= not (I15094 and I15095);
	WX4906<= not (I15107 and I15108);
	WX4913<= not (I15120 and I15121);
	WX4920<= not (I15133 and I15134);
	WX4927<= not (I15146 and I15147);
	WX4934<= not (I15159 and I15160);
	WX4941<= not (I15172 and I15173);
	WX4948<= not (I15185 and I15186);
	WX4955<= not (I15198 and I15199);
	WX4962<= not (I15211 and I15212);
	WX4969<= not (I15224 and I15225);
	WX4976<= not (I15237 and I15238);
	WX4983<= not (I15250 and I15251);
	WX4990<= not (I15263 and I15264);
	WX4997<= not (I15276 and I15277);
	WX5004<= not (I15289 and I15290);
	WX5011<= not (I15302 and I15303);
	WX5018<= not (I15315 and I15316);
	WX5025<= not (I15328 and I15329);
	WX5032<= not (I15341 and I15342);
	WX5039<= not (I15354 and I15355);
	WX5046<= not (I15367 and I15368);
	WX5053<= not (I15380 and I15381);
	WX5060<= not (I15393 and I15394);
	WX5067<= not (I15406 and I15407);
	WX5074<= not (I15419 and I15420);
	WX5081<= not (I15432 and I15433);
	WX5088<= not (I15445 and I15446);
	WX5095<= not (I15458 and I15459);
	WX5102<= not (I15471 and I15472);
	WX5110<= not (I15493 and I15494);
	WX5111<= not (I15508 and I15509);
	WX5112<= not (I15523 and I15524);
	WX5113<= not (I15530 and I15531);
	WX5114<= not (I15537 and I15538);
	WX5115<= not (I15544 and I15545);
	WX5116<= not (I15551 and I15552);
	WX5117<= not (I15558 and I15559);
	WX5118<= not (I15565 and I15566);
	WX5119<= not (I15572 and I15573);
	WX5120<= not (I15579 and I15580);
	WX5121<= not (I15586 and I15587);
	WX5122<= not (I15593 and I15594);
	WX5123<= not (I15600 and I15601);
	WX5124<= not (I15607 and I15608);
	WX5125<= not (I15614 and I15615);
	WX5126<= not (I15621 and I15622);
	WX5127<= not (I15628 and I15629);
	WX5128<= not (I15635 and I15636);
	WX5129<= not (I15642 and I15643);
	WX5130<= not (I15649 and I15650);
	WX5131<= not (I15656 and I15657);
	WX5132<= not (I15663 and I15664);
	WX5133<= not (I15670 and I15671);
	WX5134<= not (I15677 and I15678);
	WX5135<= not (I15684 and I15685);
	WX5136<= not (I15691 and I15692);
	WX5137<= not (I15698 and I15699);
	WX5138<= not (I15705 and I15706);
	WX5139<= not (I15712 and I15713);
	WX5140<= not (I15719 and I15720);
	WX5141<= not (I15726 and I15727);
	WX6072<= not (I18031 and I18032);
	WX6073<= not (I18062 and I18063);
	WX6074<= not (I18093 and I18094);
	WX6075<= not (I18124 and I18125);
	WX6076<= not (I18155 and I18156);
	WX6077<= not (I18186 and I18187);
	WX6078<= not (I18217 and I18218);
	WX6079<= not (I18248 and I18249);
	WX6080<= not (I18279 and I18280);
	WX6081<= not (I18310 and I18311);
	WX6082<= not (I18341 and I18342);
	WX6083<= not (I18372 and I18373);
	WX6084<= not (I18403 and I18404);
	WX6085<= not (I18434 and I18435);
	WX6086<= not (I18465 and I18466);
	WX6087<= not (I18496 and I18497);
	WX6088<= not (I18527 and I18528);
	WX6089<= not (I18558 and I18559);
	WX6090<= not (I18589 and I18590);
	WX6091<= not (I18620 and I18621);
	WX6092<= not (I18651 and I18652);
	WX6093<= not (I18682 and I18683);
	WX6094<= not (I18713 and I18714);
	WX6095<= not (I18744 and I18745);
	WX6096<= not (I18775 and I18776);
	WX6097<= not (I18806 and I18807);
	WX6098<= not (I18837 and I18838);
	WX6099<= not (I18868 and I18869);
	WX6100<= not (I18899 and I18900);
	WX6101<= not (I18930 and I18931);
	WX6102<= not (I18961 and I18962);
	WX6103<= not (I18992 and I18993);
	WX6178<= not (I19073 and I19074);
	WX6185<= not (I19086 and I19087);
	WX6192<= not (I19099 and I19100);
	WX6199<= not (I19112 and I19113);
	WX6206<= not (I19125 and I19126);
	WX6213<= not (I19138 and I19139);
	WX6220<= not (I19151 and I19152);
	WX6227<= not (I19164 and I19165);
	WX6234<= not (I19177 and I19178);
	WX6241<= not (I19190 and I19191);
	WX6248<= not (I19203 and I19204);
	WX6255<= not (I19216 and I19217);
	WX6262<= not (I19229 and I19230);
	WX6269<= not (I19242 and I19243);
	WX6276<= not (I19255 and I19256);
	WX6283<= not (I19268 and I19269);
	WX6290<= not (I19281 and I19282);
	WX6297<= not (I19294 and I19295);
	WX6304<= not (I19307 and I19308);
	WX6311<= not (I19320 and I19321);
	WX6318<= not (I19333 and I19334);
	WX6325<= not (I19346 and I19347);
	WX6332<= not (I19359 and I19360);
	WX6339<= not (I19372 and I19373);
	WX6346<= not (I19385 and I19386);
	WX6353<= not (I19398 and I19399);
	WX6360<= not (I19411 and I19412);
	WX6367<= not (I19424 and I19425);
	WX6374<= not (I19437 and I19438);
	WX6381<= not (I19450 and I19451);
	WX6388<= not (I19463 and I19464);
	WX6395<= not (I19476 and I19477);
	WX6403<= not (I19498 and I19499);
	WX6404<= not (I19513 and I19514);
	WX6405<= not (I19528 and I19529);
	WX6406<= not (I19535 and I19536);
	WX6407<= not (I19542 and I19543);
	WX6408<= not (I19549 and I19550);
	WX6409<= not (I19556 and I19557);
	WX6410<= not (I19563 and I19564);
	WX6411<= not (I19570 and I19571);
	WX6412<= not (I19577 and I19578);
	WX6413<= not (I19584 and I19585);
	WX6414<= not (I19591 and I19592);
	WX6415<= not (I19598 and I19599);
	WX6416<= not (I19605 and I19606);
	WX6417<= not (I19612 and I19613);
	WX6418<= not (I19619 and I19620);
	WX6419<= not (I19626 and I19627);
	WX6420<= not (I19633 and I19634);
	WX6421<= not (I19640 and I19641);
	WX6422<= not (I19647 and I19648);
	WX6423<= not (I19654 and I19655);
	WX6424<= not (I19661 and I19662);
	WX6425<= not (I19668 and I19669);
	WX6426<= not (I19675 and I19676);
	WX6427<= not (I19682 and I19683);
	WX6428<= not (I19689 and I19690);
	WX6429<= not (I19696 and I19697);
	WX6430<= not (I19703 and I19704);
	WX6431<= not (I19710 and I19711);
	WX6432<= not (I19717 and I19718);
	WX6433<= not (I19724 and I19725);
	WX6434<= not (I19731 and I19732);
	WX7365<= not (I22036 and I22037);
	WX7366<= not (I22067 and I22068);
	WX7367<= not (I22098 and I22099);
	WX7368<= not (I22129 and I22130);
	WX7369<= not (I22160 and I22161);
	WX7370<= not (I22191 and I22192);
	WX7371<= not (I22222 and I22223);
	WX7372<= not (I22253 and I22254);
	WX7373<= not (I22284 and I22285);
	WX7374<= not (I22315 and I22316);
	WX7375<= not (I22346 and I22347);
	WX7376<= not (I22377 and I22378);
	WX7377<= not (I22408 and I22409);
	WX7378<= not (I22439 and I22440);
	WX7379<= not (I22470 and I22471);
	WX7380<= not (I22501 and I22502);
	WX7381<= not (I22532 and I22533);
	WX7382<= not (I22563 and I22564);
	WX7383<= not (I22594 and I22595);
	WX7384<= not (I22625 and I22626);
	WX7385<= not (I22656 and I22657);
	WX7386<= not (I22687 and I22688);
	WX7387<= not (I22718 and I22719);
	WX7388<= not (I22749 and I22750);
	WX7389<= not (I22780 and I22781);
	WX7390<= not (I22811 and I22812);
	WX7391<= not (I22842 and I22843);
	WX7392<= not (I22873 and I22874);
	WX7393<= not (I22904 and I22905);
	WX7394<= not (I22935 and I22936);
	WX7395<= not (I22966 and I22967);
	WX7396<= not (I22997 and I22998);
	WX7471<= not (I23078 and I23079);
	WX7478<= not (I23091 and I23092);
	WX7485<= not (I23104 and I23105);
	WX7492<= not (I23117 and I23118);
	WX7499<= not (I23130 and I23131);
	WX7506<= not (I23143 and I23144);
	WX7513<= not (I23156 and I23157);
	WX7520<= not (I23169 and I23170);
	WX7527<= not (I23182 and I23183);
	WX7534<= not (I23195 and I23196);
	WX7541<= not (I23208 and I23209);
	WX7548<= not (I23221 and I23222);
	WX7555<= not (I23234 and I23235);
	WX7562<= not (I23247 and I23248);
	WX7569<= not (I23260 and I23261);
	WX7576<= not (I23273 and I23274);
	WX7583<= not (I23286 and I23287);
	WX7590<= not (I23299 and I23300);
	WX7597<= not (I23312 and I23313);
	WX7604<= not (I23325 and I23326);
	WX7611<= not (I23338 and I23339);
	WX7618<= not (I23351 and I23352);
	WX7625<= not (I23364 and I23365);
	WX7632<= not (I23377 and I23378);
	WX7639<= not (I23390 and I23391);
	WX7646<= not (I23403 and I23404);
	WX7653<= not (I23416 and I23417);
	WX7660<= not (I23429 and I23430);
	WX7667<= not (I23442 and I23443);
	WX7674<= not (I23455 and I23456);
	WX7681<= not (I23468 and I23469);
	WX7688<= not (I23481 and I23482);
	WX7696<= not (I23503 and I23504);
	WX7697<= not (I23518 and I23519);
	WX7698<= not (I23533 and I23534);
	WX7699<= not (I23540 and I23541);
	WX7700<= not (I23547 and I23548);
	WX7701<= not (I23554 and I23555);
	WX7702<= not (I23561 and I23562);
	WX7703<= not (I23568 and I23569);
	WX7704<= not (I23575 and I23576);
	WX7705<= not (I23582 and I23583);
	WX7706<= not (I23589 and I23590);
	WX7707<= not (I23596 and I23597);
	WX7708<= not (I23603 and I23604);
	WX7709<= not (I23610 and I23611);
	WX7710<= not (I23617 and I23618);
	WX7711<= not (I23624 and I23625);
	WX7712<= not (I23631 and I23632);
	WX7713<= not (I23638 and I23639);
	WX7714<= not (I23645 and I23646);
	WX7715<= not (I23652 and I23653);
	WX7716<= not (I23659 and I23660);
	WX7717<= not (I23666 and I23667);
	WX7718<= not (I23673 and I23674);
	WX7719<= not (I23680 and I23681);
	WX7720<= not (I23687 and I23688);
	WX7721<= not (I23694 and I23695);
	WX7722<= not (I23701 and I23702);
	WX7723<= not (I23708 and I23709);
	WX7724<= not (I23715 and I23716);
	WX7725<= not (I23722 and I23723);
	WX7726<= not (I23729 and I23730);
	WX7727<= not (I23736 and I23737);
	WX8658<= not (I26041 and I26042);
	WX8659<= not (I26072 and I26073);
	WX8660<= not (I26103 and I26104);
	WX8661<= not (I26134 and I26135);
	WX8662<= not (I26165 and I26166);
	WX8663<= not (I26196 and I26197);
	WX8664<= not (I26227 and I26228);
	WX8665<= not (I26258 and I26259);
	WX8666<= not (I26289 and I26290);
	WX8667<= not (I26320 and I26321);
	WX8668<= not (I26351 and I26352);
	WX8669<= not (I26382 and I26383);
	WX8670<= not (I26413 and I26414);
	WX8671<= not (I26444 and I26445);
	WX8672<= not (I26475 and I26476);
	WX8673<= not (I26506 and I26507);
	WX8674<= not (I26537 and I26538);
	WX8675<= not (I26568 and I26569);
	WX8676<= not (I26599 and I26600);
	WX8677<= not (I26630 and I26631);
	WX8678<= not (I26661 and I26662);
	WX8679<= not (I26692 and I26693);
	WX8680<= not (I26723 and I26724);
	WX8681<= not (I26754 and I26755);
	WX8682<= not (I26785 and I26786);
	WX8683<= not (I26816 and I26817);
	WX8684<= not (I26847 and I26848);
	WX8685<= not (I26878 and I26879);
	WX8686<= not (I26909 and I26910);
	WX8687<= not (I26940 and I26941);
	WX8688<= not (I26971 and I26972);
	WX8689<= not (I27002 and I27003);
	WX8764<= not (I27083 and I27084);
	WX8771<= not (I27096 and I27097);
	WX8778<= not (I27109 and I27110);
	WX8785<= not (I27122 and I27123);
	WX8792<= not (I27135 and I27136);
	WX8799<= not (I27148 and I27149);
	WX8806<= not (I27161 and I27162);
	WX8813<= not (I27174 and I27175);
	WX8820<= not (I27187 and I27188);
	WX8827<= not (I27200 and I27201);
	WX8834<= not (I27213 and I27214);
	WX8841<= not (I27226 and I27227);
	WX8848<= not (I27239 and I27240);
	WX8855<= not (I27252 and I27253);
	WX8862<= not (I27265 and I27266);
	WX8869<= not (I27278 and I27279);
	WX8876<= not (I27291 and I27292);
	WX8883<= not (I27304 and I27305);
	WX8890<= not (I27317 and I27318);
	WX8897<= not (I27330 and I27331);
	WX8904<= not (I27343 and I27344);
	WX8911<= not (I27356 and I27357);
	WX8918<= not (I27369 and I27370);
	WX8925<= not (I27382 and I27383);
	WX8932<= not (I27395 and I27396);
	WX8939<= not (I27408 and I27409);
	WX8946<= not (I27421 and I27422);
	WX8953<= not (I27434 and I27435);
	WX8960<= not (I27447 and I27448);
	WX8967<= not (I27460 and I27461);
	WX8974<= not (I27473 and I27474);
	WX8981<= not (I27486 and I27487);
	WX8989<= not (I27508 and I27509);
	WX8990<= not (I27523 and I27524);
	WX8991<= not (I27538 and I27539);
	WX8992<= not (I27545 and I27546);
	WX8993<= not (I27552 and I27553);
	WX8994<= not (I27559 and I27560);
	WX8995<= not (I27566 and I27567);
	WX8996<= not (I27573 and I27574);
	WX8997<= not (I27580 and I27581);
	WX8998<= not (I27587 and I27588);
	WX8999<= not (I27594 and I27595);
	WX9000<= not (I27601 and I27602);
	WX9001<= not (I27608 and I27609);
	WX9002<= not (I27615 and I27616);
	WX9003<= not (I27622 and I27623);
	WX9004<= not (I27629 and I27630);
	WX9005<= not (I27636 and I27637);
	WX9006<= not (I27643 and I27644);
	WX9007<= not (I27650 and I27651);
	WX9008<= not (I27657 and I27658);
	WX9009<= not (I27664 and I27665);
	WX9010<= not (I27671 and I27672);
	WX9011<= not (I27678 and I27679);
	WX9012<= not (I27685 and I27686);
	WX9013<= not (I27692 and I27693);
	WX9014<= not (I27699 and I27700);
	WX9015<= not (I27706 and I27707);
	WX9016<= not (I27713 and I27714);
	WX9017<= not (I27720 and I27721);
	WX9018<= not (I27727 and I27728);
	WX9019<= not (I27734 and I27735);
	WX9020<= not (I27741 and I27742);
	WX9951<= not (I30046 and I30047);
	WX9952<= not (I30077 and I30078);
	WX9953<= not (I30108 and I30109);
	WX9954<= not (I30139 and I30140);
	WX9955<= not (I30170 and I30171);
	WX9956<= not (I30201 and I30202);
	WX9957<= not (I30232 and I30233);
	WX9958<= not (I30263 and I30264);
	WX9959<= not (I30294 and I30295);
	WX9960<= not (I30325 and I30326);
	WX9961<= not (I30356 and I30357);
	WX9962<= not (I30387 and I30388);
	WX9963<= not (I30418 and I30419);
	WX9964<= not (I30449 and I30450);
	WX9965<= not (I30480 and I30481);
	WX9966<= not (I30511 and I30512);
	WX9967<= not (I30542 and I30543);
	WX9968<= not (I30573 and I30574);
	WX9969<= not (I30604 and I30605);
	WX9970<= not (I30635 and I30636);
	WX9971<= not (I30666 and I30667);
	WX9972<= not (I30697 and I30698);
	WX9973<= not (I30728 and I30729);
	WX9974<= not (I30759 and I30760);
	WX9975<= not (I30790 and I30791);
	WX9976<= not (I30821 and I30822);
	WX9977<= not (I30852 and I30853);
	WX9978<= not (I30883 and I30884);
	WX9979<= not (I30914 and I30915);
	WX9980<= not (I30945 and I30946);
	WX9981<= not (I30976 and I30977);
	WX9982<= not (I31007 and I31008);
	WX10057<= not (I31088 and I31089);
	WX10064<= not (I31101 and I31102);
	WX10071<= not (I31114 and I31115);
	WX10078<= not (I31127 and I31128);
	WX10085<= not (I31140 and I31141);
	WX10092<= not (I31153 and I31154);
	WX10099<= not (I31166 and I31167);
	WX10106<= not (I31179 and I31180);
	WX10113<= not (I31192 and I31193);
	WX10120<= not (I31205 and I31206);
	WX10127<= not (I31218 and I31219);
	WX10134<= not (I31231 and I31232);
	WX10141<= not (I31244 and I31245);
	WX10148<= not (I31257 and I31258);
	WX10155<= not (I31270 and I31271);
	WX10162<= not (I31283 and I31284);
	WX10169<= not (I31296 and I31297);
	WX10176<= not (I31309 and I31310);
	WX10183<= not (I31322 and I31323);
	WX10190<= not (I31335 and I31336);
	WX10197<= not (I31348 and I31349);
	WX10204<= not (I31361 and I31362);
	WX10211<= not (I31374 and I31375);
	WX10218<= not (I31387 and I31388);
	WX10225<= not (I31400 and I31401);
	WX10232<= not (I31413 and I31414);
	WX10239<= not (I31426 and I31427);
	WX10246<= not (I31439 and I31440);
	WX10253<= not (I31452 and I31453);
	WX10260<= not (I31465 and I31466);
	WX10267<= not (I31478 and I31479);
	WX10274<= not (I31491 and I31492);
	WX10282<= not (I31513 and I31514);
	WX10283<= not (I31528 and I31529);
	WX10284<= not (I31543 and I31544);
	WX10285<= not (I31550 and I31551);
	WX10286<= not (I31557 and I31558);
	WX10287<= not (I31564 and I31565);
	WX10288<= not (I31571 and I31572);
	WX10289<= not (I31578 and I31579);
	WX10290<= not (I31585 and I31586);
	WX10291<= not (I31592 and I31593);
	WX10292<= not (I31599 and I31600);
	WX10293<= not (I31606 and I31607);
	WX10294<= not (I31613 and I31614);
	WX10295<= not (I31620 and I31621);
	WX10296<= not (I31627 and I31628);
	WX10297<= not (I31634 and I31635);
	WX10298<= not (I31641 and I31642);
	WX10299<= not (I31648 and I31649);
	WX10300<= not (I31655 and I31656);
	WX10301<= not (I31662 and I31663);
	WX10302<= not (I31669 and I31670);
	WX10303<= not (I31676 and I31677);
	WX10304<= not (I31683 and I31684);
	WX10305<= not (I31690 and I31691);
	WX10306<= not (I31697 and I31698);
	WX10307<= not (I31704 and I31705);
	WX10308<= not (I31711 and I31712);
	WX10309<= not (I31718 and I31719);
	WX10310<= not (I31725 and I31726);
	WX10311<= not (I31732 and I31733);
	WX10312<= not (I31739 and I31740);
	WX10313<= not (I31746 and I31747);
	WX11244<= not (I34051 and I34052);
	WX11245<= not (I34082 and I34083);
	WX11246<= not (I34113 and I34114);
	WX11247<= not (I34144 and I34145);
	WX11248<= not (I34175 and I34176);
	WX11249<= not (I34206 and I34207);
	WX11250<= not (I34237 and I34238);
	WX11251<= not (I34268 and I34269);
	WX11252<= not (I34299 and I34300);
	WX11253<= not (I34330 and I34331);
	WX11254<= not (I34361 and I34362);
	WX11255<= not (I34392 and I34393);
	WX11256<= not (I34423 and I34424);
	WX11257<= not (I34454 and I34455);
	WX11258<= not (I34485 and I34486);
	WX11259<= not (I34516 and I34517);
	WX11260<= not (I34547 and I34548);
	WX11261<= not (I34578 and I34579);
	WX11262<= not (I34609 and I34610);
	WX11263<= not (I34640 and I34641);
	WX11264<= not (I34671 and I34672);
	WX11265<= not (I34702 and I34703);
	WX11266<= not (I34733 and I34734);
	WX11267<= not (I34764 and I34765);
	WX11268<= not (I34795 and I34796);
	WX11269<= not (I34826 and I34827);
	WX11270<= not (I34857 and I34858);
	WX11271<= not (I34888 and I34889);
	WX11272<= not (I34919 and I34920);
	WX11273<= not (I34950 and I34951);
	WX11274<= not (I34981 and I34982);
	WX11275<= not (I35012 and I35013);
	WX11350<= not (I35093 and I35094);
	WX11357<= not (I35106 and I35107);
	WX11364<= not (I35119 and I35120);
	WX11371<= not (I35132 and I35133);
	WX11378<= not (I35145 and I35146);
	WX11385<= not (I35158 and I35159);
	WX11392<= not (I35171 and I35172);
	WX11399<= not (I35184 and I35185);
	WX11406<= not (I35197 and I35198);
	WX11413<= not (I35210 and I35211);
	WX11420<= not (I35223 and I35224);
	WX11427<= not (I35236 and I35237);
	WX11434<= not (I35249 and I35250);
	WX11441<= not (I35262 and I35263);
	WX11448<= not (I35275 and I35276);
	WX11455<= not (I35288 and I35289);
	WX11462<= not (I35301 and I35302);
	WX11469<= not (I35314 and I35315);
	WX11476<= not (I35327 and I35328);
	WX11483<= not (I35340 and I35341);
	WX11490<= not (I35353 and I35354);
	WX11497<= not (I35366 and I35367);
	WX11504<= not (I35379 and I35380);
	WX11511<= not (I35392 and I35393);
	WX11518<= not (I35405 and I35406);
	WX11525<= not (I35418 and I35419);
	WX11532<= not (I35431 and I35432);
	WX11539<= not (I35444 and I35445);
	WX11546<= not (I35457 and I35458);
	WX11553<= not (I35470 and I35471);
	WX11560<= not (I35483 and I35484);
	WX11567<= not (I35496 and I35497);
	WX11575<= not (I35518 and I35519);
	WX11576<= not (I35533 and I35534);
	WX11577<= not (I35548 and I35549);
	WX11578<= not (I35555 and I35556);
	WX11579<= not (I35562 and I35563);
	WX11580<= not (I35569 and I35570);
	WX11581<= not (I35576 and I35577);
	WX11582<= not (I35583 and I35584);
	WX11583<= not (I35590 and I35591);
	WX11584<= not (I35597 and I35598);
	WX11585<= not (I35604 and I35605);
	WX11586<= not (I35611 and I35612);
	WX11587<= not (I35618 and I35619);
	WX11588<= not (I35625 and I35626);
	WX11589<= not (I35632 and I35633);
	WX11590<= not (I35639 and I35640);
	WX11591<= not (I35646 and I35647);
	WX11592<= not (I35653 and I35654);
	WX11593<= not (I35660 and I35661);
	WX11594<= not (I35667 and I35668);
	WX11595<= not (I35674 and I35675);
	WX11596<= not (I35681 and I35682);
	WX11597<= not (I35688 and I35689);
	WX11598<= not (I35695 and I35696);
	WX11599<= not (I35702 and I35703);
	WX11600<= not (I35709 and I35710);
	WX11601<= not (I35716 and I35717);
	WX11602<= not (I35723 and I35724);
	WX11603<= not (I35730 and I35731);
	WX11604<= not (I35737 and I35738);
	WX11605<= not (I35744 and I35745);
	WX11606<= not (I35751 and I35752);
	WX38<=WX36 or WX35;
	WX42<=WX40 or WX39;
	WX46<=WX44 or WX43;
	WX52<=WX50 or WX49;
	WX56<=WX54 or WX53;
	WX60<=WX58 or WX57;
	WX66<=WX64 or WX63;
	WX70<=WX68 or WX67;
	WX74<=WX72 or WX71;
	WX80<=WX78 or WX77;
	WX84<=WX82 or WX81;
	WX88<=WX86 or WX85;
	WX94<=WX92 or WX91;
	WX98<=WX96 or WX95;
	WX102<=WX100 or WX99;
	WX108<=WX106 or WX105;
	WX112<=WX110 or WX109;
	WX116<=WX114 or WX113;
	WX122<=WX120 or WX119;
	WX126<=WX124 or WX123;
	WX130<=WX128 or WX127;
	WX136<=WX134 or WX133;
	WX140<=WX138 or WX137;
	WX144<=WX142 or WX141;
	WX150<=WX148 or WX147;
	WX154<=WX152 or WX151;
	WX158<=WX156 or WX155;
	WX164<=WX162 or WX161;
	WX168<=WX166 or WX165;
	WX172<=WX170 or WX169;
	WX178<=WX176 or WX175;
	WX182<=WX180 or WX179;
	WX186<=WX184 or WX183;
	WX192<=WX190 or WX189;
	WX196<=WX194 or WX193;
	WX200<=WX198 or WX197;
	WX206<=WX204 or WX203;
	WX210<=WX208 or WX207;
	WX214<=WX212 or WX211;
	WX220<=WX218 or WX217;
	WX224<=WX222 or WX221;
	WX228<=WX226 or WX225;
	WX234<=WX232 or WX231;
	WX238<=WX236 or WX235;
	WX242<=WX240 or WX239;
	WX248<=WX246 or WX245;
	WX252<=WX250 or WX249;
	WX256<=WX254 or WX253;
	WX262<=WX260 or WX259;
	WX266<=WX264 or WX263;
	WX270<=WX268 or WX267;
	WX276<=WX274 or WX273;
	WX280<=WX278 or WX277;
	WX284<=WX282 or WX281;
	WX290<=WX288 or WX287;
	WX294<=WX292 or WX291;
	WX298<=WX296 or WX295;
	WX304<=WX302 or WX301;
	WX308<=WX306 or WX305;
	WX312<=WX310 or WX309;
	WX318<=WX316 or WX315;
	WX322<=WX320 or WX319;
	WX326<=WX324 or WX323;
	WX332<=WX330 or WX329;
	WX336<=WX334 or WX333;
	WX340<=WX338 or WX337;
	WX346<=WX344 or WX343;
	WX350<=WX348 or WX347;
	WX354<=WX352 or WX351;
	WX360<=WX358 or WX357;
	WX364<=WX362 or WX361;
	WX368<=WX366 or WX365;
	WX374<=WX372 or WX371;
	WX378<=WX376 or WX375;
	WX382<=WX380 or WX379;
	WX388<=WX386 or WX385;
	WX392<=WX390 or WX389;
	WX396<=WX394 or WX393;
	WX402<=WX400 or WX399;
	WX406<=WX404 or WX403;
	WX410<=WX408 or WX407;
	WX416<=WX414 or WX413;
	WX420<=WX418 or WX417;
	WX424<=WX422 or WX421;
	WX430<=WX428 or WX427;
	WX434<=WX432 or WX431;
	WX438<=WX436 or WX435;
	WX444<=WX442 or WX441;
	WX448<=WX446 or WX445;
	WX452<=WX450 or WX449;
	WX458<=WX456 or WX455;
	WX462<=WX460 or WX459;
	WX466<=WX464 or WX463;
	WX472<=WX470 or WX469;
	WX476<=WX474 or WX473;
	WX480<=WX478 or WX477;
	WX1010<=WX1008 or WX1007;
	WX1017<=WX1015 or WX1014;
	WX1024<=WX1022 or WX1021;
	WX1031<=WX1029 or WX1028;
	WX1038<=WX1036 or WX1035;
	WX1045<=WX1043 or WX1042;
	WX1052<=WX1050 or WX1049;
	WX1059<=WX1057 or WX1056;
	WX1066<=WX1064 or WX1063;
	WX1073<=WX1071 or WX1070;
	WX1080<=WX1078 or WX1077;
	WX1087<=WX1085 or WX1084;
	WX1094<=WX1092 or WX1091;
	WX1101<=WX1099 or WX1098;
	WX1108<=WX1106 or WX1105;
	WX1115<=WX1113 or WX1112;
	WX1122<=WX1120 or WX1119;
	WX1129<=WX1127 or WX1126;
	WX1136<=WX1134 or WX1133;
	WX1143<=WX1141 or WX1140;
	WX1150<=WX1148 or WX1147;
	WX1157<=WX1155 or WX1154;
	WX1164<=WX1162 or WX1161;
	WX1171<=WX1169 or WX1168;
	WX1178<=WX1176 or WX1175;
	WX1185<=WX1183 or WX1182;
	WX1192<=WX1190 or WX1189;
	WX1199<=WX1197 or WX1196;
	WX1206<=WX1204 or WX1203;
	WX1213<=WX1211 or WX1210;
	WX1220<=WX1218 or WX1217;
	WX1227<=WX1225 or WX1224;
	WX1331<=WX1329 or WX1328;
	WX1335<=WX1333 or WX1332;
	WX1339<=WX1337 or WX1336;
	WX1345<=WX1343 or WX1342;
	WX1349<=WX1347 or WX1346;
	WX1353<=WX1351 or WX1350;
	WX1359<=WX1357 or WX1356;
	WX1363<=WX1361 or WX1360;
	WX1367<=WX1365 or WX1364;
	WX1373<=WX1371 or WX1370;
	WX1377<=WX1375 or WX1374;
	WX1381<=WX1379 or WX1378;
	WX1387<=WX1385 or WX1384;
	WX1391<=WX1389 or WX1388;
	WX1395<=WX1393 or WX1392;
	WX1401<=WX1399 or WX1398;
	WX1405<=WX1403 or WX1402;
	WX1409<=WX1407 or WX1406;
	WX1415<=WX1413 or WX1412;
	WX1419<=WX1417 or WX1416;
	WX1423<=WX1421 or WX1420;
	WX1429<=WX1427 or WX1426;
	WX1433<=WX1431 or WX1430;
	WX1437<=WX1435 or WX1434;
	WX1443<=WX1441 or WX1440;
	WX1447<=WX1445 or WX1444;
	WX1451<=WX1449 or WX1448;
	WX1457<=WX1455 or WX1454;
	WX1461<=WX1459 or WX1458;
	WX1465<=WX1463 or WX1462;
	WX1471<=WX1469 or WX1468;
	WX1475<=WX1473 or WX1472;
	WX1479<=WX1477 or WX1476;
	WX1485<=WX1483 or WX1482;
	WX1489<=WX1487 or WX1486;
	WX1493<=WX1491 or WX1490;
	WX1499<=WX1497 or WX1496;
	WX1503<=WX1501 or WX1500;
	WX1507<=WX1505 or WX1504;
	WX1513<=WX1511 or WX1510;
	WX1517<=WX1515 or WX1514;
	WX1521<=WX1519 or WX1518;
	WX1527<=WX1525 or WX1524;
	WX1531<=WX1529 or WX1528;
	WX1535<=WX1533 or WX1532;
	WX1541<=WX1539 or WX1538;
	WX1545<=WX1543 or WX1542;
	WX1549<=WX1547 or WX1546;
	WX1555<=WX1553 or WX1552;
	WX1559<=WX1557 or WX1556;
	WX1563<=WX1561 or WX1560;
	WX1569<=WX1567 or WX1566;
	WX1573<=WX1571 or WX1570;
	WX1577<=WX1575 or WX1574;
	WX1583<=WX1581 or WX1580;
	WX1587<=WX1585 or WX1584;
	WX1591<=WX1589 or WX1588;
	WX1597<=WX1595 or WX1594;
	WX1601<=WX1599 or WX1598;
	WX1605<=WX1603 or WX1602;
	WX1611<=WX1609 or WX1608;
	WX1615<=WX1613 or WX1612;
	WX1619<=WX1617 or WX1616;
	WX1625<=WX1623 or WX1622;
	WX1629<=WX1627 or WX1626;
	WX1633<=WX1631 or WX1630;
	WX1639<=WX1637 or WX1636;
	WX1643<=WX1641 or WX1640;
	WX1647<=WX1645 or WX1644;
	WX1653<=WX1651 or WX1650;
	WX1657<=WX1655 or WX1654;
	WX1661<=WX1659 or WX1658;
	WX1667<=WX1665 or WX1664;
	WX1671<=WX1669 or WX1668;
	WX1675<=WX1673 or WX1672;
	WX1681<=WX1679 or WX1678;
	WX1685<=WX1683 or WX1682;
	WX1689<=WX1687 or WX1686;
	WX1695<=WX1693 or WX1692;
	WX1699<=WX1697 or WX1696;
	WX1703<=WX1701 or WX1700;
	WX1709<=WX1707 or WX1706;
	WX1713<=WX1711 or WX1710;
	WX1717<=WX1715 or WX1714;
	WX1723<=WX1721 or WX1720;
	WX1727<=WX1725 or WX1724;
	WX1731<=WX1729 or WX1728;
	WX1737<=WX1735 or WX1734;
	WX1741<=WX1739 or WX1738;
	WX1745<=WX1743 or WX1742;
	WX1751<=WX1749 or WX1748;
	WX1755<=WX1753 or WX1752;
	WX1759<=WX1757 or WX1756;
	WX1765<=WX1763 or WX1762;
	WX1769<=WX1767 or WX1766;
	WX1773<=WX1771 or WX1770;
	WX2303<=WX2301 or WX2300;
	WX2310<=WX2308 or WX2307;
	WX2317<=WX2315 or WX2314;
	WX2324<=WX2322 or WX2321;
	WX2331<=WX2329 or WX2328;
	WX2338<=WX2336 or WX2335;
	WX2345<=WX2343 or WX2342;
	WX2352<=WX2350 or WX2349;
	WX2359<=WX2357 or WX2356;
	WX2366<=WX2364 or WX2363;
	WX2373<=WX2371 or WX2370;
	WX2380<=WX2378 or WX2377;
	WX2387<=WX2385 or WX2384;
	WX2394<=WX2392 or WX2391;
	WX2401<=WX2399 or WX2398;
	WX2408<=WX2406 or WX2405;
	WX2415<=WX2413 or WX2412;
	WX2422<=WX2420 or WX2419;
	WX2429<=WX2427 or WX2426;
	WX2436<=WX2434 or WX2433;
	WX2443<=WX2441 or WX2440;
	WX2450<=WX2448 or WX2447;
	WX2457<=WX2455 or WX2454;
	WX2464<=WX2462 or WX2461;
	WX2471<=WX2469 or WX2468;
	WX2478<=WX2476 or WX2475;
	WX2485<=WX2483 or WX2482;
	WX2492<=WX2490 or WX2489;
	WX2499<=WX2497 or WX2496;
	WX2506<=WX2504 or WX2503;
	WX2513<=WX2511 or WX2510;
	WX2520<=WX2518 or WX2517;
	WX2624<=WX2622 or WX2621;
	WX2628<=WX2626 or WX2625;
	WX2632<=WX2630 or WX2629;
	WX2638<=WX2636 or WX2635;
	WX2642<=WX2640 or WX2639;
	WX2646<=WX2644 or WX2643;
	WX2652<=WX2650 or WX2649;
	WX2656<=WX2654 or WX2653;
	WX2660<=WX2658 or WX2657;
	WX2666<=WX2664 or WX2663;
	WX2670<=WX2668 or WX2667;
	WX2674<=WX2672 or WX2671;
	WX2680<=WX2678 or WX2677;
	WX2684<=WX2682 or WX2681;
	WX2688<=WX2686 or WX2685;
	WX2694<=WX2692 or WX2691;
	WX2698<=WX2696 or WX2695;
	WX2702<=WX2700 or WX2699;
	WX2708<=WX2706 or WX2705;
	WX2712<=WX2710 or WX2709;
	WX2716<=WX2714 or WX2713;
	WX2722<=WX2720 or WX2719;
	WX2726<=WX2724 or WX2723;
	WX2730<=WX2728 or WX2727;
	WX2736<=WX2734 or WX2733;
	WX2740<=WX2738 or WX2737;
	WX2744<=WX2742 or WX2741;
	WX2750<=WX2748 or WX2747;
	WX2754<=WX2752 or WX2751;
	WX2758<=WX2756 or WX2755;
	WX2764<=WX2762 or WX2761;
	WX2768<=WX2766 or WX2765;
	WX2772<=WX2770 or WX2769;
	WX2778<=WX2776 or WX2775;
	WX2782<=WX2780 or WX2779;
	WX2786<=WX2784 or WX2783;
	WX2792<=WX2790 or WX2789;
	WX2796<=WX2794 or WX2793;
	WX2800<=WX2798 or WX2797;
	WX2806<=WX2804 or WX2803;
	WX2810<=WX2808 or WX2807;
	WX2814<=WX2812 or WX2811;
	WX2820<=WX2818 or WX2817;
	WX2824<=WX2822 or WX2821;
	WX2828<=WX2826 or WX2825;
	WX2834<=WX2832 or WX2831;
	WX2838<=WX2836 or WX2835;
	WX2842<=WX2840 or WX2839;
	WX2848<=WX2846 or WX2845;
	WX2852<=WX2850 or WX2849;
	WX2856<=WX2854 or WX2853;
	WX2862<=WX2860 or WX2859;
	WX2866<=WX2864 or WX2863;
	WX2870<=WX2868 or WX2867;
	WX2876<=WX2874 or WX2873;
	WX2880<=WX2878 or WX2877;
	WX2884<=WX2882 or WX2881;
	WX2890<=WX2888 or WX2887;
	WX2894<=WX2892 or WX2891;
	WX2898<=WX2896 or WX2895;
	WX2904<=WX2902 or WX2901;
	WX2908<=WX2906 or WX2905;
	WX2912<=WX2910 or WX2909;
	WX2918<=WX2916 or WX2915;
	WX2922<=WX2920 or WX2919;
	WX2926<=WX2924 or WX2923;
	WX2932<=WX2930 or WX2929;
	WX2936<=WX2934 or WX2933;
	WX2940<=WX2938 or WX2937;
	WX2946<=WX2944 or WX2943;
	WX2950<=WX2948 or WX2947;
	WX2954<=WX2952 or WX2951;
	WX2960<=WX2958 or WX2957;
	WX2964<=WX2962 or WX2961;
	WX2968<=WX2966 or WX2965;
	WX2974<=WX2972 or WX2971;
	WX2978<=WX2976 or WX2975;
	WX2982<=WX2980 or WX2979;
	WX2988<=WX2986 or WX2985;
	WX2992<=WX2990 or WX2989;
	WX2996<=WX2994 or WX2993;
	WX3002<=WX3000 or WX2999;
	WX3006<=WX3004 or WX3003;
	WX3010<=WX3008 or WX3007;
	WX3016<=WX3014 or WX3013;
	WX3020<=WX3018 or WX3017;
	WX3024<=WX3022 or WX3021;
	WX3030<=WX3028 or WX3027;
	WX3034<=WX3032 or WX3031;
	WX3038<=WX3036 or WX3035;
	WX3044<=WX3042 or WX3041;
	WX3048<=WX3046 or WX3045;
	WX3052<=WX3050 or WX3049;
	WX3058<=WX3056 or WX3055;
	WX3062<=WX3060 or WX3059;
	WX3066<=WX3064 or WX3063;
	WX3596<=WX3594 or WX3593;
	WX3603<=WX3601 or WX3600;
	WX3610<=WX3608 or WX3607;
	WX3617<=WX3615 or WX3614;
	WX3624<=WX3622 or WX3621;
	WX3631<=WX3629 or WX3628;
	WX3638<=WX3636 or WX3635;
	WX3645<=WX3643 or WX3642;
	WX3652<=WX3650 or WX3649;
	WX3659<=WX3657 or WX3656;
	WX3666<=WX3664 or WX3663;
	WX3673<=WX3671 or WX3670;
	WX3680<=WX3678 or WX3677;
	WX3687<=WX3685 or WX3684;
	WX3694<=WX3692 or WX3691;
	WX3701<=WX3699 or WX3698;
	WX3708<=WX3706 or WX3705;
	WX3715<=WX3713 or WX3712;
	WX3722<=WX3720 or WX3719;
	WX3729<=WX3727 or WX3726;
	WX3736<=WX3734 or WX3733;
	WX3743<=WX3741 or WX3740;
	WX3750<=WX3748 or WX3747;
	WX3757<=WX3755 or WX3754;
	WX3764<=WX3762 or WX3761;
	WX3771<=WX3769 or WX3768;
	WX3778<=WX3776 or WX3775;
	WX3785<=WX3783 or WX3782;
	WX3792<=WX3790 or WX3789;
	WX3799<=WX3797 or WX3796;
	WX3806<=WX3804 or WX3803;
	WX3813<=WX3811 or WX3810;
	WX3917<=WX3915 or WX3914;
	WX3921<=WX3919 or WX3918;
	WX3925<=WX3923 or WX3922;
	WX3931<=WX3929 or WX3928;
	WX3935<=WX3933 or WX3932;
	WX3939<=WX3937 or WX3936;
	WX3945<=WX3943 or WX3942;
	WX3949<=WX3947 or WX3946;
	WX3953<=WX3951 or WX3950;
	WX3959<=WX3957 or WX3956;
	WX3963<=WX3961 or WX3960;
	WX3967<=WX3965 or WX3964;
	WX3973<=WX3971 or WX3970;
	WX3977<=WX3975 or WX3974;
	WX3981<=WX3979 or WX3978;
	WX3987<=WX3985 or WX3984;
	WX3991<=WX3989 or WX3988;
	WX3995<=WX3993 or WX3992;
	WX4001<=WX3999 or WX3998;
	WX4005<=WX4003 or WX4002;
	WX4009<=WX4007 or WX4006;
	WX4015<=WX4013 or WX4012;
	WX4019<=WX4017 or WX4016;
	WX4023<=WX4021 or WX4020;
	WX4029<=WX4027 or WX4026;
	WX4033<=WX4031 or WX4030;
	WX4037<=WX4035 or WX4034;
	WX4043<=WX4041 or WX4040;
	WX4047<=WX4045 or WX4044;
	WX4051<=WX4049 or WX4048;
	WX4057<=WX4055 or WX4054;
	WX4061<=WX4059 or WX4058;
	WX4065<=WX4063 or WX4062;
	WX4071<=WX4069 or WX4068;
	WX4075<=WX4073 or WX4072;
	WX4079<=WX4077 or WX4076;
	WX4085<=WX4083 or WX4082;
	WX4089<=WX4087 or WX4086;
	WX4093<=WX4091 or WX4090;
	WX4099<=WX4097 or WX4096;
	WX4103<=WX4101 or WX4100;
	WX4107<=WX4105 or WX4104;
	WX4113<=WX4111 or WX4110;
	WX4117<=WX4115 or WX4114;
	WX4121<=WX4119 or WX4118;
	WX4127<=WX4125 or WX4124;
	WX4131<=WX4129 or WX4128;
	WX4135<=WX4133 or WX4132;
	WX4141<=WX4139 or WX4138;
	WX4145<=WX4143 or WX4142;
	WX4149<=WX4147 or WX4146;
	WX4155<=WX4153 or WX4152;
	WX4159<=WX4157 or WX4156;
	WX4163<=WX4161 or WX4160;
	WX4169<=WX4167 or WX4166;
	WX4173<=WX4171 or WX4170;
	WX4177<=WX4175 or WX4174;
	WX4183<=WX4181 or WX4180;
	WX4187<=WX4185 or WX4184;
	WX4191<=WX4189 or WX4188;
	WX4197<=WX4195 or WX4194;
	WX4201<=WX4199 or WX4198;
	WX4205<=WX4203 or WX4202;
	WX4211<=WX4209 or WX4208;
	WX4215<=WX4213 or WX4212;
	WX4219<=WX4217 or WX4216;
	WX4225<=WX4223 or WX4222;
	WX4229<=WX4227 or WX4226;
	WX4233<=WX4231 or WX4230;
	WX4239<=WX4237 or WX4236;
	WX4243<=WX4241 or WX4240;
	WX4247<=WX4245 or WX4244;
	WX4253<=WX4251 or WX4250;
	WX4257<=WX4255 or WX4254;
	WX4261<=WX4259 or WX4258;
	WX4267<=WX4265 or WX4264;
	WX4271<=WX4269 or WX4268;
	WX4275<=WX4273 or WX4272;
	WX4281<=WX4279 or WX4278;
	WX4285<=WX4283 or WX4282;
	WX4289<=WX4287 or WX4286;
	WX4295<=WX4293 or WX4292;
	WX4299<=WX4297 or WX4296;
	WX4303<=WX4301 or WX4300;
	WX4309<=WX4307 or WX4306;
	WX4313<=WX4311 or WX4310;
	WX4317<=WX4315 or WX4314;
	WX4323<=WX4321 or WX4320;
	WX4327<=WX4325 or WX4324;
	WX4331<=WX4329 or WX4328;
	WX4337<=WX4335 or WX4334;
	WX4341<=WX4339 or WX4338;
	WX4345<=WX4343 or WX4342;
	WX4351<=WX4349 or WX4348;
	WX4355<=WX4353 or WX4352;
	WX4359<=WX4357 or WX4356;
	WX4889<=WX4887 or WX4886;
	WX4896<=WX4894 or WX4893;
	WX4903<=WX4901 or WX4900;
	WX4910<=WX4908 or WX4907;
	WX4917<=WX4915 or WX4914;
	WX4924<=WX4922 or WX4921;
	WX4931<=WX4929 or WX4928;
	WX4938<=WX4936 or WX4935;
	WX4945<=WX4943 or WX4942;
	WX4952<=WX4950 or WX4949;
	WX4959<=WX4957 or WX4956;
	WX4966<=WX4964 or WX4963;
	WX4973<=WX4971 or WX4970;
	WX4980<=WX4978 or WX4977;
	WX4987<=WX4985 or WX4984;
	WX4994<=WX4992 or WX4991;
	WX5001<=WX4999 or WX4998;
	WX5008<=WX5006 or WX5005;
	WX5015<=WX5013 or WX5012;
	WX5022<=WX5020 or WX5019;
	WX5029<=WX5027 or WX5026;
	WX5036<=WX5034 or WX5033;
	WX5043<=WX5041 or WX5040;
	WX5050<=WX5048 or WX5047;
	WX5057<=WX5055 or WX5054;
	WX5064<=WX5062 or WX5061;
	WX5071<=WX5069 or WX5068;
	WX5078<=WX5076 or WX5075;
	WX5085<=WX5083 or WX5082;
	WX5092<=WX5090 or WX5089;
	WX5099<=WX5097 or WX5096;
	WX5106<=WX5104 or WX5103;
	WX5210<=WX5208 or WX5207;
	WX5214<=WX5212 or WX5211;
	WX5218<=WX5216 or WX5215;
	WX5224<=WX5222 or WX5221;
	WX5228<=WX5226 or WX5225;
	WX5232<=WX5230 or WX5229;
	WX5238<=WX5236 or WX5235;
	WX5242<=WX5240 or WX5239;
	WX5246<=WX5244 or WX5243;
	WX5252<=WX5250 or WX5249;
	WX5256<=WX5254 or WX5253;
	WX5260<=WX5258 or WX5257;
	WX5266<=WX5264 or WX5263;
	WX5270<=WX5268 or WX5267;
	WX5274<=WX5272 or WX5271;
	WX5280<=WX5278 or WX5277;
	WX5284<=WX5282 or WX5281;
	WX5288<=WX5286 or WX5285;
	WX5294<=WX5292 or WX5291;
	WX5298<=WX5296 or WX5295;
	WX5302<=WX5300 or WX5299;
	WX5308<=WX5306 or WX5305;
	WX5312<=WX5310 or WX5309;
	WX5316<=WX5314 or WX5313;
	WX5322<=WX5320 or WX5319;
	WX5326<=WX5324 or WX5323;
	WX5330<=WX5328 or WX5327;
	WX5336<=WX5334 or WX5333;
	WX5340<=WX5338 or WX5337;
	WX5344<=WX5342 or WX5341;
	WX5350<=WX5348 or WX5347;
	WX5354<=WX5352 or WX5351;
	WX5358<=WX5356 or WX5355;
	WX5364<=WX5362 or WX5361;
	WX5368<=WX5366 or WX5365;
	WX5372<=WX5370 or WX5369;
	WX5378<=WX5376 or WX5375;
	WX5382<=WX5380 or WX5379;
	WX5386<=WX5384 or WX5383;
	WX5392<=WX5390 or WX5389;
	WX5396<=WX5394 or WX5393;
	WX5400<=WX5398 or WX5397;
	WX5406<=WX5404 or WX5403;
	WX5410<=WX5408 or WX5407;
	WX5414<=WX5412 or WX5411;
	WX5420<=WX5418 or WX5417;
	WX5424<=WX5422 or WX5421;
	WX5428<=WX5426 or WX5425;
	WX5434<=WX5432 or WX5431;
	WX5438<=WX5436 or WX5435;
	WX5442<=WX5440 or WX5439;
	WX5448<=WX5446 or WX5445;
	WX5452<=WX5450 or WX5449;
	WX5456<=WX5454 or WX5453;
	WX5462<=WX5460 or WX5459;
	WX5466<=WX5464 or WX5463;
	WX5470<=WX5468 or WX5467;
	WX5476<=WX5474 or WX5473;
	WX5480<=WX5478 or WX5477;
	WX5484<=WX5482 or WX5481;
	WX5490<=WX5488 or WX5487;
	WX5494<=WX5492 or WX5491;
	WX5498<=WX5496 or WX5495;
	WX5504<=WX5502 or WX5501;
	WX5508<=WX5506 or WX5505;
	WX5512<=WX5510 or WX5509;
	WX5518<=WX5516 or WX5515;
	WX5522<=WX5520 or WX5519;
	WX5526<=WX5524 or WX5523;
	WX5532<=WX5530 or WX5529;
	WX5536<=WX5534 or WX5533;
	WX5540<=WX5538 or WX5537;
	WX5546<=WX5544 or WX5543;
	WX5550<=WX5548 or WX5547;
	WX5554<=WX5552 or WX5551;
	WX5560<=WX5558 or WX5557;
	WX5564<=WX5562 or WX5561;
	WX5568<=WX5566 or WX5565;
	WX5574<=WX5572 or WX5571;
	WX5578<=WX5576 or WX5575;
	WX5582<=WX5580 or WX5579;
	WX5588<=WX5586 or WX5585;
	WX5592<=WX5590 or WX5589;
	WX5596<=WX5594 or WX5593;
	WX5602<=WX5600 or WX5599;
	WX5606<=WX5604 or WX5603;
	WX5610<=WX5608 or WX5607;
	WX5616<=WX5614 or WX5613;
	WX5620<=WX5618 or WX5617;
	WX5624<=WX5622 or WX5621;
	WX5630<=WX5628 or WX5627;
	WX5634<=WX5632 or WX5631;
	WX5638<=WX5636 or WX5635;
	WX5644<=WX5642 or WX5641;
	WX5648<=WX5646 or WX5645;
	WX5652<=WX5650 or WX5649;
	WX6182<=WX6180 or WX6179;
	WX6189<=WX6187 or WX6186;
	WX6196<=WX6194 or WX6193;
	WX6203<=WX6201 or WX6200;
	WX6210<=WX6208 or WX6207;
	WX6217<=WX6215 or WX6214;
	WX6224<=WX6222 or WX6221;
	WX6231<=WX6229 or WX6228;
	WX6238<=WX6236 or WX6235;
	WX6245<=WX6243 or WX6242;
	WX6252<=WX6250 or WX6249;
	WX6259<=WX6257 or WX6256;
	WX6266<=WX6264 or WX6263;
	WX6273<=WX6271 or WX6270;
	WX6280<=WX6278 or WX6277;
	WX6287<=WX6285 or WX6284;
	WX6294<=WX6292 or WX6291;
	WX6301<=WX6299 or WX6298;
	WX6308<=WX6306 or WX6305;
	WX6315<=WX6313 or WX6312;
	WX6322<=WX6320 or WX6319;
	WX6329<=WX6327 or WX6326;
	WX6336<=WX6334 or WX6333;
	WX6343<=WX6341 or WX6340;
	WX6350<=WX6348 or WX6347;
	WX6357<=WX6355 or WX6354;
	WX6364<=WX6362 or WX6361;
	WX6371<=WX6369 or WX6368;
	WX6378<=WX6376 or WX6375;
	WX6385<=WX6383 or WX6382;
	WX6392<=WX6390 or WX6389;
	WX6399<=WX6397 or WX6396;
	WX6503<=WX6501 or WX6500;
	WX6507<=WX6505 or WX6504;
	WX6511<=WX6509 or WX6508;
	WX6517<=WX6515 or WX6514;
	WX6521<=WX6519 or WX6518;
	WX6525<=WX6523 or WX6522;
	WX6531<=WX6529 or WX6528;
	WX6535<=WX6533 or WX6532;
	WX6539<=WX6537 or WX6536;
	WX6545<=WX6543 or WX6542;
	WX6549<=WX6547 or WX6546;
	WX6553<=WX6551 or WX6550;
	WX6559<=WX6557 or WX6556;
	WX6563<=WX6561 or WX6560;
	WX6567<=WX6565 or WX6564;
	WX6573<=WX6571 or WX6570;
	WX6577<=WX6575 or WX6574;
	WX6581<=WX6579 or WX6578;
	WX6587<=WX6585 or WX6584;
	WX6591<=WX6589 or WX6588;
	WX6595<=WX6593 or WX6592;
	WX6601<=WX6599 or WX6598;
	WX6605<=WX6603 or WX6602;
	WX6609<=WX6607 or WX6606;
	WX6615<=WX6613 or WX6612;
	WX6619<=WX6617 or WX6616;
	WX6623<=WX6621 or WX6620;
	WX6629<=WX6627 or WX6626;
	WX6633<=WX6631 or WX6630;
	WX6637<=WX6635 or WX6634;
	WX6643<=WX6641 or WX6640;
	WX6647<=WX6645 or WX6644;
	WX6651<=WX6649 or WX6648;
	WX6657<=WX6655 or WX6654;
	WX6661<=WX6659 or WX6658;
	WX6665<=WX6663 or WX6662;
	WX6671<=WX6669 or WX6668;
	WX6675<=WX6673 or WX6672;
	WX6679<=WX6677 or WX6676;
	WX6685<=WX6683 or WX6682;
	WX6689<=WX6687 or WX6686;
	WX6693<=WX6691 or WX6690;
	WX6699<=WX6697 or WX6696;
	WX6703<=WX6701 or WX6700;
	WX6707<=WX6705 or WX6704;
	WX6713<=WX6711 or WX6710;
	WX6717<=WX6715 or WX6714;
	WX6721<=WX6719 or WX6718;
	WX6727<=WX6725 or WX6724;
	WX6731<=WX6729 or WX6728;
	WX6735<=WX6733 or WX6732;
	WX6741<=WX6739 or WX6738;
	WX6745<=WX6743 or WX6742;
	WX6749<=WX6747 or WX6746;
	WX6755<=WX6753 or WX6752;
	WX6759<=WX6757 or WX6756;
	WX6763<=WX6761 or WX6760;
	WX6769<=WX6767 or WX6766;
	WX6773<=WX6771 or WX6770;
	WX6777<=WX6775 or WX6774;
	WX6783<=WX6781 or WX6780;
	WX6787<=WX6785 or WX6784;
	WX6791<=WX6789 or WX6788;
	WX6797<=WX6795 or WX6794;
	WX6801<=WX6799 or WX6798;
	WX6805<=WX6803 or WX6802;
	WX6811<=WX6809 or WX6808;
	WX6815<=WX6813 or WX6812;
	WX6819<=WX6817 or WX6816;
	WX6825<=WX6823 or WX6822;
	WX6829<=WX6827 or WX6826;
	WX6833<=WX6831 or WX6830;
	WX6839<=WX6837 or WX6836;
	WX6843<=WX6841 or WX6840;
	WX6847<=WX6845 or WX6844;
	WX6853<=WX6851 or WX6850;
	WX6857<=WX6855 or WX6854;
	WX6861<=WX6859 or WX6858;
	WX6867<=WX6865 or WX6864;
	WX6871<=WX6869 or WX6868;
	WX6875<=WX6873 or WX6872;
	WX6881<=WX6879 or WX6878;
	WX6885<=WX6883 or WX6882;
	WX6889<=WX6887 or WX6886;
	WX6895<=WX6893 or WX6892;
	WX6899<=WX6897 or WX6896;
	WX6903<=WX6901 or WX6900;
	WX6909<=WX6907 or WX6906;
	WX6913<=WX6911 or WX6910;
	WX6917<=WX6915 or WX6914;
	WX6923<=WX6921 or WX6920;
	WX6927<=WX6925 or WX6924;
	WX6931<=WX6929 or WX6928;
	WX6937<=WX6935 or WX6934;
	WX6941<=WX6939 or WX6938;
	WX6945<=WX6943 or WX6942;
	WX7475<=WX7473 or WX7472;
	WX7482<=WX7480 or WX7479;
	WX7489<=WX7487 or WX7486;
	WX7496<=WX7494 or WX7493;
	WX7503<=WX7501 or WX7500;
	WX7510<=WX7508 or WX7507;
	WX7517<=WX7515 or WX7514;
	WX7524<=WX7522 or WX7521;
	WX7531<=WX7529 or WX7528;
	WX7538<=WX7536 or WX7535;
	WX7545<=WX7543 or WX7542;
	WX7552<=WX7550 or WX7549;
	WX7559<=WX7557 or WX7556;
	WX7566<=WX7564 or WX7563;
	WX7573<=WX7571 or WX7570;
	WX7580<=WX7578 or WX7577;
	WX7587<=WX7585 or WX7584;
	WX7594<=WX7592 or WX7591;
	WX7601<=WX7599 or WX7598;
	WX7608<=WX7606 or WX7605;
	WX7615<=WX7613 or WX7612;
	WX7622<=WX7620 or WX7619;
	WX7629<=WX7627 or WX7626;
	WX7636<=WX7634 or WX7633;
	WX7643<=WX7641 or WX7640;
	WX7650<=WX7648 or WX7647;
	WX7657<=WX7655 or WX7654;
	WX7664<=WX7662 or WX7661;
	WX7671<=WX7669 or WX7668;
	WX7678<=WX7676 or WX7675;
	WX7685<=WX7683 or WX7682;
	WX7692<=WX7690 or WX7689;
	WX7796<=WX7794 or WX7793;
	WX7800<=WX7798 or WX7797;
	WX7804<=WX7802 or WX7801;
	WX7810<=WX7808 or WX7807;
	WX7814<=WX7812 or WX7811;
	WX7818<=WX7816 or WX7815;
	WX7824<=WX7822 or WX7821;
	WX7828<=WX7826 or WX7825;
	WX7832<=WX7830 or WX7829;
	WX7838<=WX7836 or WX7835;
	WX7842<=WX7840 or WX7839;
	WX7846<=WX7844 or WX7843;
	WX7852<=WX7850 or WX7849;
	WX7856<=WX7854 or WX7853;
	WX7860<=WX7858 or WX7857;
	WX7866<=WX7864 or WX7863;
	WX7870<=WX7868 or WX7867;
	WX7874<=WX7872 or WX7871;
	WX7880<=WX7878 or WX7877;
	WX7884<=WX7882 or WX7881;
	WX7888<=WX7886 or WX7885;
	WX7894<=WX7892 or WX7891;
	WX7898<=WX7896 or WX7895;
	WX7902<=WX7900 or WX7899;
	WX7908<=WX7906 or WX7905;
	WX7912<=WX7910 or WX7909;
	WX7916<=WX7914 or WX7913;
	WX7922<=WX7920 or WX7919;
	WX7926<=WX7924 or WX7923;
	WX7930<=WX7928 or WX7927;
	WX7936<=WX7934 or WX7933;
	WX7940<=WX7938 or WX7937;
	WX7944<=WX7942 or WX7941;
	WX7950<=WX7948 or WX7947;
	WX7954<=WX7952 or WX7951;
	WX7958<=WX7956 or WX7955;
	WX7964<=WX7962 or WX7961;
	WX7968<=WX7966 or WX7965;
	WX7972<=WX7970 or WX7969;
	WX7978<=WX7976 or WX7975;
	WX7982<=WX7980 or WX7979;
	WX7986<=WX7984 or WX7983;
	WX7992<=WX7990 or WX7989;
	WX7996<=WX7994 or WX7993;
	WX8000<=WX7998 or WX7997;
	WX8006<=WX8004 or WX8003;
	WX8010<=WX8008 or WX8007;
	WX8014<=WX8012 or WX8011;
	WX8020<=WX8018 or WX8017;
	WX8024<=WX8022 or WX8021;
	WX8028<=WX8026 or WX8025;
	WX8034<=WX8032 or WX8031;
	WX8038<=WX8036 or WX8035;
	WX8042<=WX8040 or WX8039;
	WX8048<=WX8046 or WX8045;
	WX8052<=WX8050 or WX8049;
	WX8056<=WX8054 or WX8053;
	WX8062<=WX8060 or WX8059;
	WX8066<=WX8064 or WX8063;
	WX8070<=WX8068 or WX8067;
	WX8076<=WX8074 or WX8073;
	WX8080<=WX8078 or WX8077;
	WX8084<=WX8082 or WX8081;
	WX8090<=WX8088 or WX8087;
	WX8094<=WX8092 or WX8091;
	WX8098<=WX8096 or WX8095;
	WX8104<=WX8102 or WX8101;
	WX8108<=WX8106 or WX8105;
	WX8112<=WX8110 or WX8109;
	WX8118<=WX8116 or WX8115;
	WX8122<=WX8120 or WX8119;
	WX8126<=WX8124 or WX8123;
	WX8132<=WX8130 or WX8129;
	WX8136<=WX8134 or WX8133;
	WX8140<=WX8138 or WX8137;
	WX8146<=WX8144 or WX8143;
	WX8150<=WX8148 or WX8147;
	WX8154<=WX8152 or WX8151;
	WX8160<=WX8158 or WX8157;
	WX8164<=WX8162 or WX8161;
	WX8168<=WX8166 or WX8165;
	WX8174<=WX8172 or WX8171;
	WX8178<=WX8176 or WX8175;
	WX8182<=WX8180 or WX8179;
	WX8188<=WX8186 or WX8185;
	WX8192<=WX8190 or WX8189;
	WX8196<=WX8194 or WX8193;
	WX8202<=WX8200 or WX8199;
	WX8206<=WX8204 or WX8203;
	WX8210<=WX8208 or WX8207;
	WX8216<=WX8214 or WX8213;
	WX8220<=WX8218 or WX8217;
	WX8224<=WX8222 or WX8221;
	WX8230<=WX8228 or WX8227;
	WX8234<=WX8232 or WX8231;
	WX8238<=WX8236 or WX8235;
	WX8768<=WX8766 or WX8765;
	WX8775<=WX8773 or WX8772;
	WX8782<=WX8780 or WX8779;
	WX8789<=WX8787 or WX8786;
	WX8796<=WX8794 or WX8793;
	WX8803<=WX8801 or WX8800;
	WX8810<=WX8808 or WX8807;
	WX8817<=WX8815 or WX8814;
	WX8824<=WX8822 or WX8821;
	WX8831<=WX8829 or WX8828;
	WX8838<=WX8836 or WX8835;
	WX8845<=WX8843 or WX8842;
	WX8852<=WX8850 or WX8849;
	WX8859<=WX8857 or WX8856;
	WX8866<=WX8864 or WX8863;
	WX8873<=WX8871 or WX8870;
	WX8880<=WX8878 or WX8877;
	WX8887<=WX8885 or WX8884;
	WX8894<=WX8892 or WX8891;
	WX8901<=WX8899 or WX8898;
	WX8908<=WX8906 or WX8905;
	WX8915<=WX8913 or WX8912;
	WX8922<=WX8920 or WX8919;
	WX8929<=WX8927 or WX8926;
	WX8936<=WX8934 or WX8933;
	WX8943<=WX8941 or WX8940;
	WX8950<=WX8948 or WX8947;
	WX8957<=WX8955 or WX8954;
	WX8964<=WX8962 or WX8961;
	WX8971<=WX8969 or WX8968;
	WX8978<=WX8976 or WX8975;
	WX8985<=WX8983 or WX8982;
	WX9089<=WX9087 or WX9086;
	WX9093<=WX9091 or WX9090;
	WX9097<=WX9095 or WX9094;
	WX9103<=WX9101 or WX9100;
	WX9107<=WX9105 or WX9104;
	WX9111<=WX9109 or WX9108;
	WX9117<=WX9115 or WX9114;
	WX9121<=WX9119 or WX9118;
	WX9125<=WX9123 or WX9122;
	WX9131<=WX9129 or WX9128;
	WX9135<=WX9133 or WX9132;
	WX9139<=WX9137 or WX9136;
	WX9145<=WX9143 or WX9142;
	WX9149<=WX9147 or WX9146;
	WX9153<=WX9151 or WX9150;
	WX9159<=WX9157 or WX9156;
	WX9163<=WX9161 or WX9160;
	WX9167<=WX9165 or WX9164;
	WX9173<=WX9171 or WX9170;
	WX9177<=WX9175 or WX9174;
	WX9181<=WX9179 or WX9178;
	WX9187<=WX9185 or WX9184;
	WX9191<=WX9189 or WX9188;
	WX9195<=WX9193 or WX9192;
	WX9201<=WX9199 or WX9198;
	WX9205<=WX9203 or WX9202;
	WX9209<=WX9207 or WX9206;
	WX9215<=WX9213 or WX9212;
	WX9219<=WX9217 or WX9216;
	WX9223<=WX9221 or WX9220;
	WX9229<=WX9227 or WX9226;
	WX9233<=WX9231 or WX9230;
	WX9237<=WX9235 or WX9234;
	WX9243<=WX9241 or WX9240;
	WX9247<=WX9245 or WX9244;
	WX9251<=WX9249 or WX9248;
	WX9257<=WX9255 or WX9254;
	WX9261<=WX9259 or WX9258;
	WX9265<=WX9263 or WX9262;
	WX9271<=WX9269 or WX9268;
	WX9275<=WX9273 or WX9272;
	WX9279<=WX9277 or WX9276;
	WX9285<=WX9283 or WX9282;
	WX9289<=WX9287 or WX9286;
	WX9293<=WX9291 or WX9290;
	WX9299<=WX9297 or WX9296;
	WX9303<=WX9301 or WX9300;
	WX9307<=WX9305 or WX9304;
	WX9313<=WX9311 or WX9310;
	WX9317<=WX9315 or WX9314;
	WX9321<=WX9319 or WX9318;
	WX9327<=WX9325 or WX9324;
	WX9331<=WX9329 or WX9328;
	WX9335<=WX9333 or WX9332;
	WX9341<=WX9339 or WX9338;
	WX9345<=WX9343 or WX9342;
	WX9349<=WX9347 or WX9346;
	WX9355<=WX9353 or WX9352;
	WX9359<=WX9357 or WX9356;
	WX9363<=WX9361 or WX9360;
	WX9369<=WX9367 or WX9366;
	WX9373<=WX9371 or WX9370;
	WX9377<=WX9375 or WX9374;
	WX9383<=WX9381 or WX9380;
	WX9387<=WX9385 or WX9384;
	WX9391<=WX9389 or WX9388;
	WX9397<=WX9395 or WX9394;
	WX9401<=WX9399 or WX9398;
	WX9405<=WX9403 or WX9402;
	WX9411<=WX9409 or WX9408;
	WX9415<=WX9413 or WX9412;
	WX9419<=WX9417 or WX9416;
	WX9425<=WX9423 or WX9422;
	WX9429<=WX9427 or WX9426;
	WX9433<=WX9431 or WX9430;
	WX9439<=WX9437 or WX9436;
	WX9443<=WX9441 or WX9440;
	WX9447<=WX9445 or WX9444;
	WX9453<=WX9451 or WX9450;
	WX9457<=WX9455 or WX9454;
	WX9461<=WX9459 or WX9458;
	WX9467<=WX9465 or WX9464;
	WX9471<=WX9469 or WX9468;
	WX9475<=WX9473 or WX9472;
	WX9481<=WX9479 or WX9478;
	WX9485<=WX9483 or WX9482;
	WX9489<=WX9487 or WX9486;
	WX9495<=WX9493 or WX9492;
	WX9499<=WX9497 or WX9496;
	WX9503<=WX9501 or WX9500;
	WX9509<=WX9507 or WX9506;
	WX9513<=WX9511 or WX9510;
	WX9517<=WX9515 or WX9514;
	WX9523<=WX9521 or WX9520;
	WX9527<=WX9525 or WX9524;
	WX9531<=WX9529 or WX9528;
	WX10061<=WX10059 or WX10058;
	WX10068<=WX10066 or WX10065;
	WX10075<=WX10073 or WX10072;
	WX10082<=WX10080 or WX10079;
	WX10089<=WX10087 or WX10086;
	WX10096<=WX10094 or WX10093;
	WX10103<=WX10101 or WX10100;
	WX10110<=WX10108 or WX10107;
	WX10117<=WX10115 or WX10114;
	WX10124<=WX10122 or WX10121;
	WX10131<=WX10129 or WX10128;
	WX10138<=WX10136 or WX10135;
	WX10145<=WX10143 or WX10142;
	WX10152<=WX10150 or WX10149;
	WX10159<=WX10157 or WX10156;
	WX10166<=WX10164 or WX10163;
	WX10173<=WX10171 or WX10170;
	WX10180<=WX10178 or WX10177;
	WX10187<=WX10185 or WX10184;
	WX10194<=WX10192 or WX10191;
	WX10201<=WX10199 or WX10198;
	WX10208<=WX10206 or WX10205;
	WX10215<=WX10213 or WX10212;
	WX10222<=WX10220 or WX10219;
	WX10229<=WX10227 or WX10226;
	WX10236<=WX10234 or WX10233;
	WX10243<=WX10241 or WX10240;
	WX10250<=WX10248 or WX10247;
	WX10257<=WX10255 or WX10254;
	WX10264<=WX10262 or WX10261;
	WX10271<=WX10269 or WX10268;
	WX10278<=WX10276 or WX10275;
	WX10382<=WX10380 or WX10379;
	WX10386<=WX10384 or WX10383;
	WX10390<=WX10388 or WX10387;
	WX10396<=WX10394 or WX10393;
	WX10400<=WX10398 or WX10397;
	WX10404<=WX10402 or WX10401;
	WX10410<=WX10408 or WX10407;
	WX10414<=WX10412 or WX10411;
	WX10418<=WX10416 or WX10415;
	WX10424<=WX10422 or WX10421;
	WX10428<=WX10426 or WX10425;
	WX10432<=WX10430 or WX10429;
	WX10438<=WX10436 or WX10435;
	WX10442<=WX10440 or WX10439;
	WX10446<=WX10444 or WX10443;
	WX10452<=WX10450 or WX10449;
	WX10456<=WX10454 or WX10453;
	WX10460<=WX10458 or WX10457;
	WX10466<=WX10464 or WX10463;
	WX10470<=WX10468 or WX10467;
	WX10474<=WX10472 or WX10471;
	WX10480<=WX10478 or WX10477;
	WX10484<=WX10482 or WX10481;
	WX10488<=WX10486 or WX10485;
	WX10494<=WX10492 or WX10491;
	WX10498<=WX10496 or WX10495;
	WX10502<=WX10500 or WX10499;
	WX10508<=WX10506 or WX10505;
	WX10512<=WX10510 or WX10509;
	WX10516<=WX10514 or WX10513;
	WX10522<=WX10520 or WX10519;
	WX10526<=WX10524 or WX10523;
	WX10530<=WX10528 or WX10527;
	WX10536<=WX10534 or WX10533;
	WX10540<=WX10538 or WX10537;
	WX10544<=WX10542 or WX10541;
	WX10550<=WX10548 or WX10547;
	WX10554<=WX10552 or WX10551;
	WX10558<=WX10556 or WX10555;
	WX10564<=WX10562 or WX10561;
	WX10568<=WX10566 or WX10565;
	WX10572<=WX10570 or WX10569;
	WX10578<=WX10576 or WX10575;
	WX10582<=WX10580 or WX10579;
	WX10586<=WX10584 or WX10583;
	WX10592<=WX10590 or WX10589;
	WX10596<=WX10594 or WX10593;
	WX10600<=WX10598 or WX10597;
	WX10606<=WX10604 or WX10603;
	WX10610<=WX10608 or WX10607;
	WX10614<=WX10612 or WX10611;
	WX10620<=WX10618 or WX10617;
	WX10624<=WX10622 or WX10621;
	WX10628<=WX10626 or WX10625;
	WX10634<=WX10632 or WX10631;
	WX10638<=WX10636 or WX10635;
	WX10642<=WX10640 or WX10639;
	WX10648<=WX10646 or WX10645;
	WX10652<=WX10650 or WX10649;
	WX10656<=WX10654 or WX10653;
	WX10662<=WX10660 or WX10659;
	WX10666<=WX10664 or WX10663;
	WX10670<=WX10668 or WX10667;
	WX10676<=WX10674 or WX10673;
	WX10680<=WX10678 or WX10677;
	WX10684<=WX10682 or WX10681;
	WX10690<=WX10688 or WX10687;
	WX10694<=WX10692 or WX10691;
	WX10698<=WX10696 or WX10695;
	WX10704<=WX10702 or WX10701;
	WX10708<=WX10706 or WX10705;
	WX10712<=WX10710 or WX10709;
	WX10718<=WX10716 or WX10715;
	WX10722<=WX10720 or WX10719;
	WX10726<=WX10724 or WX10723;
	WX10732<=WX10730 or WX10729;
	WX10736<=WX10734 or WX10733;
	WX10740<=WX10738 or WX10737;
	WX10746<=WX10744 or WX10743;
	WX10750<=WX10748 or WX10747;
	WX10754<=WX10752 or WX10751;
	WX10760<=WX10758 or WX10757;
	WX10764<=WX10762 or WX10761;
	WX10768<=WX10766 or WX10765;
	WX10774<=WX10772 or WX10771;
	WX10778<=WX10776 or WX10775;
	WX10782<=WX10780 or WX10779;
	WX10788<=WX10786 or WX10785;
	WX10792<=WX10790 or WX10789;
	WX10796<=WX10794 or WX10793;
	WX10802<=WX10800 or WX10799;
	WX10806<=WX10804 or WX10803;
	WX10810<=WX10808 or WX10807;
	WX10816<=WX10814 or WX10813;
	WX10820<=WX10818 or WX10817;
	WX10824<=WX10822 or WX10821;
	WX11354<=WX11352 or WX11351;
	WX11361<=WX11359 or WX11358;
	WX11368<=WX11366 or WX11365;
	WX11375<=WX11373 or WX11372;
	WX11382<=WX11380 or WX11379;
	WX11389<=WX11387 or WX11386;
	WX11396<=WX11394 or WX11393;
	WX11403<=WX11401 or WX11400;
	WX11410<=WX11408 or WX11407;
	WX11417<=WX11415 or WX11414;
	WX11424<=WX11422 or WX11421;
	WX11431<=WX11429 or WX11428;
	WX11438<=WX11436 or WX11435;
	WX11445<=WX11443 or WX11442;
	WX11452<=WX11450 or WX11449;
	WX11459<=WX11457 or WX11456;
	WX11466<=WX11464 or WX11463;
	WX11473<=WX11471 or WX11470;
	WX11480<=WX11478 or WX11477;
	WX11487<=WX11485 or WX11484;
	WX11494<=WX11492 or WX11491;
	WX11501<=WX11499 or WX11498;
	WX11508<=WX11506 or WX11505;
	WX11515<=WX11513 or WX11512;
	WX11522<=WX11520 or WX11519;
	WX11529<=WX11527 or WX11526;
	WX11536<=WX11534 or WX11533;
	WX11543<=WX11541 or WX11540;
	WX11550<=WX11548 or WX11547;
	WX11557<=WX11555 or WX11554;
	WX11564<=WX11562 or WX11561;
	WX11571<=WX11569 or WX11568;
end RTL;
