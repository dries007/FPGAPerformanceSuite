-- File created by Bench2VHDL
-- Name: s15850
-- File: bench/s15850.bench
-- Timestamp: 2019-05-21T22:08:29.201835
--
-- Original File
-- =============
--	# s15850.1
--	# 77 inputs
--	# 150 outputs
--	# 534 D-type flipflops
--	# 6324 inverters
--	# 3448 gates (1619 ANDs + 968 NANDs + 710 ORs + 151 NORs)
--	
--	INPUT(g18)
--	INPUT(g27)
--	INPUT(g109)
--	INPUT(g741)
--	INPUT(g742)
--	INPUT(g743)
--	INPUT(g744)
--	INPUT(g872)
--	INPUT(g873)
--	INPUT(g877)
--	INPUT(g881)
--	INPUT(g1712)
--	INPUT(g1960)
--	INPUT(g1961)
--	INPUT(g1696)
--	INPUT(g750)
--	INPUT(g85)
--	INPUT(g42)
--	INPUT(g1700)
--	INPUT(g102)
--	INPUT(g104)
--	INPUT(g101)
--	INPUT(g29)
--	INPUT(g28)
--	INPUT(g103)
--	INPUT(g83)
--	INPUT(g23)
--	INPUT(g87)
--	INPUT(g922)
--	INPUT(g892)
--	INPUT(g84)
--	INPUT(g919)
--	INPUT(g1182)
--	INPUT(g925)
--	INPUT(g48)
--	INPUT(g895)
--	INPUT(g889)
--	INPUT(g1185)
--	INPUT(g41)
--	INPUT(g43)
--	INPUT(g99)
--	INPUT(g1173)
--	INPUT(g1203)
--	INPUT(g1188)
--	INPUT(g1197)
--	INPUT(g46)
--	INPUT(g31)
--	INPUT(g45)
--	INPUT(g92)
--	INPUT(g89)
--	INPUT(g898)
--	INPUT(g91)
--	INPUT(g93)
--	INPUT(g913)
--	INPUT(g82)
--	INPUT(g88)
--	INPUT(g1194)
--	INPUT(g47)
--	INPUT(g96)
--	INPUT(g910)
--	INPUT(g95)
--	INPUT(g904)
--	INPUT(g1176)
--	INPUT(g901)
--	INPUT(g44)
--	INPUT(g916)
--	INPUT(g100)
--	INPUT(g886)
--	INPUT(g30)
--	INPUT(g86)
--	INPUT(g1170)
--	INPUT(g1200)
--	INPUT(g1191)
--	INPUT(g907)
--	INPUT(g90)
--	INPUT(g94)
--	INPUT(g1179)
--	
--	OUTPUT(g2355)
--	OUTPUT(g2601)
--	OUTPUT(g2602)
--	OUTPUT(g2603)
--	OUTPUT(g2604)
--	OUTPUT(g2605)
--	OUTPUT(g2606)
--	OUTPUT(g2607)
--	OUTPUT(g2608)
--	OUTPUT(g2609)
--	OUTPUT(g2610)
--	OUTPUT(g2611)
--	OUTPUT(g2612)
--	OUTPUT(g2648)
--	OUTPUT(g2986)
--	OUTPUT(g3007)
--	OUTPUT(g3069)
--	OUTPUT(g4172)
--	OUTPUT(g4173)
--	OUTPUT(g4174)
--	OUTPUT(g4175)
--	OUTPUT(g4176)
--	OUTPUT(g4177)
--	OUTPUT(g4178)
--	OUTPUT(g4179)
--	OUTPUT(g4180)
--	OUTPUT(g4181)
--	OUTPUT(g4887)
--	OUTPUT(g4888)
--	OUTPUT(g5101)
--	OUTPUT(g5105)
--	OUTPUT(g5658)
--	OUTPUT(g5659)
--	OUTPUT(g5816)
--	OUTPUT(g6920)
--	OUTPUT(g6926)
--	OUTPUT(g6932)
--	OUTPUT(g6942)
--	OUTPUT(g6949)
--	OUTPUT(g6955)
--	OUTPUT(g7744)
--	OUTPUT(g8061)
--	OUTPUT(g8062)
--	OUTPUT(g8271)
--	OUTPUT(g8313)
--	OUTPUT(g8316)
--	OUTPUT(g8318)
--	OUTPUT(g8323)
--	OUTPUT(g8328)
--	OUTPUT(g8331)
--	OUTPUT(g8335)
--	OUTPUT(g8340)
--	OUTPUT(g8347)
--	OUTPUT(g8349)
--	OUTPUT(g8352)
--	OUTPUT(g8561)
--	OUTPUT(g8562)
--	OUTPUT(g8563)
--	OUTPUT(g8564)
--	OUTPUT(g8565)
--	OUTPUT(g8566)
--	OUTPUT(g8976)
--	OUTPUT(g8977)
--	OUTPUT(g8978)
--	OUTPUT(g8979)
--	OUTPUT(g8980)
--	OUTPUT(g8981)
--	OUTPUT(g8982)
--	OUTPUT(g8983)
--	OUTPUT(g8984)
--	OUTPUT(g8985)
--	OUTPUT(g8986)
--	OUTPUT(g9451)
--	OUTPUT(g9961)
--	OUTPUT(g10377)
--	OUTPUT(g10379)
--	OUTPUT(g10455)
--	OUTPUT(g10457)
--	OUTPUT(g10459)
--	OUTPUT(g10461)
--	OUTPUT(g10463)
--	OUTPUT(g10465)
--	OUTPUT(g10628)
--	OUTPUT(g10801)
--	OUTPUT(g11163)
--	OUTPUT(g11206)
--	OUTPUT(g11489)
--	OUTPUT(g6842)
--	OUTPUT(g4171)
--	OUTPUT(g6267)
--	OUTPUT(g6257)
--	OUTPUT(g1957)
--	OUTPUT(g6282)
--	OUTPUT(g6284)
--	OUTPUT(g6281)
--	OUTPUT(g6253)
--	OUTPUT(g6285)
--	OUTPUT(g6283)
--	OUTPUT(g6265)
--	OUTPUT(g3327)
--	OUTPUT(g6269)
--	OUTPUT(g4204)
--	OUTPUT(g4193)
--	OUTPUT(g6266)
--	OUTPUT(g4203)
--	OUTPUT(g4212)
--	OUTPUT(g4196)
--	OUTPUT(g6263)
--	OUTPUT(g4194)
--	OUTPUT(g4192)
--	OUTPUT(g4213)
--	OUTPUT(g6256)
--	OUTPUT(g6258)
--	OUTPUT(g6279)
--	OUTPUT(g4209)
--	OUTPUT(g4208)
--	OUTPUT(g4214)
--	OUTPUT(g4206)
--	OUTPUT(g6261)
--	OUTPUT(g6255)
--	OUTPUT(g6260)
--	OUTPUT(g6274)
--	OUTPUT(g6271)
--	OUTPUT(g4195)
--	OUTPUT(g6273)
--	OUTPUT(g6275)
--	OUTPUT(g4201)
--	OUTPUT(g6264)
--	OUTPUT(g6270)
--	OUTPUT(g4216)
--	OUTPUT(g6262)
--	OUTPUT(g6278)
--	OUTPUT(g4200)
--	OUTPUT(g6277)
--	OUTPUT(g4198)
--	OUTPUT(g4210)
--	OUTPUT(g4197)
--	OUTPUT(g6259)
--	OUTPUT(g4202)
--	OUTPUT(g6280)
--	OUTPUT(g4191)
--	OUTPUT(g6254)
--	OUTPUT(g6268)
--	OUTPUT(g4205)
--	OUTPUT(g4207)
--	OUTPUT(g4215)
--	OUTPUT(g4199)
--	OUTPUT(g6272)
--	OUTPUT(g6276)
--	OUTPUT(g4211)
--	
--	g1289 = DFF(g5660)
--	g1882 = DFF(g9349)
--	g312 = DFF(g5644)
--	g452 = DFF(g11257)
--	g123 = DFF(g8272)
--	g207 = DFF(g7315)
--	g713 = DFF(g9345)
--	g1153 = DFF(g6304)
--	g1209 = DFF(g10873)
--	g1744 = DFF(g5663)
--	g1558 = DFF(g7349)
--	g695 = DFF(g9343)
--	g461 = DFF(g11467)
--	g940 = DFF(g8572)
--	g976 = DFF(g11471)
--	g709 = DFF(g8432)
--	g1092 = DFF(g6810)
--	g1574 = DFF(g7354)
--	g1864 = DFF(g7816)
--	g369 = DFF(g11439)
--	g1580 = DFF(g7356)
--	g1736 = DFF(g6846)
--	g39 = DFF(g10774)
--	g1651 = DFF(g11182)
--	g1424 = DFF(g7330)
--	g1737 = DFF(g1736)
--	g1672 = DFF(g11037)
--	g1077 = DFF(g6805)
--	g1231 = DFF(g8279)
--	g4 = DFF(g8079)
--	g774 = DFF(g7785)
--	g1104 = DFF(g6815)
--	g1304 = DFF(g7290)
--	g243 = DFF(g7325)
--	g1499 = DFF(g8447)
--	g1044 = DFF(g7789)
--	g1444 = DFF(g8987)
--	g757 = DFF(g11179)
--	g786 = DFF(g8436)
--	g1543 = DFF(g7344)
--	g552 = DFF(g11045)
--	g315 = DFF(g5645)
--	g1534 = DFF(g7341)
--	g622 = DFF(g9338)
--	g1927 = DFF(g9354)
--	g1660 = DFF(g11033)
--	g278 = DFF(g7765)
--	g1436 = DFF(g8989)
--	g718 = DFF(g8433)
--	g76 = DFF(g7775)
--	g554 = DFF(g11047)
--	g496 = DFF(g11333)
--	g981 = DFF(g11472)
--	g878 = DFF(g4896)
--	g590 = DFF(g5653)
--	g829 = DFF(g4182)
--	g1095 = DFF(g6811)
--	g704 = DFF(g9344)
--	g1265 = DFF(g7302)
--	g1786 = DFF(g7814)
--	g682 = DFF(g8429)
--	g1296 = DFF(g7292)
--	g587 = DFF(g6295)
--	g52 = DFF(g7777)
--	g646 = DFF(g8065)
--	g327 = DFF(g5649)
--	g1389 = DFF(g6836)
--	g1371 = DFF(g7311)
--	g1956 = DFF(g1955)
--	g1675 = DFF(g11038)
--	g354 = DFF(g11508)
--	g113 = DFF(g7285)
--	g639 = DFF(g8063)
--	g1684 = DFF(g11041)
--	g1639 = DFF(g8448)
--	g1791 = DFF(g8080)
--	g248 = DFF(g7323)
--	g1707 = DFF(g4907)
--	g1759 = DFF(g5668)
--	g351 = DFF(g11507)
--	g1957 = DFF(g1956)
--	g1604 = DFF(g7364)
--	g1098 = DFF(g6812)
--	g932 = DFF(g8570)
--	g126 = DFF(g5642)
--	g1896 = DFF(g8282)
--	g736 = DFF(g8435)
--	g1019 = DFF(g7807)
--	g1362 = DFF(g7305)
--	g745 = DFF(g2639)
--	g1419 = DFF(g7332)
--	g58 = DFF(g7779)
--	g32 = DFF(g11397)
--	g876 = DFF(g878)
--	g1086 = DFF(g6808)
--	g1486 = DFF(g8444)
--	g1730 = DFF(g10881)
--	g1504 = DFF(g7328)
--	g1470 = DFF(g8440)
--	g822 = DFF(g8437)
--	g583 = DFF(g6291)
--	g1678 = DFF(g11039)
--	g174 = DFF(g8423)
--	g1766 = DFF(g7810)
--	g1801 = DFF(g8450)
--	g186 = DFF(g7317)
--	g959 = DFF(g11403)
--	g1169 = DFF(g6314)
--	g1007 = DFF(g7806)
--	g1407 = DFF(g8993)
--	g1059 = DFF(g7794)
--	g1868 = DFF(g7817)
--	g758 = DFF(g6797)
--	g1718 = DFF(g6337)
--	g396 = DFF(g11265)
--	g1015 = DFF(g7808)
--	g38 = DFF(g10872)
--	g632 = DFF(g5655)
--	g1415 = DFF(g7335)
--	g1227 = DFF(g8278)
--	g1721 = DFF(g10878)
--	g882 = DFF(g883)
--	g16 = DFF(g4906)
--	g284 = DFF(g7767)
--	g426 = DFF(g11256)
--	g219 = DFF(g7310)
--	g1216 = DFF(g1360)
--	g806 = DFF(g7289)
--	g1428 = DFF(g8992)
--	g579 = DFF(g6287)
--	g1564 = DFF(g7351)
--	g1741 = DFF(g5662)
--	g225 = DFF(g7309)
--	g281 = DFF(g7766)
--	g1308 = DFF(g11627)
--	g611 = DFF(g9930)
--	g631 = DFF(g5654)
--	g1217 = DFF(g9823)
--	g1589 = DFF(g7359)
--	g1466 = DFF(g8439)
--	g1571 = DFF(g7353)
--	g1861 = DFF(g7815)
--	g1365 = DFF(g7307)
--	g1448 = DFF(g11594)
--	g1711 = DFF(g6335)
--	g1133 = DFF(g6309)
--	g1333 = DFF(g11635)
--	g153 = DFF(g8426)
--	g962 = DFF(g11404)
--	g766 = DFF(g6799)
--	g588 = DFF(g6296)
--	g486 = DFF(g11331)
--	g471 = DFF(g11469)
--	g1397 = DFF(g7322)
--	g580 = DFF(g6288)
--	g1950 = DFF(g8288)
--	g756 = DFF(g755)
--	g635 = DFF(g5656)
--	g1101 = DFF(g6814)
--	g549 = DFF(g11044)
--	g1041 = DFF(g7788)
--	g105 = DFF(g11180)
--	g1669 = DFF(g11036)
--	g1368 = DFF(g7308)
--	g1531 = DFF(g7340)
--	g1458 = DFF(g7327)
--	g572 = DFF(g10877)
--	g1011 = DFF(g7805)
--	g33 = DFF(g10867)
--	g1411 = DFF(g7331)
--	g1074 = DFF(g6813)
--	g444 = DFF(g11259)
--	g1474 = DFF(g8441)
--	g1080 = DFF(g6806)
--	g1713 = DFF(g6336)
--	g333 = DFF(g5651)
--	g269 = DFF(g7762)
--	g401 = DFF(g11266)
--	g1857 = DFF(g11409)
--	g9 = DFF(g7336)
--	g664 = DFF(g8782)
--	g965 = DFF(g11405)
--	g1400 = DFF(g7324)
--	g309 = DFF(g5652)
--	g814 = DFF(g8077)
--	g231 = DFF(g7319)
--	g557 = DFF(g11048)
--	g586 = DFF(g6294)
--	g869 = DFF(g875)
--	g1383 = DFF(g7316)
--	g158 = DFF(g8425)
--	g627 = DFF(g5657)
--	g1023 = DFF(g7799)
--	g259 = DFF(g7755)
--	g1361 = DFF(g1206)
--	g1327 = DFF(g11633)
--	g654 = DFF(g8067)
--	g293 = DFF(g7770)
--	g1346 = DFF(g11656)
--	g1633 = DFF(g8873)
--	g1753 = DFF(g5666)
--	g1508 = DFF(g7329)
--	g1240 = DFF(g7297)
--	g538 = DFF(g11326)
--	g416 = DFF(g11269)
--	g542 = DFF(g11325)
--	g1681 = DFF(g11040)
--	g374 = DFF(g11440)
--	g563 = DFF(g11050)
--	g1914 = DFF(g8284)
--	g530 = DFF(g11328)
--	g575 = DFF(g11052)
--	g1936 = DFF(g9355)
--	g55 = DFF(g7778)
--	g1117 = DFF(g6299)
--	g1317 = DFF(g1356)
--	g357 = DFF(g11509)
--	g386 = DFF(g11263)
--	g1601 = DFF(g7363)
--	g553 = DFF(g11046)
--	g166 = DFF(g7747)
--	g501 = DFF(g11334)
--	g262 = DFF(g7758)
--	g1840 = DFF(g8694)
--	g70 = DFF(g7783)
--	g318 = DFF(g5646)
--	g1356 = DFF(g6818)
--	g794 = DFF(g6800)
--	g36 = DFF(g10870)
--	g302 = DFF(g7773)
--	g342 = DFF(g11513)
--	g1250 = DFF(g7299)
--	g1163 = DFF(g6301)
--	g1810 = DFF(g2044)
--	g1032 = DFF(g7800)
--	g1432 = DFF(g8990)
--	g1053 = DFF(g7792)
--	g1453 = DFF(g7326)
--	g363 = DFF(g11511)
--	g330 = DFF(g5650)
--	g1157 = DFF(g6303)
--	g1357 = DFF(g6330)
--	g35 = DFF(g10869)
--	g928 = DFF(g8569)
--	g261 = DFF(g7757)
--	g516 = DFF(g11337)
--	g254 = DFF(g7759)
--	g778 = DFF(g8076)
--	g861 = DFF(g4190)
--	g1627 = DFF(g8871)
--	g1292 = DFF(g7293)
--	g290 = DFF(g7769)
--	g1850 = DFF(g5671)
--	g770 = DFF(g7288)
--	g1583 = DFF(g7357)
--	g466 = DFF(g11468)
--	g1561 = DFF(g7350)
--	g1527 = DFF(g4899)
--	g1546 = DFF(g7345)
--	g287 = DFF(g7768)
--	g560 = DFF(g11049)
--	g617 = DFF(g8780)
--	g17 = DFF(g4894)
--	g336 = DFF(g11653)
--	g456 = DFF(g11466)
--	g305 = DFF(g5643)
--	g345 = DFF(g11642)
--	g8 = DFF(g2613)
--	g1771 = DFF(g7811)
--	g865 = DFF(g8275)
--	g255 = DFF(g7751)
--	g1945 = DFF(g9356)
--	g1738 = DFF(g5661)
--	g1478 = DFF(g8442)
--	g1035 = DFF(g7787)
--	g1959 = DFF(g4217)
--	g1690 = DFF(g6844)
--	g1482 = DFF(g8443)
--	g1110 = DFF(g6817)
--	g296 = DFF(g7771)
--	g1663 = DFF(g11034)
--	g700 = DFF(g8431)
--	g1762 = DFF(g5669)
--	g360 = DFF(g11510)
--	g192 = DFF(g6837)
--	g1657 = DFF(g10875)
--	g722 = DFF(g9346)
--	g61 = DFF(g7780)
--	g566 = DFF(g11051)
--	g1394 = DFF(g7809)
--	g1089 = DFF(g6809)
--	g883 = DFF(g4897)
--	g1071 = DFF(g6804)
--	g986 = DFF(g11473)
--	g971 = DFF(g11470)
--	g1955 = DFF(g6338)
--	g143 = DFF(g7746)
--	g1814 = DFF(g9825)
--	g1038 = DFF(g7797)
--	g1212 = DFF(g1217)
--	g1918 = DFF(g9353)
--	g782 = DFF(g8273)
--	g1822 = DFF(g9826)
--	g237 = DFF(g7306)
--	g746 = DFF(g2638)
--	g1062 = DFF(g7795)
--	g1462 = DFF(g8438)
--	g178 = DFF(g7748)
--	g366 = DFF(g11512)
--	g837 = DFF(g4184)
--	g599 = DFF(g9819)
--	g1854 = DFF(g11408)
--	g944 = DFF(g11398)
--	g1941 = DFF(g8287)
--	g170 = DFF(g8422)
--	g1520 = DFF(g7334)
--	g686 = DFF(g9342)
--	g953 = DFF(g11401)
--	g1958 = DFF(g6339)
--	g40 = DFF(g10775)
--	g1765 = DFF(g3329)
--	g1733 = DFF(g10882)
--	g1270 = DFF(g7303)
--	g1610 = DFF(g6845)
--	g1796 = DFF(g8280)
--	g1324 = DFF(g11632)
--	g1540 = DFF(g7343)
--	g1377 = DFF(g7312)
--	g1206 = DFF(g4898)
--	g491 = DFF(g11332)
--	g1849 = DFF(g5670)
--	g213 = DFF(g7313)
--	g1781 = DFF(g7813)
--	g1900 = DFF(g9351)
--	g1245 = DFF(g7298)
--	g108 = DFF(g11593)
--	g630 = DFF(g7287)
--	g148 = DFF(g8427)
--	g833 = DFF(g4183)
--	g1923 = DFF(g8285)
--	g936 = DFF(g8571)
--	g1215 = DFF(g6315)
--	g1314 = DFF(g11629)
--	g849 = DFF(g4187)
--	g1336 = DFF(g11654)
--	g272 = DFF(g7763)
--	g1806 = DFF(g8573)
--	g826 = DFF(g8568)
--	g1065 = DFF(g7796)
--	g1887 = DFF(g8281)
--	g37 = DFF(g10871)
--	g968 = DFF(g11406)
--	g1845 = DFF(g5673)
--	g1137 = DFF(g6310)
--	g1891 = DFF(g9350)
--	g1255 = DFF(g7300)
--	g257 = DFF(g7753)
--	g874 = DFF(g9821)
--	g591 = DFF(g9818)
--	g731 = DFF(g9347)
--	g636 = DFF(g8781)
--	g1218 = DFF(g8276)
--	g605 = DFF(g9820)
--	g79 = DFF(g7776)
--	g182 = DFF(g7749)
--	g950 = DFF(g11400)
--	g1129 = DFF(g6308)
--	g857 = DFF(g4189)
--	g448 = DFF(g11258)
--	g1828 = DFF(g9827)
--	g1727 = DFF(g10880)
--	g1592 = DFF(g7360)
--	g1703 = DFF(g6843)
--	g1932 = DFF(g8286)
--	g1624 = DFF(g8870)
--	g26 = DFF(g4885)
--	g1068 = DFF(g6803)
--	g578 = DFF(g6286)
--	g440 = DFF(g11260)
--	g476 = DFF(g11338)
--	g119 = DFF(g7745)
--	g668 = DFF(g9340)
--	g139 = DFF(g8418)
--	g1149 = DFF(g6305)
--	g34 = DFF(g10868)
--	g1848 = DFF(g7366)
--	g263 = DFF(g7760)
--	g818 = DFF(g8274)
--	g1747 = DFF(g5664)
--	g802 = DFF(g6802)
--	g275 = DFF(g7764)
--	g1524 = DFF(g7338)
--	g1577 = DFF(g7355)
--	g810 = DFF(g7786)
--	g391 = DFF(g11264)
--	g658 = DFF(g9339)
--	g1386 = DFF(g7318)
--	g253 = DFF(g7750)
--	g875 = DFF(g9822)
--	g1125 = DFF(g6307)
--	g201 = DFF(g7304)
--	g1280 = DFF(g7295)
--	g1083 = DFF(g6807)
--	g650 = DFF(g8066)
--	g1636 = DFF(g8874)
--	g853 = DFF(g4188)
--	g421 = DFF(g11270)
--	g762 = DFF(g6798)
--	g956 = DFF(g11402)
--	g378 = DFF(g11441)
--	g1756 = DFF(g5667)
--	g589 = DFF(g6297)
--	g841 = DFF(g4185)
--	g1027 = DFF(g7798)
--	g1003 = DFF(g7803)
--	g1403 = DFF(g8991)
--	g1145 = DFF(g6312)
--	g1107 = DFF(g6816)
--	g1223 = DFF(g8277)
--	g406 = DFF(g11267)
--	g1811 = DFF(g11185)
--	g1642 = DFF(g11183)
--	g1047 = DFF(g7790)
--	g1654 = DFF(g10874)
--	g197 = DFF(g6835)
--	g1595 = DFF(g7361)
--	g1537 = DFF(g7342)
--	g727 = DFF(g8434)
--	g999 = DFF(g7804)
--	g798 = DFF(g6801)
--	g481 = DFF(g11324)
--	g754 = DFF(g4895)
--	g1330 = DFF(g11634)
--	g845 = DFF(g4186)
--	g790 = DFF(g8567)
--	g1512 = DFF(g8449)
--	g114 = DFF(g113)
--	g1490 = DFF(g8445)
--	g1166 = DFF(g6300)
--	g1056 = DFF(g7793)
--	g348 = DFF(g11506)
--	g868 = DFF(g874)
--	g1260 = DFF(g7301)
--	g260 = DFF(g7756)
--	g131 = DFF(g8420)
--	g7 = DFF(g2731)
--	g258 = DFF(g7754)
--	g521 = DFF(g11330)
--	g1318 = DFF(g11630)
--	g1872 = DFF(g9348)
--	g677 = DFF(g9341)
--	g582 = DFF(g6290)
--	g1393 = DFF(g7320)
--	g1549 = DFF(g7346)
--	g947 = DFF(g11399)
--	g1834 = DFF(g9895)
--	g1598 = DFF(g7362)
--	g1121 = DFF(g6306)
--	g1321 = DFF(g11631)
--	g506 = DFF(g11335)
--	g546 = DFF(g11043)
--	g1909 = DFF(g9352)
--	g755 = DFF(g6298)
--	g1552 = DFF(g7347)
--	g584 = DFF(g6292)
--	g1687 = DFF(g11042)
--	g1586 = DFF(g7358)
--	g324 = DFF(g5648)
--	g1141 = DFF(g6311)
--	g1570 = DFF(g4900)
--	g1341 = DFF(g11655)
--	g1710 = DFF(g4901)
--	g1645 = DFF(g11184)
--	g115 = DFF(g7321)
--	g135 = DFF(g8419)
--	g525 = DFF(g11329)
--	g581 = DFF(g6289)
--	g1607 = DFF(g7365)
--	g321 = DFF(g5647)
--	g67 = DFF(g7782)
--	g1275 = DFF(g11443)
--	g1311 = DFF(g11628)
--	g1615 = DFF(g8868)
--	g382 = DFF(g11442)
--	g1374 = DFF(g6825)
--	g266 = DFF(g7761)
--	g1284 = DFF(g7294)
--	g1380 = DFF(g7314)
--	g673 = DFF(g8428)
--	g1853 = DFF(g5672)
--	g162 = DFF(g8424)
--	g411 = DFF(g11268)
--	g431 = DFF(g11262)
--	g1905 = DFF(g8283)
--	g1515 = DFF(g7333)
--	g1630 = DFF(g8872)
--	g49 = DFF(g7774)
--	g991 = DFF(g7802)
--	g1300 = DFF(g7291)
--	g339 = DFF(g11505)
--	g256 = DFF(g7752)
--	g1750 = DFF(g5665)
--	g585 = DFF(g6293)
--	g1440 = DFF(g8988)
--	g1666 = DFF(g11035)
--	g1528 = DFF(g7339)
--	g1351 = DFF(g11657)
--	g1648 = DFF(g11181)
--	g127 = DFF(g8421)
--	g1618 = DFF(g11611)
--	g1235 = DFF(g7296)
--	g299 = DFF(g7772)
--	g435 = DFF(g11261)
--	g64 = DFF(g7781)
--	g1555 = DFF(g7348)
--	g995 = DFF(g7801)
--	g1621 = DFF(g8869)
--	g1113 = DFF(g6313)
--	g643 = DFF(g8064)
--	g1494 = DFF(g8446)
--	g1567 = DFF(g7352)
--	g691 = DFF(g8430)
--	g534 = DFF(g11327)
--	g1776 = DFF(g7812)
--	g569 = DFF(g10876)
--	g1160 = DFF(g6302)
--	g1360 = DFF(g9824)
--	g1050 = DFF(g7791)
--	g1 = DFF(g8078)
--	g511 = DFF(g11336)
--	g1724 = DFF(g10879)
--	g12 = DFF(g7337)
--	g1878 = DFF(g8695)
--	g73 = DFF(g7784)
--	
--	I8854 = NOT(g4500)
--	g5652 = NOT(I9117)
--	I12913 = NOT(g7845)
--	g11354 = NOT(I17179)
--	g6837 = NOT(I10891)
--	I10941 = NOT(g6555)
--	I6979 = NOT(g2888)
--	g5843 = NOT(I9458)
--	g2771 = NOT(I5854)
--	g3537 = NOT(g3164)
--	g6062 = NOT(I9699)
--	I9984 = NOT(g5529)
--	I14382 = NOT(g8886)
--	g7706 = NOT(I12335)
--	I13618 = NOT(g8345)
--	I15181 = NOT(g9968)
--	g6620 = NOT(I10573)
--	I12436 = NOT(g7659)
--	g5193 = NOT(g4682)
--	g6462 = NOT(I10394)
--	g8925 = NOT(I14252)
--	I14519 = NOT(g9106)
--	g10289 = NOT(I15691)
--	I14176 = NOT(g8784)
--	I14185 = NOT(g8790)
--	g11181 = NOT(I16944)
--	I14675 = NOT(g9263)
--	g2299 = NOT(g1707)
--	I12607 = NOT(g7633)
--	g3272 = NOT(g2450)
--	g2547 = NOT(g23)
--	g9291 = NOT(g8892)
--	I6001 = NOT(g2548)
--	I7048 = NOT(g2807)
--	g10309 = NOT(I15733)
--	g7029 = NOT(I11180)
--	g4440 = NOT(g4130)
--	I9544 = NOT(g5024)
--	g10288 = NOT(I15688)
--	I12274 = NOT(g7110)
--	I9483 = NOT(g5050)
--	g7787 = NOT(I12526)
--	I6676 = NOT(g2759)
--	I8520 = NOT(g4338)
--	g10571 = NOT(I16236)
--	I17692 = NOT(g11596)
--	I17761 = NOT(g11652)
--	I13469 = NOT(g8147)
--	g9344 = NOT(I14537)
--	g7956 = NOT(g7432)
--	g3417 = NOT(I6624)
--	g4323 = NOT(g4130)
--	I11286 = NOT(g6551)
--	I8031 = NOT(g3540)
--	g7675 = NOT(I12300)
--	g8320 = NOT(I13344)
--	I12565 = NOT(g7388)
--	I16644 = NOT(g10865)
--	I11306 = NOT(g6731)
--	g1981 = NOT(g650)
--	I7333 = NOT(g3729)
--	I13039 = NOT(g8054)
--	g3982 = NOT(g3052)
--	g6249 = NOT(I10006)
--	g9259 = NOT(g8892)
--	I15190 = NOT(g9974)
--	g11426 = NOT(I17331)
--	g9819 = NOT(I14958)
--	g8277 = NOT(I13203)
--	I5050 = NOT(g1216)
--	I5641 = NOT(g546)
--	g5121 = NOT(g4682)
--	g1997 = NOT(g798)
--	g3629 = NOT(g3228)
--	g3328 = NOT(I6501)
--	I12641 = NOT(g7709)
--	g5670 = NOT(I9171)
--	g6842 = NOT(I10898)
--	g8617 = NOT(g8465)
--	I15520 = NOT(g10035)
--	I7396 = NOT(g4102)
--	I7803 = NOT(g3820)
--	g3330 = NOT(I6507)
--	g2991 = NOT(I6233)
--	I9461 = NOT(g4940)
--	g2244 = NOT(I5251)
--	g6192 = NOT(I9923)
--	g6298 = NOT(I10153)
--	g6085 = NOT(I9734)
--	I12153 = NOT(g6874)
--	g4351 = NOT(I7630)
--	I11677 = NOT(g7056)
--	g10687 = NOT(I16356)
--	g4530 = NOT(I7935)
--	g8516 = NOT(I13717)
--	g5232 = NOT(g4640)
--	I13975 = NOT(g8588)
--	g2078 = NOT(g135)
--	I8911 = NOT(g4565)
--	g2340 = NOT(g1918)
--	g7684 = NOT(g7148)
--	I12409 = NOT(g7501)
--	g7745 = NOT(I12400)
--	g8987 = NOT(I14382)
--	g11546 = NOT(g11519)
--	I10729 = NOT(g5935)
--	g5253 = NOT(g4346)
--	g7338 = NOT(I11662)
--	I7509 = NOT(g3566)
--	I9427 = NOT(g4963)
--	g3800 = NOT(g3292)
--	I15088 = NOT(g9832)
--	g2907 = NOT(I6074)
--	g7791 = NOT(I12538)
--	I11143 = NOT(g6446)
--	g6854 = NOT(I10920)
--	g11088 = NOT(I16871)
--	g7309 = NOT(I11575)
--	g8299 = NOT(I13255)
--	I9046 = NOT(g4736)
--	g6941 = NOT(g6503)
--	g2435 = NOT(g201)
--	I14439 = NOT(g8969)
--	g4010 = NOT(g3144)
--	g2082 = NOT(g1371)
--	I6932 = NOT(g2850)
--	I7662 = NOT(g3336)
--	I9446 = NOT(g5052)
--	g5519 = NOT(g4811)
--	g5740 = NOT(I9302)
--	I5289 = NOT(g49)
--	I9514 = NOT(g5094)
--	g7808 = NOT(I12589)
--	g2482 = NOT(I5565)
--	I5658 = NOT(g560)
--	I15497 = NOT(g10119)
--	I6624 = NOT(g2629)
--	g8892 = NOT(I14242)
--	I11169 = NOT(g6481)
--	g3213 = NOT(I6388)
--	I6068 = NOT(g2227)
--	g11497 = NOT(I17510)
--	I13791 = NOT(g8518)
--	I16867 = NOT(g10913)
--	I10349 = NOT(g6215)
--	g10260 = NOT(g10125)
--	g7759 = NOT(I12442)
--	I8473 = NOT(g4577)
--	I14349 = NOT(g8958)
--	g6708 = NOT(I10689)
--	g10668 = NOT(g10563)
--	I5271 = NOT(g70)
--	I9191 = NOT(g5546)
--	I9391 = NOT(g5013)
--	g6219 = NOT(g5426)
--	I15250 = NOT(g9980)
--	I17100 = NOT(g11221)
--	I14906 = NOT(g9508)
--	g9825 = NOT(I14976)
--	g7201 = NOT(I11427)
--	I14083 = NOT(g8747)
--	g10195 = NOT(I15559)
--	I8324 = NOT(g4794)
--	g6031 = NOT(I9642)
--	g2915 = NOT(I6094)
--	I13666 = NOT(g8292)
--	I9695 = NOT(g5212)
--	I11363 = NOT(g6595)
--	I11217 = NOT(g6529)
--	g6431 = NOT(g6145)
--	g6252 = NOT(I10015)
--	g4172 = NOT(I7333)
--	g6812 = NOT(I10846)
--	g8991 = NOT(I14394)
--	g4372 = NOT(I7677)
--	g7049 = NOT(I11228)
--	I6576 = NOT(g2617)
--	g10525 = NOT(g10499)
--	g10488 = NOT(I16101)
--	I10566 = NOT(g5904)
--	I13478 = NOT(g8191)
--	g5586 = NOT(I8996)
--	g8709 = NOT(g8674)
--	g2214 = NOT(g115)
--	I9536 = NOT(g5008)
--	g6176 = NOT(I9905)
--	g4618 = NOT(g3829)
--	I15296 = NOT(g9995)
--	g4143 = NOT(I7291)
--	I7381 = NOT(g4078)
--	I9159 = NOT(g5033)
--	g11339 = NOT(I17142)
--	g8140 = NOT(I13017)
--	I16979 = NOT(g11088)
--	I16496 = NOT(g10707)
--	g8078 = NOT(I12936)
--	I7847 = NOT(g3435)
--	I9359 = NOT(g5576)
--	g8340 = NOT(I13400)
--	g2110 = NOT(I5002)
--	I15338 = NOT(g10013)
--	g6405 = NOT(g6133)
--	g8478 = NOT(I13678)
--	I16111 = NOT(g10385)
--	g4282 = NOT(g4013)
--	g11644 = NOT(I17736)
--	g7604 = NOT(I12162)
--	g9768 = NOT(g9432)
--	g4566 = NOT(g3753)
--	g7098 = NOT(I11333)
--	g10893 = NOT(I16641)
--	I4961 = NOT(g254)
--	g4988 = NOT(I8358)
--	g6286 = NOT(I10117)
--	g8959 = NOT(I14326)
--	I13580 = NOT(g8338)
--	I9016 = NOT(g4722)
--	I6398 = NOT(g2335)
--	g8517 = NOT(I13720)
--	g3348 = NOT(g2733)
--	I15060 = NOT(g9696)
--	I15968 = NOT(g10408)
--	I5332 = NOT(g756)
--	g8482 = NOT(g8329)
--	g2002 = NOT(g818)
--	I10138 = NOT(g5677)
--	g11060 = NOT(g10937)
--	I17407 = NOT(g11417)
--	I12303 = NOT(g7242)
--	g5645 = NOT(I9096)
--	I15855 = NOT(g10336)
--	g2824 = NOT(I5932)
--	g11197 = NOT(g11112)
--	g4555 = NOT(I7964)
--	g5691 = NOT(g5236)
--	I9642 = NOT(g5229)
--	g7539 = NOT(I11953)
--	g7896 = NOT(I12678)
--	g8656 = NOT(I13941)
--	g9887 = NOT(I15068)
--	I8199 = NOT(g4013)
--	g6974 = NOT(g6365)
--	g6270 = NOT(I10069)
--	I14415 = NOT(g8940)
--	g3260 = NOT(I6428)
--	g11411 = NOT(I17274)
--	I10852 = NOT(g6751)
--	g10042 = NOT(I15253)
--	g10255 = NOT(g10139)
--	g6073 = NOT(I9712)
--	g10189 = NOT(I15545)
--	I4903 = NOT(g259)
--	g2877 = NOT(I6025)
--	I11531 = NOT(g7126)
--	g10679 = NOT(g10584)
--	g6796 = NOT(g6252)
--	I8900 = NOT(g4560)
--	I16735 = NOT(g10855)
--	g1968 = NOT(g369)
--	g5879 = NOT(I9498)
--	I10963 = NOT(g6793)
--	g10270 = NOT(g10156)
--	g3463 = NOT(g3256)
--	g7268 = NOT(I11505)
--	g7362 = NOT(I11734)
--	I11740 = NOT(g7030)
--	g10188 = NOT(I15542)
--	I12174 = NOT(g6939)
--	I12796 = NOT(g7543)
--	g5659 = NOT(I9138)
--	g7419 = NOT(g7206)
--	I15503 = NOT(g10044)
--	I17441 = NOT(g11445)
--	g6980 = NOT(I11127)
--	I17206 = NOT(g11323)
--	g4113 = NOT(I7255)
--	g6069 = NOT(I9706)
--	g11503 = NOT(I17528)
--	g7052 = NOT(I11235)
--	g8110 = NOT(g7996)
--	g2556 = NOT(g186)
--	g4313 = NOT(g3586)
--	I16196 = NOT(g10496)
--	I7817 = NOT(g3399)
--	g8310 = NOT(I13314)
--	g10460 = NOT(I15971)
--	g2222 = NOT(g158)
--	I11953 = NOT(g6907)
--	I13373 = NOT(g8226)
--	I6818 = NOT(g2758)
--	g4202 = NOT(I7423)
--	I6867 = NOT(g2949)
--	I9880 = NOT(g5405)
--	g10093 = NOT(I15326)
--	I10484 = NOT(g6155)
--	g9845 = NOT(g9679)
--	g3720 = NOT(I6888)
--	g10267 = NOT(g10130)
--	g10294 = NOT(I15704)
--	I11800 = NOT(g7246)
--	g4908 = NOT(g4396)
--	g5111 = NOT(I8499)
--	g11450 = NOT(I17407)
--	I13800 = NOT(g8500)
--	g5275 = NOT(g4371)
--	I11417 = NOT(g6638)
--	I17758 = NOT(g11647)
--	g3318 = NOT(g2245)
--	g11315 = NOT(I17108)
--	g4094 = NOT(g2744)
--	I17435 = NOT(g11454)
--	g10065 = NOT(I15293)
--	I5092 = NOT(g32)
--	g8002 = NOT(I12832)
--	g5615 = NOT(I9043)
--	g4567 = NOT(g3374)
--	I8259 = NOT(g4590)
--	g11202 = NOT(g11112)
--	g7728 = NOT(I12369)
--	g6287 = NOT(I10120)
--	I14312 = NOT(g8814)
--	I9612 = NOT(g5149)
--	g10875 = NOT(I16595)
--	I9243 = NOT(g5245)
--	g11055 = NOT(g10950)
--	g3393 = NOT(g3144)
--	g9807 = NOT(g9490)
--	g11111 = NOT(g10974)
--	g4776 = NOT(g3586)
--	I9935 = NOT(g5477)
--	g4593 = NOT(I8004)
--	I11964 = NOT(g6910)
--	I7441 = NOT(g3473)
--	I15986 = NOT(g10417)
--	g3971 = NOT(I7104)
--	g7070 = NOT(I11289)
--	g2237 = NOT(g713)
--	g6399 = NOT(I10305)
--	g5284 = NOT(g4376)
--	I11423 = NOT(g6488)
--	g7470 = NOT(g6927)
--	I15741 = NOT(g10260)
--	g7897 = NOT(g7712)
--	g7025 = NOT(g6400)
--	I6370 = NOT(g2356)
--	g7425 = NOT(g7214)
--	I11587 = NOT(g6828)
--	g2844 = NOT(I5966)
--	I12553 = NOT(g7676)
--	I12862 = NOT(g7638)
--	I8215 = NOT(g3981)
--	I10813 = NOT(g6397)
--	g11384 = NOT(I17209)
--	I14799 = NOT(g9661)
--	I6821 = NOT(g3015)
--	g2194 = NOT(g47)
--	g10160 = NOT(I15476)
--	g6797 = NOT(I10801)
--	g11067 = NOT(g10974)
--	g9342 = NOT(I14531)
--	I12326 = NOT(g7246)
--	g8928 = NOT(I14257)
--	g3121 = NOT(g2462)
--	I16280 = NOT(g10537)
--	g4160 = NOT(I7303)
--	g3321 = NOT(I6484)
--	g2089 = NOT(I4917)
--	g4933 = NOT(I8298)
--	I14973 = NOT(g9733)
--	g2731 = NOT(I5789)
--	I16688 = NOT(g10800)
--	I11543 = NOT(g6881)
--	g5420 = NOT(g4300)
--	I15801 = NOT(g10282)
--	I12948 = NOT(g8019)
--	g10455 = NOT(I15956)
--	g8064 = NOT(I12910)
--	g4521 = NOT(g3586)
--	I14805 = NOT(g9360)
--	g6291 = NOT(I10132)
--	g2557 = NOT(g1840)
--	g4050 = NOT(I7163)
--	I13117 = NOT(g7904)
--	I12904 = NOT(g7985)
--	I4873 = NOT(g105)
--	g8785 = NOT(I14090)
--	g4450 = NOT(g3914)
--	g5794 = NOT(I9394)
--	g9097 = NOT(g8892)
--	g2071 = NOT(I4873)
--	g7678 = NOT(I12307)
--	g6144 = NOT(I9857)
--	I11569 = NOT(g6821)
--	g3253 = NOT(I6417)
--	I7743 = NOT(g3762)
--	g6344 = NOT(I10251)
--	g3938 = NOT(g2991)
--	g7331 = NOT(I11641)
--	I15196 = NOT(g9974)
--	g9354 = NOT(I14567)
--	g10201 = NOT(g10175)
--	g7406 = NOT(I11786)
--	g10277 = NOT(I15675)
--	g2242 = NOT(I5245)
--	I9213 = NOT(g4944)
--	g3909 = NOT(g2920)
--	I6106 = NOT(g2116)
--	g7635 = NOT(I12245)
--	I4869 = NOT(g253)
--	I13568 = NOT(g8343)
--	I13747 = NOT(g8299)
--	I15526 = NOT(g10051)
--	g8563 = NOT(I13782)
--	g10075 = NOT(I15302)
--	g4724 = NOT(g3586)
--	g6259 = NOT(I10036)
--	g4179 = NOT(I7354)
--	g7766 = NOT(I12463)
--	I5722 = NOT(g2075)
--	g7682 = NOT(g7148)
--	I13242 = NOT(g8267)
--	I17500 = NOT(g11478)
--	g6694 = NOT(I10663)
--	g4379 = NOT(g3698)
--	g3519 = NOT(g3164)
--	g7801 = NOT(I12568)
--	g7305 = NOT(I11563)
--	I7411 = NOT(g4140)
--	g8295 = NOT(I13239)
--	g2955 = NOT(I6156)
--	I8136 = NOT(g4144)
--	g5628 = NOT(I9062)
--	I6061 = NOT(g2246)
--	I12183 = NOT(g7007)
--	g6852 = NOT(I10914)
--	I11814 = NOT(g7196)
--	g5515 = NOT(g4429)
--	I6461 = NOT(g2261)
--	g5630 = NOT(I9068)
--	I12397 = NOT(g7284)
--	I4917 = NOT(g584)
--	g2254 = NOT(g131)
--	g2814 = NOT(I5916)
--	g11402 = NOT(I17249)
--	g4289 = NOT(g4013)
--	g7748 = NOT(I12409)
--	g4777 = NOT(g3992)
--	I11807 = NOT(g6854)
--	g11457 = NOT(I17424)
--	I9090 = NOT(g5567)
--	g4835 = NOT(I8192)
--	I14400 = NOT(g8891)
--	g2350 = NOT(I5424)
--	g7755 = NOT(I12430)
--	g9267 = NOT(g8892)
--	g9312 = NOT(I14509)
--	I13639 = NOT(g8321)
--	g2038 = NOT(g1776)
--	I8943 = NOT(g4585)
--	I16763 = NOT(g10890)
--	I12933 = NOT(g7899)
--	g7226 = NOT(I11464)
--	g8089 = NOT(g7934)
--	g10352 = NOT(I15820)
--	g2438 = NOT(g243)
--	I11293 = NOT(g6516)
--	I13230 = NOT(g8244)
--	g2773 = NOT(I5858)
--	g4271 = NOT(g3971)
--	I6904 = NOT(g2820)
--	I12508 = NOT(g7731)
--	I11638 = NOT(g6948)
--	I12634 = NOT(g7727)
--	g10155 = NOT(I15461)
--	I17613 = NOT(g11550)
--	g10822 = NOT(I16534)
--	I4786 = NOT(g109)
--	I6046 = NOT(g2218)
--	I9056 = NOT(g4753)
--	g6951 = NOT(I11097)
--	g10266 = NOT(g10129)
--	I8228 = NOT(g4468)
--	I14005 = NOT(g8631)
--	g10170 = NOT(g10118)
--	I8465 = NOT(g4807)
--	I16660 = NOT(g10793)
--	g7045 = NOT(g6435)
--	I10538 = NOT(g5910)
--	I8934 = NOT(g4271)
--	I5424 = NOT(g910)
--	I5795 = NOT(g2462)
--	g7445 = NOT(I11845)
--	g6114 = NOT(I9795)
--	I5737 = NOT(g2100)
--	I6403 = NOT(g2337)
--	I5809 = NOT(g2356)
--	g6314 = NOT(I10201)
--	I7713 = NOT(g3750)
--	g9761 = NOT(g9454)
--	I11841 = NOT(g7226)
--	I11992 = NOT(g7058)
--	I11391 = NOT(g6387)
--	I9851 = NOT(g5405)
--	g2212 = NOT(g686)
--	I13391 = NOT(g8178)
--	g6870 = NOT(I10952)
--	g4674 = NOT(I8050)
--	g8948 = NOT(I14299)
--	g3141 = NOT(g2563)
--	I6391 = NOT(g2478)
--	I5672 = NOT(g569)
--	I15688 = NOT(g10207)
--	g5040 = NOT(I8421)
--	I5077 = NOT(g35)
--	g1983 = NOT(g750)
--	g6825 = NOT(I10873)
--	g3710 = NOT(g3215)
--	g7369 = NOT(g7273)
--	g7602 = NOT(I12156)
--	g10167 = NOT(I15497)
--	g10194 = NOT(g10062)
--	g10589 = NOT(I16252)
--	I16550 = NOT(g10726)
--	g4541 = NOT(I7946)
--	g7007 = NOT(I11146)
--	I17371 = NOT(g11410)
--	I17234 = NOT(g11353)
--	g7920 = NOT(g7516)
--	I11578 = NOT(g6824)
--	I12574 = NOT(g7522)
--	g10524 = NOT(g10458)
--	g2229 = NOT(g162)
--	I15157 = NOT(g9931)
--	I16307 = NOT(g10589)
--	g4332 = NOT(g4130)
--	I12205 = NOT(g6993)
--	g7767 = NOT(I12466)
--	I6159 = NOT(g2123)
--	g11157 = NOT(g10950)
--	g4680 = NOT(g3829)
--	g6136 = NOT(I9845)
--	g8150 = NOT(I13039)
--	g4209 = NOT(I7444)
--	g4353 = NOT(I7636)
--	g5666 = NOT(I9159)
--	g6336 = NOT(I10231)
--	g8350 = NOT(I13430)
--	I13586 = NOT(g8356)
--	g10119 = NOT(I15365)
--	I8337 = NOT(g4352)
--	g8438 = NOT(I13612)
--	g6594 = NOT(I10560)
--	g11066 = NOT(g10974)
--	g4802 = NOT(g3337)
--	I13442 = NOT(g8182)
--	g8009 = NOT(I12849)
--	I5304 = NOT(g79)
--	g10118 = NOT(I15362)
--	I6016 = NOT(g2201)
--	I6757 = NOT(g2732)
--	g7793 = NOT(I12544)
--	I9279 = NOT(g5314)
--	g5648 = NOT(I9105)
--	g6806 = NOT(I10828)
--	g5875 = NOT(g5361)
--	g6943 = NOT(I11079)
--	I16269 = NOT(g10558)
--	I9720 = NOT(g5248)
--	I12592 = NOT(g7445)
--	g10616 = NOT(I16289)
--	g4558 = NOT(g3880)
--	g5655 = NOT(I9126)
--	I13615 = NOT(g8333)
--	g7415 = NOT(I11797)
--	g7227 = NOT(I11467)
--	I9872 = NOT(g5557)
--	g10313 = NOT(I15741)
--	I5926 = NOT(g2172)
--	I13720 = NOT(g8358)
--	I9652 = NOT(g5426)
--	I5754 = NOT(g2304)
--	I10991 = NOT(g6759)
--	I15763 = NOT(g10244)
--	I11275 = NOT(g6502)
--	g10276 = NOT(I15672)
--	g11511 = NOT(I17552)
--	g4901 = NOT(I8268)
--	I7760 = NOT(g3768)
--	I16670 = NOT(g10797)
--	I11746 = NOT(g6857)
--	I13430 = NOT(g8241)
--	g10305 = NOT(I15725)
--	g10254 = NOT(g10196)
--	g4511 = NOT(g3586)
--	g10900 = NOT(I16656)
--	g9576 = NOT(I14713)
--	g2837 = NOT(g2130)
--	g10466 = NOT(I15989)
--	g5884 = NOT(I9505)
--	I5044 = NOT(g1182)
--	g6433 = NOT(I10349)
--	g5839 = NOT(I9452)
--	g8229 = NOT(g7826)
--	I6654 = NOT(g2952)
--	g8993 = NOT(I14400)
--	g2620 = NOT(g1998)
--	I12846 = NOT(g7685)
--	g2462 = NOT(I5555)
--	g9349 = NOT(I14552)
--	I8815 = NOT(g4471)
--	g10101 = NOT(I15335)
--	g10177 = NOT(I15523)
--	I16667 = NOT(g10780)
--	I13806 = NOT(g8478)
--	I7220 = NOT(g3213)
--	I5862 = NOT(g2537)
--	I9598 = NOT(g5120)
--	I7779 = NOT(g3774)
--	I17724 = NOT(g11625)
--	g6845 = NOT(I10907)
--	g7502 = NOT(I11882)
--	I8154 = NOT(g3636)
--	I10584 = NOT(g5864)
--	I17359 = NOT(g11372)
--	g3545 = NOT(I6733)
--	I15314 = NOT(g10007)
--	g11550 = NOT(I17591)
--	I15287 = NOT(g9980)
--	g6195 = NOT(g5426)
--	I7423 = NOT(g3331)
--	g6137 = NOT(I9848)
--	g5667 = NOT(I9162)
--	g6395 = NOT(I10293)
--	g3380 = NOT(I6576)
--	g5143 = NOT(g4682)
--	g6337 = NOT(I10234)
--	I16487 = NOT(g10771)
--	g6913 = NOT(I11021)
--	g10064 = NOT(I15290)
--	g11287 = NOT(g11207)
--	I15085 = NOT(g9720)
--	g2249 = NOT(g127)
--	I9625 = NOT(g5405)
--	g4580 = NOT(g3880)
--	I10759 = NOT(g5803)
--	g11307 = NOT(I17092)
--	g11076 = NOT(I16843)
--	I9232 = NOT(g4944)
--	g7188 = NOT(I11408)
--	g7689 = NOT(I12322)
--	I17121 = NOT(g11231)
--	g11596 = NOT(g11580)
--	g7388 = NOT(I11773)
--	I10114 = NOT(g5768)
--	I9253 = NOT(g5052)
--	I9938 = NOT(g5478)
--	g10874 = NOT(I16592)
--	g11054 = NOT(g10950)
--	g6807 = NOT(I10831)
--	I9813 = NOT(g5241)
--	I6417 = NOT(g2344)
--	g5693 = NOT(I9224)
--	g11243 = NOT(g11112)
--	I17344 = NOT(g11369)
--	g3507 = NOT(g3307)
--	g4262 = NOT(g4013)
--	g2298 = NOT(I5336)
--	g2085 = NOT(I4903)
--	I7665 = NOT(g3732)
--	g10630 = NOT(I16311)
--	g11431 = NOT(I17344)
--	g6859 = NOT(I10937)
--	g7028 = NOT(g6407)
--	I6982 = NOT(g2889)
--	g6266 = NOT(I10057)
--	I15269 = NOT(g9993)
--	g10166 = NOT(I15494)
--	g7030 = NOT(I11183)
--	I12583 = NOT(g7546)
--	I9519 = NOT(g4998)
--	g8062 = NOT(I12904)
--	g7430 = NOT(g7221)
--	I15341 = NOT(g10019)
--	I5414 = NOT(g904)
--	I16286 = NOT(g10540)
--	I7999 = NOT(g4114)
--	g2854 = NOT(I5986)
--	I17173 = NOT(g11293)
--	I5946 = NOT(g2176)
--	I10849 = NOT(g6734)
--	g11341 = NOT(I17146)
--	I7633 = NOT(g3474)
--	g4889 = NOT(I8240)
--	g2941 = NOT(I6118)
--	g6248 = NOT(I10003)
--	g11655 = NOT(I17767)
--	g9258 = NOT(g8892)
--	g3905 = NOT(g2920)
--	g10892 = NOT(I16638)
--	g9818 = NOT(I14955)
--	g9352 = NOT(I14561)
--	I7303 = NOT(g3262)
--	I8293 = NOT(g4779)
--	I10398 = NOT(g5820)
--	I13475 = NOT(g8173)
--	g11180 = NOT(I16941)
--	g7826 = NOT(I12627)
--	g3628 = NOT(g3111)
--	g6255 = NOT(I10024)
--	g4175 = NOT(I7342)
--	g6081 = NOT(g4977)
--	g6815 = NOT(I10855)
--	I10141 = NOT(g5683)
--	g4375 = NOT(g3638)
--	I10804 = NOT(g6388)
--	I5513 = NOT(g255)
--	g3630 = NOT(I6789)
--	g8788 = NOT(I14097)
--	I11222 = NOT(g6533)
--	I12282 = NOT(g7113)
--	I15335 = NOT(g10007)
--	I16601 = NOT(g10806)
--	g5113 = NOT(I8503)
--	g6692 = NOT(I10659)
--	I16187 = NOT(g10492)
--	g6097 = NOT(I9754)
--	I7732 = NOT(g3758)
--	g7910 = NOT(g7460)
--	I12357 = NOT(g7147)
--	g2219 = NOT(g94)
--	g9893 = NOT(I15082)
--	g2640 = NOT(g1984)
--	g6154 = NOT(I9875)
--	g4285 = NOT(g3688)
--	g6354 = NOT(g5867)
--	g2031 = NOT(g1690)
--	g10907 = NOT(I16673)
--	g5202 = NOT(g4640)
--	g6960 = NOT(I11112)
--	I15694 = NOT(g10234)
--	I5378 = NOT(g1857)
--	g2431 = NOT(I5510)
--	I15965 = NOT(g10405)
--	g2252 = NOT(I5271)
--	g2812 = NOT(g2158)
--	I7240 = NOT(g2824)
--	g7609 = NOT(I12177)
--	I10135 = NOT(g6249)
--	g7308 = NOT(I11572)
--	g8192 = NOT(I13117)
--	g2958 = NOT(I6163)
--	g8085 = NOT(g7932)
--	g10074 = NOT(I15299)
--	g5094 = NOT(I8462)
--	I13347 = NOT(g8122)
--	g2176 = NOT(g82)
--	g9026 = NOT(I14415)
--	g8485 = NOT(g8341)
--	g4184 = NOT(I7369)
--	g5494 = NOT(g4412)
--	g3750 = NOT(I6941)
--	g2005 = NOT(g928)
--	g7883 = NOT(g7689)
--	I7043 = NOT(g2908)
--	g4384 = NOT(I7707)
--	I9141 = NOT(g5402)
--	I9860 = NOT(g5405)
--	g5567 = NOT(I8982)
--	g4339 = NOT(g4144)
--	I9341 = NOT(g5013)
--	g10238 = NOT(g10191)
--	I16169 = NOT(g10448)
--	I9525 = NOT(g5001)
--	I14361 = NOT(g8951)
--	g2829 = NOT(I5943)
--	g11619 = NOT(I17675)
--	g2765 = NOT(g2184)
--	g9821 = NOT(I14964)
--	g11502 = NOT(I17525)
--	g7758 = NOT(I12439)
--	I5916 = NOT(g2217)
--	I13236 = NOT(g8245)
--	g7066 = NOT(I11275)
--	g7589 = NOT(I12099)
--	g4424 = NOT(g3688)
--	g3040 = NOT(g2135)
--	g4737 = NOT(g3440)
--	I11351 = NOT(g6698)
--	I13952 = NOT(g8451)
--	g5593 = NOT(I9013)
--	g6112 = NOT(I9789)
--	I13351 = NOT(g8214)
--	g6218 = NOT(I9965)
--	g6267 = NOT(I10060)
--	g3440 = NOT(g3041)
--	g6312 = NOT(I10195)
--	g11618 = NOT(I17672)
--	g9984 = NOT(I15184)
--	I11821 = NOT(g7205)
--	g10176 = NOT(I15520)
--	g10185 = NOT(g10040)
--	g10675 = NOT(g10574)
--	I16479 = NOT(g10767)
--	g10092 = NOT(I15323)
--	I10048 = NOT(g5734)
--	I16363 = NOT(g10599)
--	I16217 = NOT(g10501)
--	g3323 = NOT(g2157)
--	I15278 = NOT(g10033)
--	g7571 = NOT(I12035)
--	g7365 = NOT(I11743)
--	g2733 = NOT(I5795)
--	g4077 = NOT(I7202)
--	g6001 = NOT(I9625)
--	g7048 = NOT(I11225)
--	g10154 = NOT(I15458)
--	g2270 = NOT(I5311)
--	I5798 = NOT(g2085)
--	I17240 = NOT(g11395)
--	g7711 = NOT(I12344)
--	g4523 = NOT(g3546)
--	I10221 = NOT(g6117)
--	I11790 = NOT(g7246)
--	g8520 = NOT(I13729)
--	g6293 = NOT(I10138)
--	g11469 = NOT(I17444)
--	g8219 = NOT(g7826)
--	g2225 = NOT(I5210)
--	g8640 = NOT(g8512)
--	g10935 = NOT(g10827)
--	g2610 = NOT(I5731)
--	g2073 = NOT(I4879)
--	g2796 = NOT(g2276)
--	g11468 = NOT(I17441)
--	g11039 = NOT(I16778)
--	I6851 = NOT(g2937)
--	g4205 = NOT(I7432)
--	I7697 = NOT(g3743)
--	I10613 = NOT(g6000)
--	I11873 = NOT(g6863)
--	g10883 = NOT(g10809)
--	I17755 = NOT(g11646)
--	g7333 = NOT(I11647)
--	g9106 = NOT(I14439)
--	I7210 = NOT(g2798)
--	g7774 = NOT(I12487)
--	g5521 = NOT(g4530)
--	g3528 = NOT(g3164)
--	g8958 = NOT(I14323)
--	I16580 = NOT(g10826)
--	I17770 = NOT(g11649)
--	g11038 = NOT(I16775)
--	g5050 = NOT(I8429)
--	g2124 = NOT(I5050)
--	g3351 = NOT(I6535)
--	g5641 = NOT(I9084)
--	I17563 = NOT(g11492)
--	g2980 = NOT(g1983)
--	g6727 = NOT(g5997)
--	g8376 = NOT(I13478)
--	I5632 = NOT(g932)
--	I5095 = NOT(g37)
--	I6260 = NOT(g2025)
--	g2069 = NOT(I4869)
--	I9111 = NOT(g5596)
--	g7196 = NOT(I11420)
--	g4551 = NOT(g3946)
--	I15601 = NOT(g10173)
--	I9311 = NOT(g4915)
--	I15187 = NOT(g9968)
--	g7803 = NOT(I12574)
--	I12248 = NOT(g7098)
--	I13209 = NOT(g8198)
--	g4499 = NOT(g3546)
--	I8848 = NOT(g4490)
--	g2540 = NOT(I5655)
--	g7538 = NOT(I11950)
--	I13834 = NOT(g8488)
--	I5579 = NOT(g1197)
--	g7780 = NOT(I12505)
--	g5724 = NOT(I9268)
--	g9027 = NOT(I14418)
--	g2206 = NOT(I5171)
--	I12779 = NOT(g7608)
--	g10729 = NOT(g10630)
--	g6703 = NOT(I10678)
--	I9174 = NOT(g4903)
--	I5719 = NOT(g2072)
--	g10577 = NOT(g10526)
--	I17767 = NOT(g11648)
--	g7509 = NOT(I11889)
--	g9427 = NOT(g9079)
--	I10033 = NOT(g5693)
--	I7820 = NOT(g3811)
--	I10234 = NOT(g6114)
--	g4754 = NOT(g3440)
--	I16531 = NOT(g10720)
--	g10439 = NOT(g10334)
--	I11021 = NOT(g6398)
--	I12081 = NOT(g6934)
--	g5878 = NOT(g5309)
--	g6932 = NOT(I11058)
--	g7662 = NOT(I12279)
--	g4273 = NOT(g4013)
--	I16178 = NOT(g10490)
--	I12786 = NOT(g7622)
--	I17633 = NOT(g11578)
--	g5658 = NOT(I9135)
--	g5777 = NOT(I9365)
--	I10795 = NOT(g6123)
--	I13726 = NOT(g8375)
--	g7467 = NOT(g7148)
--	g1990 = NOT(g774)
--	I6118 = NOT(g2248)
--	g8225 = NOT(g7826)
--	I17191 = NOT(g11315)
--	I17719 = NOT(g11623)
--	I11614 = NOT(g6838)
--	g8610 = NOT(g8483)
--	I6367 = NOT(g2045)
--	I9180 = NOT(g4905)
--	I12647 = NOT(g7711)
--	I16676 = NOT(g10798)
--	I16685 = NOT(g10785)
--	I11436 = NOT(g6488)
--	I9380 = NOT(g5013)
--	g10349 = NOT(I15811)
--	g9345 = NOT(I14540)
--	I16953 = NOT(g11082)
--	I13436 = NOT(g8187)
--	I9591 = NOT(g5095)
--	I16373 = NOT(g10593)
--	g4444 = NOT(I7800)
--	g8473 = NOT(I13669)
--	g2199 = NOT(g48)
--	g11410 = NOT(I17271)
--	g2399 = NOT(g605)
--	g9763 = NOT(I14906)
--	g7093 = NOT(I11326)
--	I12999 = NOT(g7844)
--	g3372 = NOT(g3121)
--	I10514 = NOT(g6154)
--	I12380 = NOT(g7204)
--	g10906 = NOT(I16670)
--	I15479 = NOT(g10091)
--	I13320 = NOT(g8096)
--	g10083 = NOT(I15311)
--	I9020 = NOT(g4773)
--	g8124 = NOT(g8011)
--	g10284 = NOT(g10167)
--	g7256 = NOT(I11489)
--	g8980 = NOT(I14361)
--	g7816 = NOT(I12613)
--	g8324 = NOT(I13354)
--	g11479 = NOT(I17470)
--	I6193 = NOT(g2155)
--	I11593 = NOT(g6830)
--	g3143 = NOT(I6363)
--	g11363 = NOT(I17188)
--	g3343 = NOT(g2779)
--	I11122 = NOT(g6450)
--	g2797 = NOT(g2524)
--	I13122 = NOT(g7966)
--	I6549 = NOT(g2838)
--	g4543 = NOT(g3946)
--	I10421 = NOT(g5826)
--	I11464 = NOT(g6443)
--	g3566 = NOT(I6738)
--	I6971 = NOT(g2882)
--	g6716 = NOT(g5949)
--	I14421 = NOT(g8944)
--	g2245 = NOT(I5254)
--	g6149 = NOT(I9866)
--	g3988 = NOT(g3121)
--	I6686 = NOT(g3015)
--	g6349 = NOT(I10258)
--	g7847 = NOT(I12638)
--	g3693 = NOT(g2920)
--	I11034 = NOT(g6629)
--	I10012 = NOT(g5543)
--	g3334 = NOT(I6517)
--	I5725 = NOT(g2079)
--	g7685 = NOT(g7148)
--	g7197 = NOT(I11423)
--	I11641 = NOT(g6960)
--	I11797 = NOT(g6852)
--	g5997 = NOT(I9617)
--	I15580 = NOT(g10155)
--	I13797 = NOT(g8473)
--	I6598 = NOT(g2623)
--	g7021 = NOT(I11162)
--	g4729 = NOT(g3586)
--	g4961 = NOT(I8333)
--	g7421 = NOT(I11807)
--	g10139 = NOT(I15415)
--	g2344 = NOT(I5410)
--	I8211 = NOT(g3566)
--	I9905 = NOT(g5300)
--	g6398 = NOT(I10302)
--	I10541 = NOT(g6176)
--	I6121 = NOT(g2121)
--	g1963 = NOT(g110)
--	I17324 = NOT(g11347)
--	g7263 = NOT(I11498)
--	I14473 = NOT(g8921)
--	g2207 = NOT(I5174)
--	g10138 = NOT(I15412)
--	I17701 = NOT(g11617)
--	I10789 = NOT(g5867)
--	I12448 = NOT(g7530)
--	I13409 = NOT(g8141)
--	I17534 = NOT(g11495)
--	g3792 = NOT(I7017)
--	g5353 = NOT(I8820)
--	g8849 = NOT(g8745)
--	g2259 = NOT(I5292)
--	g6241 = NOT(I9992)
--	g2819 = NOT(g2159)
--	I11408 = NOT(g6405)
--	I12505 = NOT(g7728)
--	I11635 = NOT(g6947)
--	I10724 = NOT(g6096)
--	g11084 = NOT(I16863)
--	g4885 = NOT(I8228)
--	g4414 = NOT(I7752)
--	I10325 = NOT(g6003)
--	g11110 = NOT(g10974)
--	g3621 = NOT(I6754)
--	I6938 = NOT(g2854)
--	I7668 = NOT(g3733)
--	g2852 = NOT(I5982)
--	I7840 = NOT(g3431)
--	I16543 = NOT(g10747)
--	g10852 = NOT(g10740)
--	g8781 = NOT(I14080)
--	I8614 = NOT(g4414)
--	I10920 = NOT(g6733)
--	I10535 = NOT(g5867)
--	I12026 = NOT(g7119)
--	I10434 = NOT(g5843)
--	g11179 = NOT(I16938)
--	g2701 = NOT(g2040)
--	g3113 = NOT(I6343)
--	g7562 = NOT(g6984)
--	I14358 = NOT(g8950)
--	I7390 = NOT(g4087)
--	I10828 = NOT(g6708)
--	I10946 = NOT(g6548)
--	g8797 = NOT(I14116)
--	g6644 = NOT(I10601)
--	g4513 = NOT(g3546)
--	g7631 = NOT(I12235)
--	I5171 = NOT(g1419)
--	g7723 = NOT(I12354)
--	g6119 = NOT(I9810)
--	I9973 = NOT(g5502)
--	g7817 = NOT(I12616)
--	g5901 = NOT(g5361)
--	I4920 = NOT(g260)
--	g8291 = NOT(I13227)
--	g11373 = NOT(I17198)
--	g3094 = NOT(I6302)
--	g6258 = NOT(I10033)
--	g4178 = NOT(I7351)
--	g4436 = NOT(g3638)
--	g6818 = NOT(I10864)
--	g4679 = NOT(g4013)
--	g11654 = NOT(I17764)
--	g4378 = NOT(I7697)
--	g7605 = NOT(I12165)
--	g5511 = NOT(I8934)
--	I11575 = NOT(g6823)
--	g3518 = NOT(g3164)
--	I10682 = NOT(g6051)
--	g10576 = NOT(g10524)
--	I9040 = NOT(g4794)
--	g8144 = NOT(I13027)
--	g8344 = NOT(I13412)
--	g6717 = NOT(I10706)
--	I9440 = NOT(g5078)
--	g11417 = NOT(I17302)
--	I13711 = NOT(g8342)
--	I16814 = NOT(g10910)
--	I12433 = NOT(g7657)
--	g4335 = NOT(I7612)
--	I9123 = NOT(g4890)
--	I11109 = NOT(g6464)
--	g7751 = NOT(I12418)
--	g4182 = NOT(I7363)
--	I9323 = NOT(g5620)
--	I13109 = NOT(g7981)
--	g4288 = NOT(g4130)
--	I11537 = NOT(g7144)
--	g4382 = NOT(g3638)
--	I16772 = NOT(g10887)
--	g3776 = NOT(g2579)
--	g6893 = NOT(I10991)
--	g5574 = NOT(g4300)
--	g5864 = NOT(I9483)
--	g10200 = NOT(g10169)
--	g8694 = NOT(I13975)
--	g2825 = NOT(I5935)
--	g2650 = NOT(g2006)
--	g10608 = NOT(I16283)
--	g10115 = NOT(I15353)
--	g6386 = NOT(I10282)
--	g7585 = NOT(I12081)
--	I17447 = NOT(g11457)
--	I5684 = NOT(g572)
--	I8061 = NOT(g3381)
--	g4805 = NOT(g3337)
--	I7163 = NOT(g2643)
--	I5963 = NOT(g2179)
--	I7810 = NOT(g3799)
--	g7041 = NOT(g6427)
--	I7363 = NOT(g4005)
--	I16638 = NOT(g10863)
--	g2008 = NOT(g971)
--	I13606 = NOT(g8311)
--	I12971 = NOT(g8039)
--	I11303 = NOT(g6526)
--	g6274 = NOT(I10081)
--	I7432 = NOT(g3663)
--	g6426 = NOT(I10340)
--	g11423 = NOT(I17324)
--	g2336 = NOT(g1900)
--	I16416 = NOT(g10664)
--	I12369 = NOT(g7189)
--	I9875 = NOT(g5278)
--	I7453 = NOT(g3708)
--	g6170 = NOT(g5426)
--	I14506 = NOT(g8923)
--	g7673 = NOT(I12296)
--	I9655 = NOT(g5173)
--	g6125 = NOT(I9822)
--	I5707 = NOT(g2418)
--	g8886 = NOT(I14228)
--	g3521 = NOT(g3164)
--	g8951 = NOT(I14306)
--	I16510 = NOT(g10712)
--	g5262 = NOT(g4353)
--	g3050 = NOT(I6260)
--	I11091 = NOT(g6657)
--	g10973 = NOT(I16720)
--	g5736 = NOT(I9296)
--	g6984 = NOT(g6382)
--	g6280 = NOT(I10099)
--	g6939 = NOT(I11071)
--	g7669 = NOT(I12286)
--	I17246 = NOT(g11341)
--	g11543 = NOT(g11519)
--	g3996 = NOT(g3144)
--	g10184 = NOT(g10039)
--	I12412 = NOT(g7520)
--	I8403 = NOT(g4264)
--	g10674 = NOT(g10584)
--	g8314 = NOT(I13326)
--	g5623 = NOT(I9053)
--	g7772 = NOT(I12481)
--	I7157 = NOT(g3015)
--	g7058 = NOT(I11255)
--	I12133 = NOT(g6870)
--	I5957 = NOT(g2178)
--	I7357 = NOT(g4077)
--	g2122 = NOT(I5044)
--	g2228 = NOT(g28)
--	g7531 = NOT(I11929)
--	g4095 = NOT(I7233)
--	g9554 = NOT(I14697)
--	g8870 = NOT(I14182)
--	g2322 = NOT(I5378)
--	I10927 = NOT(g6755)
--	g7458 = NOT(g7123)
--	g5889 = NOT(I9514)
--	I12229 = NOT(g7070)
--	I6962 = NOT(g2791)
--	g4495 = NOT(I7886)
--	I9839 = NOT(g5226)
--	g2230 = NOT(g704)
--	g4437 = NOT(g3345)
--	g4102 = NOT(I7244)
--	I17591 = NOT(g11514)
--	g4208 = NOT(I7441)
--	g7890 = NOT(g7479)
--	g8650 = NOT(I13933)
--	I13840 = NOT(g8488)
--	I16586 = NOT(g10850)
--	g3379 = NOT(g3121)
--	I15568 = NOT(g10094)
--	g10934 = NOT(g10827)
--	g6106 = NOT(I9773)
--	g5175 = NOT(g4682)
--	g6306 = NOT(I10177)
--	g7505 = NOT(g7148)
--	g3878 = NOT(g2920)
--	g11242 = NOT(g11112)
--	I5098 = NOT(g38)
--	g8008 = NOT(I12846)
--	I10240 = NOT(g5937)
--	g7011 = NOT(g6503)
--	g4719 = NOT(g3586)
--	g10692 = NOT(I16363)
--	g5651 = NOT(I9114)
--	I6587 = NOT(g2620)
--	I10648 = NOT(g6030)
--	I15814 = NOT(g10202)
--	g8336 = NOT(I13388)
--	I14903 = NOT(g9507)
--	I5833 = NOT(g2103)
--	g6387 = NOT(g6121)
--	g5285 = NOT(g4355)
--	g6461 = NOT(I10391)
--	I15807 = NOT(g10284)
--	I15974 = NOT(g10411)
--	I8858 = NOT(g4506)
--	g2550 = NOT(g1834)
--	g7074 = NOT(I11299)
--	I16720 = NOT(g10854)
--	g3271 = NOT(I6443)
--	g10400 = NOT(g10348)
--	g2845 = NOT(g2168)
--	I9282 = NOT(g5633)
--	I15639 = NOT(g10179)
--	I10563 = NOT(g6043)
--	I5584 = NOT(g1200)
--	g10214 = NOT(I15586)
--	g9490 = NOT(g9324)
--	g9823 = NOT(I14970)
--	g2195 = NOT(g83)
--	g4265 = NOT(g3664)
--	I15293 = NOT(g10001)
--	I9988 = NOT(g5526)
--	g6427 = NOT(I10343)
--	I12627 = NOT(g7697)
--	g2395 = NOT(g231)
--	g2891 = NOT(I6055)
--	g5184 = NOT(g4682)
--	g2337 = NOT(I5395)
--	I11483 = NOT(g6567)
--	g2913 = NOT(I6088)
--	g10329 = NOT(I15775)
--	g10207 = NOT(g10186)
--	g4442 = NOT(g3638)
--	I6985 = NOT(g2890)
--	g6904 = NOT(I11008)
--	g6200 = NOT(I9935)
--	g11638 = NOT(I17724)
--	g10539 = NOT(I16184)
--	g4786 = NOT(I8154)
--	g6046 = NOT(I9669)
--	g8065 = NOT(I12913)
--	g3799 = NOT(I7022)
--	I8315 = NOT(g4788)
--	I8811 = NOT(g4465)
--	g6446 = NOT(I10370)
--	g8122 = NOT(I12981)
--	g3981 = NOT(I7118)
--	g8465 = NOT(g8289)
--	g9529 = NOT(I14672)
--	g4164 = NOT(I7311)
--	g10538 = NOT(I16181)
--	g4233 = NOT(g3698)
--	g5424 = NOT(I8865)
--	g9348 = NOT(I14549)
--	I11326 = NOT(g6660)
--	I13949 = NOT(g8451)
--	g6403 = NOT(g6128)
--	I13326 = NOT(g8203)
--	I9804 = NOT(g5417)
--	g6145 = NOT(I9860)
--	g2859 = NOT(I5995)
--	g3997 = NOT(I7131)
--	I15510 = NOT(g10035)
--	g9355 = NOT(I14570)
--	I9792 = NOT(g5403)
--	I6832 = NOT(g2909)
--	g4454 = NOT(g3914)
--	g8033 = NOT(I12875)
--	g11510 = NOT(I17549)
--	g6191 = NOT(g5446)
--	g7569 = NOT(I12029)
--	g5672 = NOT(I9177)
--	g4296 = NOT(I7559)
--	I11904 = NOT(g6902)
--	I10633 = NOT(g6015)
--	I10898 = NOT(g6735)
--	g5231 = NOT(g4640)
--	I17318 = NOT(g11340)
--	g3332 = NOT(I6513)
--	I11252 = NOT(g6542)
--	g10241 = NOT(g10192)
--	g9260 = NOT(g8892)
--	g6695 = NOT(I10666)
--	I10719 = NOT(g6003)
--	I13621 = NOT(g8315)
--	g5643 = NOT(I9090)
--	g3353 = NOT(g3121)
--	I7735 = NOT(g3759)
--	I6507 = NOT(g2808)
--	I14191 = NOT(g8795)
--	g8096 = NOT(I12953)
--	g2248 = NOT(g99)
--	g11578 = NOT(I17616)
--	g2342 = NOT(I5406)
--	I7782 = NOT(g3775)
--	g6107 = NOT(I9776)
--	I17540 = NOT(g11498)
--	I12857 = NOT(g7638)
--	g11014 = NOT(I16735)
--	g6307 = NOT(I10180)
--	g3744 = NOT(g3307)
--	g6536 = NOT(I10456)
--	I4883 = NOT(g581)
--	g5205 = NOT(g4366)
--	I15586 = NOT(g10159)
--	I8880 = NOT(g4537)
--	g2255 = NOT(I5276)
--	I5728 = NOT(g2084)
--	g7688 = NOT(g7148)
--	I12793 = NOT(g7619)
--	g2481 = NOT(g882)
--	I9202 = NOT(g4915)
--	g8195 = NOT(I13122)
--	g7976 = NOT(I12776)
--	g8137 = NOT(I13010)
--	g8891 = NOT(I14239)
--	g8337 = NOT(I13391)
--	g10235 = NOT(g10189)
--	g4012 = NOT(I7154)
--	I11183 = NOT(g6507)
--	I16193 = NOT(g10485)
--	g11442 = NOT(I17377)
--	g2097 = NOT(I4935)
--	I12765 = NOT(g7638)
--	g10683 = NOT(g10612)
--	g5742 = NOT(I9308)
--	g2726 = NOT(g2021)
--	g4412 = NOT(I7746)
--	I11397 = NOT(g6713)
--	I13397 = NOT(g8138)
--	g2154 = NOT(I5067)
--	g6016 = NOT(I9632)
--	I12690 = NOT(g7555)
--	g4189 = NOT(I7384)
--	I5070 = NOT(g1194)
--	g2960 = NOT(I6173)
--	I10861 = NOT(g6694)
--	I10573 = NOT(g5980)
--	I9567 = NOT(g5556)
--	g8807 = NOT(I14140)
--	I14573 = NOT(g9029)
--	g4888 = NOT(I8237)
--	g7126 = NOT(I11367)
--	I13933 = NOT(g8505)
--	I17377 = NOT(g11412)
--	g7326 = NOT(I11626)
--	I10045 = NOT(g5727)
--	g6115 = NOT(I9798)
--	g6251 = NOT(I10012)
--	g4171 = NOT(I7330)
--	g6315 = NOT(I10204)
--	g6811 = NOT(I10843)
--	I15275 = NOT(g9994)
--	g4371 = NOT(I7674)
--	I14045 = NOT(g8603)
--	I17739 = NOT(g11641)
--	g4429 = NOT(I7779)
--	g4787 = NOT(g3423)
--	I8982 = NOT(g4728)
--	g11041 = NOT(I16784)
--	g10882 = NOT(I16616)
--	g5754 = NOT(I9332)
--	I9776 = NOT(g5353)
--	I10099 = NOT(g5800)
--	I16475 = NOT(g10765)
--	g6447 = NOT(g6166)
--	I10388 = NOT(g5830)
--	I8234 = NOT(g4232)
--	g7760 = NOT(I12445)
--	I14388 = NOT(g8924)
--	I8328 = NOT(g4801)
--	I17146 = NOT(g11305)
--	I16863 = NOT(g10972)
--	g3092 = NOT(g2181)
--	I14701 = NOT(g9291)
--	I10251 = NOT(g6126)
--	I14534 = NOT(g9290)
--	g4281 = NOT(g3586)
--	I9965 = NOT(g5493)
--	g5613 = NOT(g4840)
--	g6874 = NOT(I10958)
--	g8142 = NOT(I13023)
--	g2112 = NOT(g639)
--	g8342 = NOT(I13406)
--	g2218 = NOT(g85)
--	I15983 = NOT(g10414)
--	g2267 = NOT(I5304)
--	I17698 = NOT(g11616)
--	g11035 = NOT(I16766)
--	g8255 = NOT(g7986)
--	g8081 = NOT(g8000)
--	g8481 = NOT(g8324)
--	g2001 = NOT(g814)
--	g7608 = NOT(I12174)
--	g7924 = NOT(g7470)
--	I5406 = NOT(g898)
--	g7220 = NOT(I11456)
--	g5572 = NOT(I8989)
--	g5862 = NOT(I9479)
--	I12245 = NOT(g7093)
--	g7779 = NOT(I12502)
--	I4780 = NOT(g872)
--	I6040 = NOT(g2216)
--	g6595 = NOT(I10563)
--	g10584 = NOT(g10522)
--	I15517 = NOT(g10051)
--	I13574 = NOT(g8360)
--	g2329 = NOT(I5383)
--	g8354 = NOT(I13442)
--	I14140 = NOT(g8717)
--	g7023 = NOT(I11166)
--	I7952 = NOT(g3664)
--	g4963 = NOT(I8337)
--	g10206 = NOT(g10178)
--	I5801 = NOT(g1984)
--	I7276 = NOT(g2861)
--	g9670 = NOT(I14799)
--	I16781 = NOT(g10893)
--	g4791 = NOT(I8161)
--	g7977 = NOT(I12779)
--	g2828 = NOT(I5940)
--	g6272 = NOT(I10075)
--	I16236 = NOT(g10535)
--	g3262 = NOT(I6432)
--	g2727 = NOT(g2022)
--	g3736 = NOT(I6924)
--	g5534 = NOT(g4545)
--	g5729 = NOT(I9279)
--	g7361 = NOT(I11731)
--	g10114 = NOT(I15350)
--	I16175 = NOT(g10488)
--	g9813 = NOT(I14948)
--	I15193 = NOT(g9968)
--	g6417 = NOT(g6136)
--	I13051 = NOT(g8060)
--	I15362 = NOT(g9987)
--	g6935 = NOT(I11065)
--	g11193 = NOT(g11112)
--	g7051 = NOT(I11232)
--	g10107 = NOT(I15341)
--	I11756 = NOT(g7191)
--	g2221 = NOT(I5198)
--	g3076 = NOT(I6282)
--	I13592 = NOT(g8362)
--	g8783 = NOT(g8746)
--	I15523 = NOT(g10058)
--	g7327 = NOT(I11629)
--	I12232 = NOT(g7072)
--	I6528 = NOT(g3274)
--	I16264 = NOT(g10557)
--	g8979 = NOT(I14358)
--	I16790 = NOT(g10900)
--	I8490 = NOT(g4526)
--	g4201 = NOT(I7420)
--	I6648 = NOT(g2635)
--	g8218 = NOT(g7826)
--	I9658 = NOT(g5150)
--	g8312 = NOT(I13320)
--	I7546 = NOT(g4105)
--	g6128 = NOT(I9829)
--	g6629 = NOT(I10584)
--	g5885 = NOT(g5361)
--	g10345 = NOT(I15801)
--	g7999 = NOT(I12825)
--	g7146 = NOT(I11391)
--	g5660 = NOT(I9141)
--	I5445 = NOT(g922)
--	g6330 = NOT(I10221)
--	g7346 = NOT(I11686)
--	I10162 = NOT(g5943)
--	g7633 = NOT(I12239)
--	g4049 = NOT(g3144)
--	g3375 = NOT(I6569)
--	g8001 = NOT(I12829)
--	I12261 = NOT(g7078)
--	g4449 = NOT(g4144)
--	g3722 = NOT(I6894)
--	I8456 = NOT(g4472)
--	g7103 = NOT(I11338)
--	g5903 = NOT(I9536)
--	g4575 = NOT(g3880)
--	g10848 = NOT(I16546)
--	g11475 = NOT(I17466)
--	g8293 = NOT(I13233)
--	g8129 = NOT(g8015)
--	I6010 = NOT(g2256)
--	g2068 = NOT(I4866)
--	I11152 = NOT(g6469)
--	g8329 = NOT(I13367)
--	g10141 = NOT(I15421)
--	g7696 = NOT(g7148)
--	g10804 = NOT(I16514)
--	g6800 = NOT(I10810)
--	g4098 = NOT(I7240)
--	g3500 = NOT(I6690)
--	I15437 = NOT(g10050)
--	I16209 = NOT(g10452)
--	I8851 = NOT(g4498)
--	I11731 = NOT(g7021)
--	g8828 = NOT(g8744)
--	g11437 = NOT(I17362)
--	g2677 = NOT(g2034)
--	g10263 = NOT(g10127)
--	g7753 = NOT(I12424)
--	I9981 = NOT(g5514)
--	g8727 = NOT(g8592)
--	g5679 = NOT(I9194)
--	g7508 = NOT(g6950)
--	g3384 = NOT(g3143)
--	g10332 = NOT(I15782)
--	g6213 = NOT(g5426)
--	g8592 = NOT(I13837)
--	g7944 = NOT(g7410)
--	I15347 = NOT(g9995)
--	g7072 = NOT(I11293)
--	I15253 = NOT(g9987)
--	g10135 = NOT(I15403)
--	I12445 = NOT(g7521)
--	g11347 = NOT(I17164)
--	g4896 = NOT(I8253)
--	I7906 = NOT(g3907)
--	g2349 = NOT(I5421)
--	g7043 = NOT(I11214)
--	I12499 = NOT(g7725)
--	I11405 = NOT(g6627)
--	g5288 = NOT(g4438)
--	g9341 = NOT(I14528)
--	g3424 = NOT(g2896)
--	I9132 = NOT(g4893)
--	g10361 = NOT(g10268)
--	g3737 = NOT(g2834)
--	g7443 = NOT(I11841)
--	I9332 = NOT(g4935)
--	g9525 = NOT(g9257)
--	I9153 = NOT(g5027)
--	I9680 = NOT(g5194)
--	I10147 = NOT(g5697)
--	I6343 = NOT(g1963)
--	I10355 = NOT(g6003)
--	g7116 = NOT(I11351)
--	g5805 = NOT(I9409)
--	g5916 = NOT(I9550)
--	g7316 = NOT(I11596)
--	g2198 = NOT(g668)
--	I6282 = NOT(g2231)
--	g4268 = NOT(I7523)
--	I7771 = NOT(g3418)
--	I16607 = NOT(g10787)
--	g2855 = NOT(I5989)
--	g4362 = NOT(I7651)
--	I11929 = NOT(g6901)
--	I14355 = NOT(g8948)
--	I12989 = NOT(g8043)
--	g11351 = NOT(I17170)
--	g3077 = NOT(g2213)
--	g5422 = NOT(g4470)
--	g7034 = NOT(I11191)
--	I10825 = NOT(g6588)
--	g4419 = NOT(I7763)
--	I9744 = NOT(g5263)
--	I12056 = NOT(g6929)
--	I10370 = NOT(g5857)
--	g6166 = NOT(I9893)
--	g8624 = NOT(g8486)
--	g3523 = NOT(g2971)
--	I14370 = NOT(g8954)
--	g8953 = NOT(I14312)
--	I10858 = NOT(g6688)
--	I13020 = NOT(g8049)
--	I13583 = NOT(g8344)
--	g4452 = NOT(g3365)
--	I8872 = NOT(g4529)
--	I15063 = NOT(g9699)
--	g2241 = NOT(g722)
--	g7147 = NOT(I11394)
--	g6056 = NOT(g5426)
--	g5947 = NOT(I9585)
--	g7347 = NOT(I11689)
--	g11063 = NOT(g10974)
--	I11046 = NOT(g6635)
--	I10996 = NOT(g6786)
--	I12271 = NOT(g7218)
--	g7681 = NOT(g7148)
--	g6649 = NOT(I10610)
--	I8989 = NOT(g4746)
--	g8677 = NOT(I13962)
--	g110 = NOT(I4786)
--	I10367 = NOT(g6234)
--	I10394 = NOT(g5824)
--	I9901 = NOT(g5557)
--	g7697 = NOT(g7101)
--	I14367 = NOT(g8953)
--	I14394 = NOT(g8884)
--	I16641 = NOT(g10864)
--	g3742 = NOT(I6929)
--	g7914 = NOT(g7651)
--	g8576 = NOT(I13819)
--	g2524 = NOT(g986)
--	g7210 = NOT(I11440)
--	g4728 = NOT(I8080)
--	I16292 = NOT(g10551)
--	g2644 = NOT(g1990)
--	g6698 = NOT(I10671)
--	g4730 = NOT(g3546)
--	g8716 = NOT(g8576)
--	I17546 = NOT(g11500)
--	g8149 = NOT(I13036)
--	g10947 = NOT(I16708)
--	g4504 = NOT(I7899)
--	I11357 = NOT(g6594)
--	g6964 = NOT(g6509)
--	g8349 = NOT(I13427)
--	g2119 = NOT(I5031)
--	g5095 = NOT(I8465)
--	g6260 = NOT(I10039)
--	g5037 = NOT(I8414)
--	I13357 = NOT(g8125)
--	I12199 = NOT(g7278)
--	g4185 = NOT(I7372)
--	I7244 = NOT(g3226)
--	g9311 = NOT(I14506)
--	g11422 = NOT(I17321)
--	I11743 = NOT(g7035)
--	I13105 = NOT(g7929)
--	g5653 = NOT(I9120)
--	g4385 = NOT(I7710)
--	g7413 = NOT(g7197)
--	g5102 = NOT(I8476)
--	g2258 = NOT(I5289)
--	I14319 = NOT(g8816)
--	g2352 = NOT(I5430)
--	g2818 = NOT(I5922)
--	I7140 = NOT(g2641)
--	g6063 = NOT(g5446)
--	I12529 = NOT(g7589)
--	I5940 = NOT(g2175)
--	g2867 = NOT(I6007)
--	I16635 = NOT(g10862)
--	g10463 = NOT(I15980)
--	g11208 = NOT(g11077)
--	g4470 = NOT(I7843)
--	g8198 = NOT(I13131)
--	g4897 = NOT(I8256)
--	g8747 = NOT(I14040)
--	I7478 = NOT(g3566)
--	g5719 = NOT(I9259)
--	g4425 = NOT(I7771)
--	I12843 = NOT(g7683)
--	I15542 = NOT(g10065)
--	g10972 = NOT(I16717)
--	g10033 = NOT(I15235)
--	I5388 = NOT(g889)
--	g10234 = NOT(g10188)
--	I7435 = NOT(g3459)
--	g7936 = NOT(g7712)
--	g11542 = NOT(g11519)
--	g11453 = NOT(I17416)
--	g5752 = NOT(I9326)
--	I6094 = NOT(g2110)
--	I13803 = NOT(g8476)
--	g3044 = NOT(I6256)
--	g2211 = NOT(g153)
--	I14540 = NOT(g9310)
--	g6279 = NOT(I10096)
--	g2186 = NOT(g90)
--	g7317 = NOT(I11599)
--	g6720 = NOT(I10713)
--	I8253 = NOT(g4637)
--	g6118 = NOT(I9807)
--	g3983 = NOT(g3222)
--	g11614 = NOT(I17662)
--	g7601 = NOT(I12153)
--	I5430 = NOT(g916)
--	g5265 = NOT(g4362)
--	g11436 = NOT(I17359)
--	g3862 = NOT(g2920)
--	g5042 = NOT(g4840)
--	I15320 = NOT(g10013)
--	g9832 = NOT(I14989)
--	g6652 = NOT(I10613)
--	g4678 = NOT(g3546)
--	g6057 = NOT(g5446)
--	g6843 = NOT(I10901)
--	I15530 = NOT(g10107)
--	g11073 = NOT(g10913)
--	g4331 = NOT(I7606)
--	g3543 = NOT(g3101)
--	g2170 = NOT(g30)
--	g2614 = NOT(g1994)
--	g7775 = NOT(I12490)
--	g11593 = NOT(I17633)
--	g7922 = NOT(I12712)
--	g2125 = NOT(I5053)
--	g8319 = NOT(I13341)
--	g11346 = NOT(I17161)
--	I15565 = NOT(g10101)
--	g2821 = NOT(I5929)
--	g9507 = NOT(g9268)
--	I15464 = NOT(g10094)
--	I6965 = NOT(g2880)
--	I10120 = NOT(g6248)
--	g4766 = NOT(g3440)
--	I11662 = NOT(g7033)
--	I10739 = NOT(g5942)
--	g4087 = NOT(I7220)
--	g4105 = NOT(I7249)
--	g8152 = NOT(I13043)
--	g10421 = NOT(g10331)
--	I16537 = NOT(g10721)
--	g8352 = NOT(I13436)
--	g4305 = NOT(g4013)
--	g6971 = NOT(g6517)
--	I13027 = NOT(g8051)
--	I12258 = NOT(g7103)
--	g3729 = NOT(I6907)
--	I6264 = NOT(g2118)
--	I16108 = NOT(g10383)
--	g6686 = NOT(I10651)
--	g10163 = NOT(I15485)
--	g8717 = NOT(I14010)
--	g11034 = NOT(I16763)
--	g7460 = NOT(g7148)
--	g7597 = NOT(I12133)
--	g5296 = NOT(g4444)
--	I11249 = NOT(g6541)
--	I5638 = NOT(g936)
--	I14645 = NOT(g9088)
--	I16283 = NOT(g10538)
--	g2083 = NOT(g139)
--	I6360 = NOT(g2261)
--	g4748 = NOT(g3546)
--	I16492 = NOT(g10773)
--	I13482 = NOT(g8193)
--	I5308 = NOT(g97)
--	I11710 = NOT(g7020)
--	g7784 = NOT(I12517)
--	I4992 = NOT(g1170)
--	g4755 = NOT(g3440)
--	g10541 = NOT(I16190)
--	I10698 = NOT(g5856)
--	g6121 = NOT(I9816)
--	I15409 = NOT(g10065)
--	I7002 = NOT(g2907)
--	g8186 = NOT(I13109)
--	g10473 = NOT(g10380)
--	g4226 = NOT(g3698)
--	I11204 = NOT(g6523)
--	g6670 = NOT(I10633)
--	I7402 = NOT(g4121)
--	g11409 = NOT(I17268)
--	I6996 = NOT(g2904)
--	g3946 = NOT(I7099)
--	I13779 = NOT(g8514)
--	I7236 = NOT(g3219)
--	I15635 = NOT(g10185)
--	I16982 = NOT(g11088)
--	g8599 = NOT(g8546)
--	g7995 = NOT(I12817)
--	g2790 = NOT(g2276)
--	g11408 = NOT(I17265)
--	g7079 = NOT(I11312)
--	g11635 = NOT(I17719)
--	I11778 = NOT(g7210)
--	g3903 = NOT(I7070)
--	g5012 = NOT(I8388)
--	g9100 = NOT(g8892)
--	g8274 = NOT(I13194)
--	I10427 = NOT(g5839)
--	g7479 = NOT(I11873)
--	g8426 = NOT(I13592)
--	g1994 = NOT(g794)
--	g4445 = NOT(I7803)
--	g6253 = NOT(I10018)
--	g2061 = NOT(g1828)
--	g2187 = NOT(g746)
--	g6938 = NOT(I11068)
--	g4173 = NOT(I7336)
--	g6813 = NOT(I10849)
--	g4373 = NOT(I7680)
--	I11786 = NOT(g7246)
--	I16796 = NOT(g11016)
--	g10535 = NOT(I16172)
--	g4491 = NOT(g3546)
--	g8125 = NOT(I12986)
--	g7190 = NOT(I11412)
--	g8325 = NOT(I13357)
--	I11647 = NOT(g6925)
--	g7390 = NOT(g6847)
--	I12878 = NOT(g7638)
--	g5888 = NOT(g5102)
--	I13945 = NOT(g8488)
--	I12171 = NOT(g6885)
--	g10121 = NOT(I15371)
--	g8984 = NOT(I14373)
--	g3436 = NOT(g3144)
--	g4369 = NOT(I7668)
--	g8280 = NOT(I13212)
--	I7556 = NOT(g4080)
--	g4602 = NOT(I8011)
--	g7501 = NOT(I11879)
--	I17450 = NOT(g11450)
--	g3378 = NOT(I6572)
--	g5787 = NOT(I9383)
--	I9424 = NOT(g4963)
--	I9795 = NOT(g5404)
--	I17315 = NOT(g11393)
--	g10344 = NOT(I15798)
--	I9737 = NOT(g5258)
--	g2904 = NOT(I6065)
--	g2200 = NOT(g92)
--	g6552 = NOT(g5733)
--	g7356 = NOT(I11716)
--	g2046 = NOT(g1845)
--	I17707 = NOT(g11619)
--	g4920 = NOT(I8293)
--	I5827 = NOT(g2271)
--	g2446 = NOT(g1400)
--	g4459 = NOT(I7820)
--	I17202 = NOT(g11322)
--	g3335 = NOT(I6520)
--	I13233 = NOT(g8265)
--	g8483 = NOT(g8332)
--	g4767 = NOT(I8123)
--	I7064 = NOT(g2984)
--	g11575 = NOT(g11561)
--	g2003 = NOT(g822)
--	g5281 = NOT(g4428)
--	g3382 = NOT(I6580)
--	I9077 = NOT(g4765)
--	I7899 = NOT(g3380)
--	g4535 = NOT(g3946)
--	I8358 = NOT(g4794)
--	I6611 = NOT(g2626)
--	I8506 = NOT(g4334)
--	g2345 = NOT(g1936)
--	g10173 = NOT(g10120)
--	I17070 = NOT(g11233)
--	g8106 = NOT(g7950)
--	g11109 = NOT(g10974)
--	g8306 = NOT(I13290)
--	g2763 = NOT(I5847)
--	g2191 = NOT(g1696)
--	g2391 = NOT(I5478)
--	g6586 = NOT(g5949)
--	I12919 = NOT(g8003)
--	I6799 = NOT(g2750)
--	I11932 = NOT(g6908)
--	g3749 = NOT(I6938)
--	g8790 = NOT(I14101)
--	I9205 = NOT(g5309)
--	g11108 = NOT(g10974)
--	g2695 = NOT(g2039)
--	g9666 = NOT(I14793)
--	g8061 = NOT(I12901)
--	g5684 = NOT(I9205)
--	I8275 = NOT(g4351)
--	I8311 = NOT(g4794)
--	g4415 = NOT(g3914)
--	g5639 = NOT(I9080)
--	I14127 = NOT(g8768)
--	I17384 = NOT(g11437)
--	g7810 = NOT(I12595)
--	g7363 = NOT(I11737)
--	g10134 = NOT(I15400)
--	I7295 = NOT(g3260)
--	I11961 = NOT(g7053)
--	I16553 = NOT(g10754)
--	g5109 = NOT(I8495)
--	g5791 = NOT(I9391)
--	g3798 = NOT(g3228)
--	I13448 = NOT(g8150)
--	I9099 = NOT(g5572)
--	g2159 = NOT(I5080)
--	g7432 = NOT(I11824)
--	I14490 = NOT(g8885)
--	g6141 = NOT(I9854)
--	g8622 = NOT(g8485)
--	g6570 = NOT(g5949)
--	g6860 = NOT(g6475)
--	g7053 = NOT(I11238)
--	I11505 = NOT(g6585)
--	g9351 = NOT(I14558)
--	I5662 = NOT(g563)
--	g9875 = NOT(I15036)
--	g8427 = NOT(I13595)
--	I5067 = NOT(g33)
--	g9530 = NOT(I14675)
--	g6710 = NOT(I10693)
--	g5808 = NOT(g5320)
--	I5418 = NOT(g907)
--	g2858 = NOT(I5992)
--	I12598 = NOT(g7628)
--	I7194 = NOT(g2629)
--	I14376 = NOT(g8959)
--	I14385 = NOT(g8890)
--	g4203 = NOT(I7426)
--	I8985 = NOT(g4733)
--	I13717 = NOT(g8354)
--	g11381 = NOT(I17206)
--	g4721 = NOT(g3546)
--	g2016 = NOT(g1361)
--	I13212 = NOT(g8195)
--	g2757 = NOT(I5837)
--	g8446 = NOT(I13636)
--	g7568 = NOT(I12026)
--	g5759 = NOT(I9341)
--	I9754 = NOT(g5271)
--	I10888 = NOT(g6333)
--	g8514 = NOT(I13711)
--	I6802 = NOT(g2751)
--	g3632 = NOT(I6799)
--	g3095 = NOT(g2482)
--	g3037 = NOT(g2135)
--	g8003 = NOT(I12835)
--	I14888 = NOT(g9454)
--	I16252 = NOT(g10515)
--	g3437 = NOT(I6654)
--	I12817 = NOT(g7692)
--	I9273 = NOT(g5091)
--	I10671 = NOT(g6045)
--	I17695 = NOT(g11614)
--	g3102 = NOT(g2482)
--	I4924 = NOT(g123)
--	g3208 = NOT(I6381)
--	I12322 = NOT(g7246)
--	g7912 = NOT(g7651)
--	g8145 = NOT(I13030)
--	g8345 = NOT(I13415)
--	g2251 = NOT(g731)
--	g2642 = NOT(g1988)
--	I12159 = NOT(g7243)
--	g7357 = NOT(I11719)
--	g2047 = NOT(g1857)
--	I12532 = NOT(g7594)
--	I12901 = NOT(g7984)
--	g8191 = NOT(I13114)
--	g10927 = NOT(g10827)
--	g9884 = NOT(I15063)
--	g6158 = NOT(I9883)
--	g3719 = NOT(g2920)
--	I12783 = NOT(g7590)
--	g11390 = NOT(I17219)
--	I13723 = NOT(g8359)
--	g5865 = NOT(I9486)
--	g8695 = NOT(I13978)
--	I5847 = NOT(g2275)
--	I6901 = NOT(g2818)
--	I11149 = NOT(g6468)
--	g2874 = NOT(I6022)
--	g7929 = NOT(g7519)
--	g3752 = NOT(I6947)
--	I16673 = NOT(g10782)
--	I11433 = NOT(g6424)
--	I16847 = NOT(g10886)
--	I11387 = NOT(g6672)
--	g5604 = NOT(I9032)
--	I13433 = NOT(g8181)
--	g5098 = NOT(g4840)
--	g2654 = NOT(g2012)
--	I11620 = NOT(g6840)
--	g4188 = NOT(I7381)
--	g5498 = NOT(I8919)
--	I9712 = NOT(g5230)
--	g6587 = NOT(g5827)
--	g4388 = NOT(I7719)
--	g10491 = NOT(I16108)
--	g10903 = NOT(g10809)
--	I11097 = NOT(g6748)
--	I5421 = NOT(g549)
--	g8359 = NOT(I13457)
--	g6111 = NOT(I9786)
--	g6275 = NOT(I10084)
--	g6311 = NOT(I10192)
--	g4216 = NOT(I7465)
--	g10604 = NOT(I16280)
--	g9343 = NOT(I14534)
--	g8858 = NOT(g8743)
--	g4671 = NOT(g3354)
--	g2880 = NOT(I6028)
--	g4428 = NOT(I7776)
--	g2537 = NOT(I5646)
--	I10546 = NOT(g5914)
--	g5896 = NOT(I9525)
--	g4430 = NOT(I7782)
--	I14546 = NOT(g9312)
--	I7438 = NOT(g3461)
--	g3164 = NOT(I6370)
--	g3364 = NOT(g3121)
--	I7009 = NOT(g2913)
--	I10024 = NOT(g5700)
--	I8204 = NOT(g3976)
--	I12631 = NOT(g7705)
--	g8115 = NOT(g7953)
--	g4564 = NOT(g3880)
--	g8251 = NOT(I13166)
--	g8315 = NOT(I13329)
--	g2612 = NOT(I5737)
--	I15326 = NOT(g10025)
--	g2017 = NOT(g1218)
--	g6284 = NOT(I10111)
--	g2243 = NOT(I5248)
--	g8447 = NOT(I13639)
--	I6580 = NOT(g3186)
--	g3770 = NOT(I6985)
--	g6239 = NOT(I9988)
--	g10794 = NOT(I16496)
--	I15536 = NOT(g10111)
--	g10395 = NOT(g10320)
--	g5419 = NOT(I8858)
--	g9804 = NOT(I14939)
--	g10262 = NOT(g10142)
--	g7683 = NOT(g7148)
--	g11040 = NOT(I16781)
--	g10899 = NOT(g10803)
--	g6591 = NOT(I10553)
--	I11412 = NOT(g6411)
--	g5052 = NOT(g4394)
--	I13412 = NOT(g8142)
--	I5101 = NOT(g1960)
--	g8874 = NOT(I14194)
--	g3532 = NOT(g3164)
--	g7778 = NOT(I12499)
--	g2234 = NOT(g87)
--	g6853 = NOT(I10917)
--	I10126 = NOT(g5682)
--	I10659 = NOT(g6038)
--	I16574 = NOT(g10821)
--	g2629 = NOT(g2001)
--	g4638 = NOT(g3354)
--	g2328 = NOT(g1882)
--	I12289 = NOT(g7142)
--	I6968 = NOT(g2881)
--	g6420 = NOT(I10334)
--	g11621 = NOT(I17681)
--	g2130 = NOT(I5057)
--	g10191 = NOT(I15551)
--	g2542 = NOT(g1868)
--	I8973 = NOT(g4488)
--	g2330 = NOT(g1891)
--	g7735 = NOT(I12384)
--	I16311 = NOT(g10584)
--	g4308 = NOT(g3863)
--	I11228 = NOT(g6471)
--	I17231 = NOT(g11303)
--	g7782 = NOT(I12511)
--	g6559 = NOT(g5758)
--	I12571 = NOT(g7509)
--	g3012 = NOT(I6247)
--	I11011 = NOT(g6340)
--	I5751 = NOT(g2296)
--	g8595 = NOT(I13840)
--	g6931 = NOT(I11055)
--	g5728 = NOT(I9276)
--	g5486 = NOT(g4395)
--	I10296 = NOT(g6242)
--	I11716 = NOT(g7026)
--	g5730 = NOT(I9282)
--	g5504 = NOT(g4419)
--	g7949 = NOT(g7422)
--	g4217 = NOT(I7468)
--	g11183 = NOT(I16950)
--	I8123 = NOT(g3630)
--	g3990 = NOT(g3121)
--	g2554 = NOT(I5672)
--	g4758 = NOT(g3586)
--	g4066 = NOT(I7191)
--	g8272 = NOT(I13188)
--	I16592 = NOT(g10781)
--	g4589 = NOT(I7996)
--	g5185 = NOT(g4682)
--	g11397 = NOT(I17234)
--	g5881 = NOT(g5361)
--	g7627 = NOT(I12223)
--	g9094 = NOT(g8892)
--	I5041 = NOT(g1179)
--	I9135 = NOT(g5198)
--	g4466 = NOT(I7833)
--	g1992 = NOT(g782)
--	g6905 = NOT(I11011)
--	g8978 = NOT(I14355)
--	I5441 = NOT(g919)
--	g3371 = NOT(g2837)
--	g11062 = NOT(g10937)
--	I10060 = NOT(g5752)
--	g2213 = NOT(g1110)
--	g11509 = NOT(I17546)
--	g7998 = NOT(I12822)
--	g10247 = NOT(I15639)
--	g4165 = NOT(g3164)
--	g4365 = NOT(g3880)
--	I13627 = NOT(g8326)
--	g5425 = NOT(g4300)
--	g10389 = NOT(g10307)
--	g10926 = NOT(g10827)
--	I10855 = NOT(g6685)
--	I13959 = NOT(g8451)
--	I13379 = NOT(g8133)
--	g11508 = NOT(I17543)
--	g4711 = NOT(I8061)
--	g6100 = NOT(I9759)
--	I11112 = NOT(g6445)
--	g8982 = NOT(I14367)
--	g11634 = NOT(I17716)
--	g10612 = NOT(I16286)
--	g6300 = NOT(I10159)
--	g7603 = NOT(I12159)
--	g4055 = NOT(g3144)
--	g7039 = NOT(I11204)
--	I9749 = NOT(g5266)
--	g10388 = NOT(g10305)
--	I8351 = NOT(g4794)
--	g8234 = NOT(g7826)
--	g2902 = NOT(I6061)
--	g7439 = NOT(I11833)
--	g8128 = NOT(I12993)
--	g8328 = NOT(I13364)
--	g7850 = NOT(I12647)
--	g10534 = NOT(I16169)
--	g10098 = NOT(I15332)
--	I17456 = NOT(g11453)
--	g4333 = NOT(g4144)
--	I7837 = NOT(g4158)
--	g8330 = NOT(I13370)
--	g10251 = NOT(g10195)
--	g10272 = NOT(g10168)
--	g2090 = NOT(I4920)
--	g4774 = NOT(I8136)
--	I7462 = NOT(g3721)
--	I9798 = NOT(g5415)
--	I13096 = NOT(g7925)
--	g2166 = NOT(I5101)
--	g6750 = NOT(I10759)
--	g9264 = NOT(I14477)
--	I6424 = NOT(g2462)
--	g7702 = NOT(g7079)
--	g4196 = NOT(I7405)
--	g5678 = NOT(I9191)
--	I10503 = NOT(g5858)
--	I16413 = NOT(g10663)
--	g10462 = NOT(I15977)
--	g4396 = NOT(I7735)
--	g3138 = NOT(I6356)
--	g8800 = NOT(I14123)
--	I14503 = NOT(g8920)
--	I8410 = NOT(g4283)
--	g2056 = NOT(I4859)
--	I16691 = NOT(g10788)
--	g9360 = NOT(I14579)
--	g3109 = NOT(g2482)
--	g3791 = NOT(I7014)
--	g2456 = NOT(g1397)
--	g7919 = NOT(g7512)
--	g10032 = NOT(I15232)
--	g2529 = NOT(I5638)
--	g2649 = NOT(g2005)
--	g10140 = NOT(I15418)
--	g4780 = NOT(g3440)
--	I8839 = NOT(g4484)
--	g6040 = NOT(I9655)
--	g2348 = NOT(I5418)
--	I6077 = NOT(g2349)
--	g11574 = NOT(g11561)
--	g11452 = NOT(I17413)
--	g11047 = NOT(I16802)
--	g5682 = NOT(I9199)
--	g5766 = NOT(I9346)
--	g5105 = NOT(I8487)
--	g4509 = NOT(I7906)
--	g6440 = NOT(g6150)
--	g1976 = NOT(g643)
--	g11205 = NOT(g11112)
--	I6477 = NOT(g2069)
--	I9632 = NOT(g5557)
--	g7952 = NOT(g7427)
--	I15311 = NOT(g10013)
--	g9450 = NOT(g9097)
--	g5305 = NOT(g4378)
--	g5801 = NOT(g5320)
--	I5734 = NOT(g2097)
--	I6523 = NOT(g2819)
--	g2155 = NOT(I5070)
--	I4820 = NOT(g865)
--	I17243 = NOT(g11396)
--	g2355 = NOT(I5435)
--	g2851 = NOT(I5979)
--	I7249 = NOT(g2833)
--	I12559 = NOT(g7477)
--	I14315 = NOT(g8815)
--	I6643 = NOT(g3008)
--	g8213 = NOT(g7826)
--	I10819 = NOT(g6706)
--	g11311 = NOT(I17100)
--	I10910 = NOT(g6703)
--	I12424 = NOT(g7635)
--	I9102 = NOT(g5586)
--	I9208 = NOT(g5047)
--	g3707 = NOT(g2920)
--	I9302 = NOT(g5576)
--	I14910 = NOT(g9532)
--	g7616 = NOT(I12196)
--	g7561 = NOT(I12015)
--	g4067 = NOT(I7194)
--	g3759 = NOT(I6958)
--	I8278 = NOT(g4495)
--	I14257 = NOT(g8805)
--	g5748 = NOT(I9320)
--	I10979 = NOT(g6565)
--	g2964 = NOT(I6193)
--	g4418 = NOT(I7760)
--	I9869 = NOT(g5405)
--	g4467 = NOT(g3829)
--	I15072 = NOT(g9713)
--	I14979 = NOT(g9671)
--	g4290 = NOT(g3586)
--	I10111 = NOT(g5754)
--	I14055 = NOT(g8650)
--	g10871 = NOT(I16583)
--	g11051 = NOT(I16814)
--	I5992 = NOT(g2195)
--	g7004 = NOT(I11143)
--	I16583 = NOT(g10848)
--	g11072 = NOT(g10913)
--	I17773 = NOT(g11650)
--	I15592 = NOT(g10163)
--	I15756 = NOT(g10266)
--	g7527 = NOT(g7148)
--	I17268 = NOT(g11351)
--	I6742 = NOT(g3326)
--	I12544 = NOT(g7669)
--	g4093 = NOT(g2965)
--	I8282 = NOT(g4770)
--	g6151 = NOT(I9872)
--	g7764 = NOT(I12457)
--	g4256 = NOT(g3664)
--	g6648 = NOT(I10607)
--	g9777 = NOT(g9474)
--	g7546 = NOT(I11970)
--	I5080 = NOT(g36)
--	I15350 = NOT(g10001)
--	I10384 = NOT(g5842)
--	g10162 = NOT(I15482)
--	g3715 = NOT(g2920)
--	I9265 = NOT(g5085)
--	I16787 = NOT(g10896)
--	g11350 = NOT(g11287)
--	I5713 = NOT(g2436)
--	I15820 = NOT(g10204)
--	g5091 = NOT(g4385)
--	g8056 = NOT(g7671)
--	I13317 = NOT(g8093)
--	I12610 = NOT(g7627)
--	g4181 = NOT(I7360)
--	I6754 = NOT(g2906)
--	g8529 = NOT(I13738)
--	I14094 = NOT(g8700)
--	g4381 = NOT(g3914)
--	g7925 = NOT(g7476)
--	I9786 = NOT(g5396)
--	g2118 = NOT(g1854)
--	g8348 = NOT(I13424)
--	I12255 = NOT(g7203)
--	I6273 = NOT(g2482)
--	g2872 = NOT(I6016)
--	I16105 = NOT(g10382)
--	g10629 = NOT(g10583)
--	I10150 = NOT(g5705)
--	g5169 = NOT(g4596)
--	g4197 = NOT(I7408)
--	I10801 = NOT(g6536)
--	g8155 = NOT(I13048)
--	g11396 = NOT(I17231)
--	I13002 = NOT(g8045)
--	g8355 = NOT(I13445)
--	g10220 = NOT(I15592)
--	g5007 = NOT(I8379)
--	I13057 = NOT(g7843)
--	g2652 = NOT(g2008)
--	g2057 = NOT(g754)
--	g10628 = NOT(I16307)
--	I12678 = NOT(g7376)
--	I13128 = NOT(g7976)
--	g2843 = NOT(I5963)
--	g10911 = NOT(I16685)
--	g7320 = NOT(I11608)
--	g2989 = NOT(g2135)
--	g3539 = NOT(g3015)
--	g4263 = NOT(g3586)
--	I13245 = NOT(g8269)
--	I11626 = NOT(g7042)
--	I16769 = NOT(g10894)
--	g5718 = NOT(I9256)
--	I12460 = NOT(g7569)
--	I12939 = NOT(g7977)
--	g5767 = NOT(I9349)
--	I15691 = NOT(g10233)
--	I9296 = NOT(g4908)
--	I10018 = NOT(g5862)
--	I11299 = NOT(g6727)
--	I13323 = NOT(g8203)
--	I7176 = NOT(g2623)
--	I5976 = NOT(g2186)
--	g2549 = NOT(g1386)
--	I6572 = NOT(g2853)
--	I10526 = NOT(g6161)
--	g8063 = NOT(I12907)
--	g2834 = NOT(I5952)
--	g2971 = NOT(g2046)
--	g6172 = NOT(I9901)
--	g6278 = NOT(I10093)
--	g7617 = NOT(I12199)
--	I7405 = NOT(g3861)
--	g7906 = NOT(I12694)
--	g7789 = NOT(I12532)
--	g11405 = NOT(I17258)
--	g5261 = NOT(g4640)
--	g10591 = NOT(I16258)
--	I6543 = NOT(g3186)
--	g3362 = NOT(I6546)
--	g3419 = NOT(g3104)
--	I7829 = NOT(g3425)
--	g6667 = NOT(I10630)
--	g7516 = NOT(g7148)
--	g4562 = NOT(I7973)
--	g6343 = NOT(I10248)
--	g10754 = NOT(I16439)
--	g9353 = NOT(I14564)
--	g3052 = NOT(I6264)
--	g10355 = NOT(I15829)
--	g5415 = NOT(I8848)
--	g6282 = NOT(I10105)
--	g7771 = NOT(I12478)
--	g6566 = NOT(g5791)
--	I11737 = NOT(g7027)
--	g8279 = NOT(I13209)
--	g2121 = NOT(I5041)
--	g4631 = NOT(g3820)
--	I12875 = NOT(g7638)
--	g10825 = NOT(I16537)
--	I10917 = NOT(g6732)
--	I15583 = NOT(g10157)
--	g9802 = NOT(g9490)
--	g1999 = NOT(g806)
--	I11232 = NOT(g6537)
--	g4257 = NOT(g3664)
--	g6134 = NOT(I9839)
--	g5664 = NOT(I9153)
--	g8318 = NOT(I13338)
--	g8872 = NOT(I14188)
--	I9706 = NOT(g5221)
--	g2232 = NOT(I5221)
--	g10172 = NOT(I15510)
--	g11046 = NOT(I16799)
--	g3086 = NOT(g2276)
--	g5203 = NOT(g4640)
--	g2253 = NOT(g100)
--	g3728 = NOT(I6904)
--	g2813 = NOT(I5913)
--	I9029 = NOT(g4781)
--	g8989 = NOT(I14388)
--	I14077 = NOT(g8758)
--	I9171 = NOT(g4902)
--	g6555 = NOT(g5740)
--	I10706 = NOT(g6080)
--	I9371 = NOT(g5075)
--	g6804 = NOT(I10822)
--	I15787 = NOT(g10269)
--	I6414 = NOT(g2342)
--	g3730 = NOT(g3015)
--	g2909 = NOT(I6080)
--	I9956 = NOT(g5485)
--	I10689 = NOT(g6059)
--	g3385 = NOT(g3121)
--	I5383 = NOT(g886)
--	I15302 = NOT(g10007)
--	g11357 = NOT(I17182)
--	g7991 = NOT(I12809)
--	I6513 = NOT(g2812)
--	g2606 = NOT(I5719)
--	g10319 = NOT(g10270)
--	g4441 = NOT(g3914)
--	g6113 = NOT(I9792)
--	g6313 = NOT(I10198)
--	g7078 = NOT(I11309)
--	g7340 = NOT(I11668)
--	I10102 = NOT(g5730)
--	I16778 = NOT(g10891)
--	I13831 = NOT(g8560)
--	g10318 = NOT(I15752)
--	I8050 = NOT(g4089)
--	I13445 = NOT(g8149)
--	I5588 = NOT(g1203)
--	g8121 = NOT(I12978)
--	g10227 = NOT(I15601)
--	g7907 = NOT(g7664)
--	I6436 = NOT(g2351)
--	I6679 = NOT(g2902)
--	g8321 = NOT(I13347)
--	g4673 = NOT(g4013)
--	g6202 = NOT(g5426)
--	g8670 = NOT(g8551)
--	g5689 = NOT(I9216)
--	I8996 = NOT(g4757)
--	I9684 = NOT(g5426)
--	g7035 = NOT(I11194)
--	I15768 = NOT(g10249)
--	I9138 = NOT(g5210)
--	I9639 = NOT(g5126)
--	g7959 = NOT(I12751)
--	I10066 = NOT(g5778)
--	I9338 = NOT(g5576)
--	I10231 = NOT(g6111)
--	g8625 = NOT(g8487)
--	g7082 = NOT(I11315)
--	g2586 = NOT(g1972)
--	g5216 = NOT(g4445)
--	g10540 = NOT(I16187)
--	I17410 = NOT(g11419)
--	g6094 = NOT(I9749)
--	I11498 = NOT(g6578)
--	I12595 = NOT(g7706)
--	I16647 = NOT(g10866)
--	g10058 = NOT(I15281)
--	I16356 = NOT(g10597)
--	g4669 = NOT(g4013)
--	I8724 = NOT(g4791)
--	g6567 = NOT(I10495)
--	g5671 = NOT(I9174)
--	g4368 = NOT(I7665)
--	I11989 = NOT(g6919)
--	I17666 = NOT(g11603)
--	I10885 = NOT(g6332)
--	I8379 = NOT(g4231)
--	g3331 = NOT(I6510)
--	g10203 = NOT(g10177)
--	I14876 = NOT(g9526)
--	I11611 = NOT(g6913)
--	g7656 = NOT(I12265)
--	g4772 = NOT(g3440)
--	g3406 = NOT(I6611)
--	I11722 = NOT(g7034)
--	I7399 = NOT(g4113)
--	g10044 = NOT(I15263)
--	g3635 = NOT(I6812)
--	I6022 = NOT(g2258)
--	g4458 = NOT(I7817)
--	g2570 = NOT(g207)
--	g2860 = NOT(I5998)
--	g2341 = NOT(I5403)
--	g9262 = NOT(I14473)
--	g3682 = NOT(g2920)
--	g6593 = NOT(I10557)
--	I9759 = NOT(g5344)
--	g8519 = NOT(I13726)
--	g3105 = NOT(g2482)
--	g7915 = NOT(g7473)
--	g3305 = NOT(I6474)
--	g10281 = NOT(g10162)
--	g98 = NOT(I4783)
--	g2645 = NOT(g1991)
--	I8835 = NOT(g4791)
--	g5826 = NOT(I9440)
--	I12418 = NOT(g7568)
--	I12822 = NOT(g7677)
--	g10902 = NOT(I16660)
--	g10377 = NOT(I15855)
--	g8606 = NOT(g8481)
--	g7214 = NOT(I11450)
--	I6947 = NOT(g2860)
--	g10120 = NOT(I15368)
--	g4011 = NOT(I7151)
--	g9076 = NOT(g8892)
--	g5741 = NOT(I9305)
--	g3748 = NOT(g2971)
--	g4411 = NOT(I7743)
--	g4734 = NOT(g3586)
--	I11342 = NOT(g6686)
--	g9889 = NOT(I15072)
--	g7110 = NOT(I11345)
--	g6264 = NOT(I10051)
--	g7310 = NOT(I11578)
--	I6560 = NOT(g2845)
--	I7291 = NOT(g3212)
--	I8611 = NOT(g4562)
--	I10456 = NOT(g5844)
--	I15482 = NOT(g10115)
--	g5638 = NOT(I9077)
--	g3226 = NOT(I6403)
--	g6933 = NOT(I11061)
--	g7663 = NOT(I12282)
--	I11650 = NOT(g6938)
--	g10699 = NOT(I16376)
--	g2607 = NOT(I5722)
--	I12853 = NOT(g7638)
--	I16897 = NOT(g10947)
--	I5240 = NOT(g64)
--	g2962 = NOT(I6183)
--	g6521 = NOT(I10437)
--	I17084 = NOT(g11249)
--	g4474 = NOT(g3820)
--	g10290 = NOT(I15694)
--	g2158 = NOT(I5077)
--	g6050 = NOT(I9677)
--	g6641 = NOT(I10598)
--	I11198 = NOT(g6521)
--	I9498 = NOT(g5081)
--	I12589 = NOT(g7571)
--	g10698 = NOT(I16373)
--	g2506 = NOT(g636)
--	g6450 = NOT(I10378)
--	I6037 = NOT(g2560)
--	I17321 = NOT(g11348)
--	g5883 = NOT(g5309)
--	I10314 = NOT(g6251)
--	g7402 = NOT(g6860)
--	I6495 = NOT(g2076)
--	I9833 = NOT(g5197)
--	I17179 = NOT(g11307)
--	I11528 = NOT(g6796)
--	I6102 = NOT(g2240)
--	I16717 = NOT(g10779)
--	I17531 = NOT(g11488)
--	I7694 = NOT(g3742)
--	I11330 = NOT(g6571)
--	I6302 = NOT(g2243)
--	g3373 = NOT(I6565)
--	I15778 = NOT(g10255)
--	g7762 = NOT(I12451)
--	g3491 = NOT(g2669)
--	g4080 = NOT(g2903)
--	I5116 = NOT(g40)
--	g11081 = NOT(I16856)
--	I7852 = NOT(g3438)
--	I7923 = NOT(g3394)
--	g5758 = NOT(I9338)
--	g8141 = NOT(I13020)
--	g8570 = NOT(I13803)
--	g5066 = NOT(I8436)
--	g5589 = NOT(I9001)
--	g6724 = NOT(I10719)
--	g8341 = NOT(I13403)
--	I10054 = NOT(g5728)
--	g2275 = NOT(g757)
--	I9539 = NOT(g5354)
--	I9896 = NOT(g5295)
--	g4713 = NOT(g3546)
--	I10243 = NOT(g5918)
--	I11132 = NOT(g6451)
--	I11869 = NOT(g6894)
--	g7877 = NOT(g7479)
--	I7701 = NOT(g3513)
--	g3369 = NOT(I6557)
--	I5565 = NOT(g1713)
--	g3007 = NOT(I6240)
--	g9339 = NOT(I14522)
--	I15356 = NOT(g10013)
--	g7657 = NOT(I12268)
--	g6878 = NOT(I10966)
--	I15826 = NOT(g10205)
--	I6917 = NOT(g2832)
--	I15380 = NOT(g10098)
--	I4894 = NOT(g258)
--	g2174 = NOT(g31)
--	g3459 = NOT(I6661)
--	g6289 = NOT(I10126)
--	g9024 = NOT(I14409)
--	g2374 = NOT(g591)
--	I12616 = NOT(g7534)
--	I9162 = NOT(g5035)
--	g7556 = NOT(I11992)
--	I9268 = NOT(g5305)
--	I16723 = NOT(g10851)
--	g3767 = NOT(I6976)
--	g10547 = NOT(I16206)
--	g9424 = NOT(g9076)
--	g10895 = NOT(I16647)
--	I7886 = NOT(g4076)
--	I9362 = NOT(g5013)
--	g6835 = NOT(I10885)
--	g2985 = NOT(I6217)
--	g9809 = NOT(I14944)
--	g5827 = NOT(I9443)
--	g6882 = NOT(I10974)
--	g7928 = NOT(g7508)
--	I10156 = NOT(g6100)
--	I10655 = NOT(g6036)
--	I15672 = NOT(g10132)
--	g3582 = NOT(g3164)
--	I16387 = NOT(g10629)
--	I17334 = NOT(g11360)
--	g6271 = NOT(I10072)
--	I11225 = NOT(g6534)
--	g10226 = NOT(I15598)
--	I9452 = NOT(g5085)
--	g11182 = NOT(I16947)
--	g11651 = NOT(I17755)
--	g7064 = NOT(I11269)
--	I5210 = NOT(g58)
--	g2239 = NOT(I5240)
--	I10180 = NOT(g6107)
--	g9672 = NOT(I14805)
--	I13708 = NOT(g8337)
--	g5774 = NOT(I9362)
--	g7899 = NOT(I12683)
--	g3793 = NOT(g2593)
--	g7464 = NOT(I11858)
--	I12053 = NOT(g6928)
--	g8358 = NOT(I13454)
--	I12809 = NOT(g7686)
--	g7785 = NOT(I12520)
--	I16811 = NOT(g10908)
--	g10551 = NOT(I16214)
--	I6233 = NOT(g2299)
--	g2832 = NOT(I5946)
--	I12466 = NOT(g7585)
--	g3415 = NOT(g3121)
--	g3227 = NOT(I6406)
--	I7825 = NOT(g3414)
--	g6799 = NOT(I10807)
--	g2853 = NOT(g2171)
--	I11043 = NOT(g6412)
--	I6454 = NOT(g2368)
--	I13043 = NOT(g8055)
--	I17216 = NOT(g11291)
--	g2420 = NOT(g237)
--	g6674 = NOT(I10639)
--	I9486 = NOT(g5066)
--	g11513 = NOT(I17558)
--	I12177 = NOT(g7259)
--	g10127 = NOT(I15383)
--	g3664 = NOT(g3209)
--	g8275 = NOT(I13197)
--	g2507 = NOT(I5584)
--	g8311 = NOT(I13317)
--	g3246 = NOT(g2482)
--	I15448 = NOT(g10056)
--	g5509 = NOT(g4739)
--	g4326 = NOT(g3863)
--	I14694 = NOT(g9259)
--	I7408 = NOT(g4125)
--	g7237 = NOT(I11477)
--	g10490 = NOT(I16105)
--	I9185 = NOT(g4915)
--	I7336 = NOT(g3997)
--	g3721 = NOT(I6891)
--	g11505 = NOT(I17534)
--	I11602 = NOT(g6833)
--	I11810 = NOT(g7246)
--	g11404 = NOT(I17255)
--	g6132 = NOT(I9833)
--	g5662 = NOT(I9147)
--	I6553 = NOT(g3186)
--	I4850 = NOT(g1958)
--	g7844 = NOT(I12631)
--	I17543 = NOT(g11499)
--	I11068 = NOT(g6426)
--	I13068 = NOT(g7906)
--	g6680 = NOT(I10643)
--	g6209 = NOT(I9956)
--	g8985 = NOT(I14376)
--	I11879 = NOT(g6893)
--	g5994 = NOT(I9612)
--	g10889 = NOT(I16629)
--	I16850 = NOT(g10905)
--	I11970 = NOT(g6918)
--	g7394 = NOT(I11778)
--	I10557 = NOT(g6197)
--	g10354 = NOT(I15826)
--	g2905 = NOT(I6068)
--	g7089 = NOT(I11322)
--	g7731 = NOT(I12376)
--	g10888 = NOT(I16626)
--	g6802 = NOT(I10816)
--	g8239 = NOT(g7826)
--	g4183 = NOT(I7366)
--	g9273 = NOT(I14490)
--	g4608 = NOT(g3829)
--	g5816 = NOT(I9424)
--	I5922 = NOT(g2170)
--	I7465 = NOT(g3726)
--	g7966 = NOT(I12762)
--	g2100 = NOT(I4948)
--	I10278 = NOT(g5815)
--	g3940 = NOT(g2920)
--	g6558 = NOT(I10484)
--	I12009 = NOT(g6915)
--	I6888 = NOT(g2960)
--	I8262 = NOT(g4636)
--	I11967 = NOT(g6911)
--	g8020 = NOT(I12862)
--	I10286 = NOT(g6237)
--	g8420 = NOT(I13574)
--	I5060 = NOT(g1191)
--	g10931 = NOT(g10827)
--	g3388 = NOT(I6590)
--	I10039 = NOT(g5718)
--	I14306 = NOT(g8812)
--	I11459 = NOT(g6488)
--	g11433 = NOT(I17350)
--	g9572 = NOT(I14709)
--	g5685 = NOT(I9208)
--	g5197 = NOT(I8611)
--	g5700 = NOT(I9237)
--	g8794 = NOT(I14109)
--	g5397 = NOT(I8835)
--	g2750 = NOT(I5818)
--	I8889 = NOT(g4553)
--	g11620 = NOT(I17678)
--	g10190 = NOT(I15548)
--	I8476 = NOT(g4577)
--	g4361 = NOT(I7648)
--	I9766 = NOT(g5348)
--	I15811 = NOT(g10200)
--	g3428 = NOT(I6639)
--	I7096 = NOT(g3186)
--	I12454 = NOT(g7544)
--	I9087 = NOT(g5113)
--	I9105 = NOT(g5589)
--	I9305 = NOT(g4970)
--	I9801 = NOT(g5416)
--	g3430 = NOT(I6643)
--	g7814 = NOT(I12607)
--	I12712 = NOT(g7441)
--	g11646 = NOT(I17742)
--	g4051 = NOT(I7166)
--	I10601 = NOT(g5996)
--	I13010 = NOT(g8047)
--	g11343 = NOT(I17152)
--	I13918 = NOT(g8451)
--	I16379 = NOT(g10598)
--	g4127 = NOT(I7276)
--	g4451 = NOT(g3638)
--	I15971 = NOT(g10408)
--	g4327 = NOT(I7600)
--	I17265 = NOT(g11352)
--	g7350 = NOT(I11698)
--	g2040 = NOT(g1786)
--	g6574 = NOT(I10514)
--	I12907 = NOT(g7959)
--	I5995 = NOT(g2196)
--	I11079 = NOT(g6649)
--	g10546 = NOT(I16203)
--	g7038 = NOT(I11201)
--	I11444 = NOT(g6653)
--	I17416 = NOT(g11420)
--	g10211 = NOT(I15583)
--	g9534 = NOT(I14687)
--	g9961 = NOT(I15162)
--	g6714 = NOT(g5867)
--	g7438 = NOT(g7232)
--	g7773 = NOT(I12484)
--	I11599 = NOT(g6832)
--	g7009 = NOT(I11152)
--	g11369 = NOT(I17194)
--	g2123 = NOT(I5047)
--	I6639 = NOT(g2632)
--	g4346 = NOT(I7625)
--	g8515 = NOT(I13714)
--	g10088 = NOT(I15317)
--	I8285 = NOT(g4771)
--	I10937 = NOT(g6552)
--	I12239 = NOT(g7073)
--	I5840 = NOT(g2432)
--	I15368 = NOT(g9990)
--	I17510 = NOT(g11481)
--	I16742 = NOT(g10857)
--	g8100 = NOT(g7947)
--	I16944 = NOT(g11079)
--	g3910 = NOT(g3015)
--	I13086 = NOT(g7924)
--	g7769 = NOT(I12472)
--	I15412 = NOT(g10075)
--	g3638 = NOT(I6821)
--	I8139 = NOT(g3681)
--	g7212 = NOT(I11444)
--	g5723 = NOT(I9265)
--	I14884 = NOT(g9454)
--	g11412 = NOT(I17277)
--	I11817 = NOT(g7246)
--	I10168 = NOT(g5982)
--	g5101 = NOT(I8473)
--	g5817 = NOT(I9427)
--	I11322 = NOT(g6652)
--	g7918 = NOT(g7505)
--	g5301 = NOT(g4373)
--	g7967 = NOT(I12765)
--	g6262 = NOT(I10045)
--	I15229 = NOT(g9968)
--	g2351 = NOT(I5427)
--	I11159 = NOT(g6478)
--	g10700 = NOT(I16379)
--	g2648 = NOT(I5765)
--	I9491 = NOT(g5072)
--	g10126 = NOT(I15380)
--	I8024 = NOT(g4117)
--	I11901 = NOT(g6897)
--	I16802 = NOT(g10902)
--	g2530 = NOT(I5641)
--	g6736 = NOT(I10739)
--	I13125 = NOT(g7975)
--	g8750 = NOT(I14045)
--	I10666 = NOT(g6042)
--	g4508 = NOT(g3946)
--	g10250 = NOT(g10136)
--	g2655 = NOT(g2013)
--	g4944 = NOT(g4430)
--	g4240 = NOT(g3664)
--	I11783 = NOT(g7246)
--	I16793 = NOT(g11014)
--	I7342 = NOT(g4011)
--	I9602 = NOT(g5013)
--	g4472 = NOT(I7847)
--	I10015 = NOT(g5641)
--	I5704 = NOT(g2056)
--	g7993 = NOT(I12813)
--	I7255 = NOT(g3227)
--	g6076 = NOT(I9717)
--	I4906 = NOT(g119)
--	I11656 = NOT(g7122)
--	I6049 = NOT(g2219)
--	g5751 = NOT(I9323)
--	g3758 = NOT(I6955)
--	g3066 = NOT(g2135)
--	I8231 = NOT(g4170)
--	g4443 = NOT(g3359)
--	g10296 = NOT(I15708)
--	g8440 = NOT(I13618)
--	I11680 = NOT(g7064)
--	g8969 = NOT(I14340)
--	I17116 = NOT(g11229)
--	g2410 = NOT(g1453)
--	g9679 = NOT(g9452)
--	I7726 = NOT(g3378)
--	g6175 = NOT(g5320)
--	g4116 = NOT(I7260)
--	I7154 = NOT(g2617)
--	g8323 = NOT(I13351)
--	g6871 = NOT(g6724)
--	g2884 = NOT(I6040)
--	I7354 = NOT(g4066)
--	g2839 = NOT(I5957)
--	g3365 = NOT(I6553)
--	g3861 = NOT(I7054)
--	I6498 = NOT(g2958)
--	I17746 = NOT(g11643)
--	g3055 = NOT(g2135)
--	I5053 = NOT(g1188)
--	I15959 = NOT(g10402)
--	g6285 = NOT(I10114)
--	g11627 = NOT(I17695)
--	g7921 = NOT(g7463)
--	g10197 = NOT(I15565)
--	g5673 = NOT(I9180)
--	g4347 = NOT(g3880)
--	I8551 = NOT(g4342)
--	I10084 = NOT(g5742)
--	g2172 = NOT(g43)
--	g3333 = NOT(g2779)
--	I9415 = NOT(g5047)
--	g11112 = NOT(I16897)
--	I17237 = NOT(g11394)
--	g4681 = NOT(g3546)
--	g10870 = NOT(I16580)
--	g11050 = NOT(I16811)
--	I8499 = NOT(g4330)
--	I12577 = NOT(g7532)
--	g8151 = NOT(g8036)
--	g10527 = NOT(g10462)
--	g3774 = NOT(I6999)
--	g8351 = NOT(I13433)
--	I17340 = NOT(g11366)
--	g4533 = NOT(I7938)
--	I13017 = NOT(g7848)
--	I13364 = NOT(g8221)
--	I15386 = NOT(g10101)
--	g6184 = NOT(I9915)
--	g2235 = NOT(g96)
--	g2343 = NOT(g1927)
--	I12439 = NOT(g7663)
--	g5669 = NOT(I9168)
--	I10531 = NOT(g6169)
--	I17684 = NOT(g11609)
--	g6339 = NOT(I10240)
--	I14179 = NOT(g8785)
--	g4210 = NOT(I7447)
--	I14531 = NOT(g9273)
--	I7112 = NOT(g3186)
--	I17142 = NOT(g11301)
--	g11096 = NOT(I16879)
--	g7620 = NOT(I12208)
--	g4596 = NOT(I8007)
--	g3538 = NOT(I6726)
--	I6019 = NOT(g2554)
--	g4013 = NOT(I7157)
--	g6424 = NOT(g6140)
--	I16626 = NOT(g10859)
--	I10186 = NOT(g6110)
--	g6737 = NOT(g6016)
--	g10867 = NOT(I16571)
--	g2334 = NOT(I5388)
--	g10894 = NOT(I16644)
--	g6809 = NOT(I10837)
--	I10685 = NOT(g6054)
--	g5743 = NOT(I9311)
--	g4413 = NOT(I7749)
--	g5890 = NOT(g5361)
--	I11289 = NOT(g6508)
--	I6052 = NOT(g2220)
--	g2548 = NOT(I5667)
--	I14373 = NOT(g8956)
--	I11309 = NOT(g6531)
--	I5929 = NOT(g2225)
--	I13023 = NOT(g8050)
--	g8884 = NOT(I14224)
--	I16298 = NOT(g10553)
--	I13224 = NOT(g8261)
--	g7788 = NOT(I12529)
--	g6077 = NOT(I9720)
--	g11429 = NOT(I17340)
--	g5011 = NOT(I8385)
--	I16775 = NOT(g10889)
--	g3067 = NOT(I6273)
--	I13571 = NOT(g8355)
--	g10315 = NOT(g10243)
--	g5856 = NOT(g5245)
--	g5734 = NOT(I9290)
--	g10819 = NOT(I16525)
--	g11428 = NOT(I17337)
--	g10910 = NOT(I16682)
--	g3290 = NOT(I6461)
--	I17362 = NOT(g11376)
--	g10202 = NOT(g10171)
--	I10334 = NOT(g6003)
--	g10257 = NOT(g10197)
--	g4317 = NOT(I7586)
--	g8278 = NOT(I13206)
--	I4876 = NOT(g580)
--	g3093 = NOT(I6299)
--	g1998 = NOT(g802)
--	g5474 = NOT(I8889)
--	g10111 = NOT(I15347)
--	g7192 = NOT(g6742)
--	g5992 = NOT(I9608)
--	g7085 = NOT(I11318)
--	g3256 = NOT(I6424)
--	I7746 = NOT(g3763)
--	g6634 = NOT(I10589)
--	I9188 = NOT(g4908)
--	I10762 = NOT(g6127)
--	g8667 = NOT(I13952)
--	g3816 = NOT(g3228)
--	g8143 = NOT(g8029)
--	I13816 = NOT(g8559)
--	I15548 = NOT(g10083)
--	I6504 = NOT(g3214)
--	I9388 = NOT(g5576)
--	g8235 = NOT(g7967)
--	g8343 = NOT(I13409)
--	g6742 = NOT(g5830)
--	g11548 = NOT(g11519)
--	g6104 = NOT(I9769)
--	I14964 = NOT(g9762)
--	g10590 = NOT(I16255)
--	I9216 = NOT(g4935)
--	I6385 = NOT(g2260)
--	g6304 = NOT(I10171)
--	I16856 = NOT(g10909)
--	g8566 = NOT(I13791)
--	g6499 = NOT(g5867)
--	I16261 = NOT(g10556)
--	g2202 = NOT(g148)
--	g11504 = NOT(I17531)
--	g8988 = NOT(I14385)
--	g4775 = NOT(I8139)
--	I11752 = NOT(g7032)
--	g8134 = NOT(I13005)
--	g7941 = NOT(g7406)
--	I15317 = NOT(g10025)
--	I6025 = NOT(g2259)
--	g2908 = NOT(I6077)
--	g8334 = NOT(I13382)
--	g9265 = NOT(g8892)
--	g6926 = NOT(I11046)
--	g2094 = NOT(I4924)
--	I12415 = NOT(g7631)
--	g11317 = NOT(I17112)
--	g10094 = NOT(I15329)
--	g3397 = NOT(g2896)
--	g8548 = NOT(g8390)
--	g2518 = NOT(g590)
--	g4060 = NOT(g3144)
--	g4460 = NOT(g3820)
--	I9564 = NOT(g5109)
--	I7468 = NOT(g3697)
--	g6273 = NOT(I10078)
--	I8885 = NOT(g4548)
--	g8804 = NOT(I14133)
--	I14543 = NOT(g9311)
--	I8414 = NOT(g4293)
--	g10150 = NOT(I15448)
--	g10801 = NOT(I16507)
--	I9826 = NOT(g5390)
--	I10117 = NOT(g6241)
--	g7708 = NOT(I12339)
--	I13669 = NOT(g8294)
--	g10735 = NOT(I16416)
--	g10877 = NOT(I16601)
--	g11057 = NOT(g10937)
--	g7520 = NOT(I11898)
--	g8792 = NOT(I14105)
--	I17347 = NOT(g11373)
--	I7677 = NOT(g3735)
--	I11668 = NOT(g7043)
--	g6044 = NOT(I9665)
--	g2593 = NOT(g1973)
--	g7031 = NOT(g6413)
--	g4739 = NOT(g4117)
--	I8903 = NOT(g4561)
--	g6444 = NOT(g6158)
--	g11245 = NOT(g11112)
--	g7431 = NOT(I11821)
--	I15323 = NOT(g10019)
--	g6269 = NOT(I10066)
--	I15299 = NOT(g9995)
--	g7812 = NOT(I12601)
--	g11626 = NOT(I17692)
--	g9770 = NOT(g9432)
--	g10196 = NOT(I15562)
--	I11489 = NOT(g6569)
--	g10695 = NOT(I16366)
--	g5688 = NOT(I9213)
--	g11323 = NOT(I17124)
--	I13489 = NOT(g8233)
--	g2965 = NOT(I6196)
--	I6406 = NOT(g2339)
--	I5475 = NOT(g1289)
--	I7716 = NOT(g3751)
--	g6572 = NOT(g5805)
--	g6862 = NOT(g6720)
--	g7376 = NOT(I11756)
--	I5949 = NOT(g2540)
--	g10526 = NOT(g10460)
--	g8313 = NOT(I13323)
--	I12484 = NOT(g7580)
--	I14242 = NOT(g8787)
--	I9108 = NOT(g5593)
--	I15775 = NOT(g10253)
--	I13424 = NOT(g8200)
--	g4479 = NOT(I7858)
--	g9532 = NOT(I14681)
--	I9308 = NOT(g5494)
--	g6712 = NOT(g5984)
--	I8036 = NOT(g3820)
--	g4294 = NOT(g3664)
--	I10123 = NOT(g5676)
--	g6543 = NOT(g5888)
--	g4840 = NOT(I8199)
--	I8436 = NOT(g4462)
--	g9553 = NOT(I14694)
--	I5292 = NOT(g76)
--	I9883 = NOT(g5557)
--	I14123 = NOT(g8767)
--	g3723 = NOT(g3071)
--	g7765 = NOT(I12460)
--	g7286 = NOT(I11534)
--	g4190 = NOT(I7387)
--	I5998 = NOT(g2197)
--	g4390 = NOT(g3914)
--	I10807 = NOT(g6396)
--	g10457 = NOT(I15962)
--	g3817 = NOT(I7043)
--	g7911 = NOT(g7664)
--	I5646 = NOT(g940)
--	I10974 = NOT(g6563)
--	g8094 = NOT(g7987)
--	g2050 = NOT(g1861)
--	g2641 = NOT(g1987)
--	I8831 = NOT(g4480)
--	I15232 = NOT(g9974)
--	I10639 = NOT(g5830)
--	I17516 = NOT(g11483)
--	g2450 = NOT(g1351)
--	I16432 = NOT(g10702)
--	g4501 = NOT(g3946)
--	g8518 = NOT(I13723)
--	g6729 = NOT(I10724)
--	g6961 = NOT(I11115)
--	g8567 = NOT(I13794)
--	I10293 = NOT(g5863)
--	g4156 = NOT(I7295)
--	I11713 = NOT(g7023)
--	g7733 = NOT(I12380)
--	I5850 = NOT(g2273)
--	g7270 = NOT(I11515)
--	g9990 = NOT(I15190)
--	g6927 = NOT(I11049)
--	g3751 = NOT(I6944)
--	I9165 = NOT(g5037)
--	I16461 = NOT(g10735)
--	I9571 = NOT(g5509)
--	I9365 = NOT(g5392)
--	g7610 = NOT(I12180)
--	g2179 = NOT(g89)
--	g4942 = NOT(I8308)
--	g9029 = NOT(I14424)
--	g6014 = NOT(g5309)
--	g7073 = NOT(I11296)
--	I12799 = NOT(g7556)
--	g7796 = NOT(I12553)
--	I12813 = NOT(g7688)
--	g6885 = NOT(I10979)
--	g9429 = NOT(g9082)
--	g22 = NOT(I4777)
--	g7473 = NOT(g7148)
--	I10391 = NOT(g5838)
--	I17209 = NOT(g11289)
--	g6660 = NOT(I10623)
--	I11255 = NOT(g6547)
--	g10256 = NOT(g10140)
--	I6173 = NOT(g2125)
--	g11512 = NOT(I17555)
--	I13255 = NOT(g8270)
--	I14391 = NOT(g8928)
--	I16650 = NOT(g10776)
--	I6373 = NOT(g2024)
--	I6091 = NOT(g2270)
--	g5183 = NOT(g4640)
--	g7124 = NOT(I11363)
--	g7980 = NOT(I12786)
--	g7324 = NOT(I11620)
--	g10280 = NOT(g10160)
--	g6903 = NOT(I11005)
--	g2777 = NOT(g2276)
--	I5919 = NOT(g2530)
--	I11188 = NOT(g6513)
--	g7069 = NOT(I11286)
--	I12805 = NOT(g7684)
--	I13188 = NOT(g8171)
--	g5779 = NOT(I9371)
--	I13678 = NOT(g8306)
--	I14579 = NOT(g9272)
--	g4954 = NOT(g4509)
--	g4250 = NOT(g3698)
--	g4163 = NOT(I7308)
--	I5952 = NOT(g2506)
--	g2882 = NOT(I6034)
--	g7540 = NOT(I11956)
--	g8160 = NOT(I13057)
--	g4363 = NOT(I7654)
--	I11686 = NOT(g7039)
--	I16528 = NOT(g10732)
--	I7577 = NOT(g4124)
--	I5276 = NOT(g1411)
--	g8360 = NOT(I13460)
--	I16843 = NOT(g10898)
--	I6007 = NOT(g2199)
--	g5423 = NOT(g4300)
--	I13460 = NOT(g8155)
--	I17453 = NOT(g11451)
--	I11383 = NOT(g6385)
--	g2271 = NOT(g877)
--	g7377 = NOT(I11759)
--	g7206 = NOT(I11436)
--	g10157 = NOT(I15467)
--	g11445 = NOT(I17384)
--	g6036 = NOT(I9647)
--	I5561 = NOT(g869)
--	I13030 = NOT(g8052)
--	g2611 = NOT(I5734)
--	g4453 = NOT(I7810)
--	g8450 = NOT(I13648)
--	g6178 = NOT(g4977)
--	I6767 = NOT(g2914)
--	g11499 = NOT(I17516)
--	I8495 = NOT(g4325)
--	g3368 = NOT(g3138)
--	g9745 = NOT(g9454)
--	I11065 = NOT(g6750)
--	I6535 = NOT(g2826)
--	g1987 = NOT(g762)
--	g9338 = NOT(I14519)
--	g7287 = NOT(I11537)
--	g2799 = NOT(g2276)
--	g11498 = NOT(I17513)
--	I5986 = NOT(g2194)
--	g6135 = NOT(I9842)
--	g5665 = NOT(I9156)
--	g9109 = NOT(I14452)
--	g6335 = NOT(I10228)
--	I15989 = NOT(g10417)
--	g9309 = NOT(g8892)
--	g3531 = NOT(g2971)
--	I8869 = NOT(g4421)
--	g5127 = NOT(I8535)
--	g3458 = NOT(g3144)
--	g6182 = NOT(g5446)
--	g6288 = NOT(I10123)
--	I17274 = NOT(g11389)
--	g6382 = NOT(I10278)
--	I9662 = NOT(g5319)
--	g8179 = NOT(I13086)
--	g7849 = NOT(I12644)
--	g10876 = NOT(I16598)
--	g10885 = NOT(g10809)
--	g11056 = NOT(g10950)
--	g3743 = NOT(I6932)
--	g8379 = NOT(I13485)
--	g4912 = NOT(I8282)
--	I14116 = NOT(g8766)
--	g2997 = NOT(g2135)
--	g11611 = NOT(I17657)
--	I12400 = NOT(g7537)
--	g2541 = NOT(I5658)
--	g11080 = NOT(I16853)
--	I7426 = NOT(g3334)
--	I9290 = NOT(g5052)
--	g5146 = NOT(g4596)
--	g10854 = NOT(g10708)
--	g6805 = NOT(I10825)
--	g5633 = NOT(g4388)
--	g3505 = NOT(I6694)
--	g7781 = NOT(I12508)
--	I5970 = NOT(g2185)
--	g6749 = NOT(I10756)
--	I16708 = NOT(g10822)
--	g2238 = NOT(I5237)
--	g11432 = NOT(I17347)
--	I13837 = NOT(g8488)
--	g3411 = NOT(I6616)
--	I9093 = NOT(g5397)
--	g7900 = NOT(g7712)
--	I16258 = NOT(g10555)
--	I4948 = NOT(g586)
--	g2209 = NOT(g93)
--	g7797 = NOT(I12556)
--	I9256 = NOT(g5078)
--	I8265 = NOT(g4602)
--	I9816 = NOT(g5576)
--	g5696 = NOT(I9229)
--	I15461 = NOT(g10074)
--	g6947 = NOT(I11085)
--	I7984 = NOT(g3621)
--	I5224 = NOT(g61)
--	I7280 = NOT(g3208)
--	I10237 = NOT(g6120)
--	g6798 = NOT(I10804)
--	I8442 = NOT(g4464)
--	I12538 = NOT(g7658)
--	g8271 = NOT(I13185)
--	g2802 = NOT(g2276)
--	g11342 = NOT(I17149)
--	I10340 = NOT(g6205)
--	g1991 = NOT(g778)
--	I5120 = NOT(g622)
--	g3474 = NOT(I6679)
--	g9449 = NOT(g9094)
--	g6560 = NOT(g5759)
--	I14340 = NOT(g8820)
--	g5753 = NOT(I9329)
--	I8164 = NOT(g3566)
--	I15736 = NOT(g10258)
--	g10456 = NOT(I15959)
--	g5508 = NOT(I8929)
--	g11199 = NOT(g11112)
--	I14684 = NOT(g9124)
--	g11650 = NOT(I17752)
--	g7144 = NOT(I11387)
--	I11617 = NOT(g6839)
--	g7344 = NOT(I11680)
--	g5072 = NOT(I8442)
--	I7636 = NOT(g3330)
--	I13915 = NOT(g8451)
--	g5472 = NOT(I8885)
--	g8981 = NOT(I14364)
--	I9421 = NOT(g5063)
--	g8674 = NOT(I13959)
--	I5789 = NOT(g2162)
--	g5043 = NOT(g4840)
--	I11201 = NOT(g6522)
--	g10314 = NOT(I15744)
--	g7259 = NOT(I11494)
--	g5443 = NOT(I8872)
--	g6208 = NOT(I9953)
--	I7790 = NOT(g3782)
--	I16879 = NOT(g10936)
--	g6302 = NOT(I10165)
--	g10307 = NOT(I15729)
--	I15365 = NOT(g10025)
--	I7061 = NOT(g3050)
--	g6579 = NOT(g5949)
--	g5116 = NOT(g4682)
--	g6869 = NOT(I10949)
--	g7852 = NOT(g7479)
--	g7923 = NOT(g7527)
--	I17164 = NOT(g11320)
--	I7387 = NOT(g4083)
--	g10596 = NOT(I16269)
--	I11467 = NOT(g6488)
--	I11494 = NOT(g6574)
--	I13595 = NOT(g8339)
--	g8132 = NOT(I12999)
--	g6719 = NOT(I10710)
--	I12235 = NOT(g7082)
--	g8332 = NOT(I13376)
--	g10243 = NOT(I15635)
--	I11623 = NOT(g6841)
--	I12683 = NOT(g7387)
--	I6388 = NOT(g2329)
--	g8680 = NOT(I13965)
--	g10431 = NOT(g10328)
--	I11037 = NOT(g6629)
--	g8353 = NOT(I13439)
--	I14130 = NOT(g8769)
--	I10362 = NOT(g6224)
--	g2864 = NOT(g2298)
--	I10165 = NOT(g5948)
--	I13782 = NOT(g8515)
--	g6917 = NOT(I11029)
--	g4894 = NOT(I8247)
--	I6028 = NOT(g2208)
--	g10269 = NOT(g10154)
--	g8802 = NOT(I14127)
--	I6671 = NOT(g2757)
--	I6428 = NOT(g2348)
--	g7886 = NOT(g7479)
--	g4735 = NOT(g3546)
--	I17327 = NOT(g11349)
--	g6265 = NOT(I10054)
--	g3976 = NOT(I7109)
--	I6247 = NOT(g2462)
--	g4782 = NOT(g4089)
--	I11155 = NOT(g6470)
--	g10156 = NOT(I15464)
--	I15708 = NOT(g10241)
--	I17537 = NOT(g11497)
--	I13418 = NOT(g8145)
--	I13822 = NOT(g8488)
--	g5697 = NOT(I9232)
--	I10006 = NOT(g5633)
--	g6442 = NOT(I10362)
--	g9452 = NOT(I14645)
--	g7314 = NOT(I11590)
--	g5210 = NOT(I8631)
--	I17108 = NOT(g11225)
--	g11471 = NOT(I17450)
--	I7345 = NOT(g4050)
--	I16458 = NOT(g10734)
--	I8429 = NOT(g4458)
--	I9605 = NOT(g5620)
--	g4475 = NOT(I7852)
--	g5596 = NOT(I9020)
--	g6164 = NOT(g5426)
--	I7763 = NOT(g3769)
--	I7191 = NOT(g2646)
--	g10734 = NOT(I16413)
--	I10437 = NOT(g5755)
--	g10335 = NOT(I15787)
--	g7650 = NOT(I12261)
--	g3326 = NOT(I6495)
--	I15244 = NOT(g10031)
--	g4292 = NOT(g3863)
--	g10930 = NOT(g10827)
--	g11043 = NOT(I16790)
--	g6454 = NOT(I10388)
--	g11244 = NOT(g11112)
--	g4526 = NOT(I7931)
--	I5478 = NOT(g1212)
--	g6296 = NOT(I10147)
--	I11194 = NOT(g6515)
--	g3760 = NOT(g3003)
--	g7008 = NOT(I11149)
--	I13194 = NOT(g8140)
--	I13589 = NOT(g8361)
--	g2623 = NOT(g1999)
--	I17381 = NOT(g11436)
--	I7536 = NOT(g4098)
--	I9585 = NOT(g5241)
--	g2076 = NOT(I4886)
--	g10131 = NOT(I15395)
--	g2889 = NOT(I6049)
--	I11524 = NOT(g6593)
--	I16598 = NOT(g10804)
--	g11069 = NOT(g10974)
--	g4084 = NOT(g3119)
--	I11836 = NOT(g7220)
--	I5435 = NOT(g18)
--	g4603 = NOT(g3829)
--	g5936 = NOT(I9564)
--	g7336 = NOT(I11656)
--	g8600 = NOT(g8475)
--	I15068 = NOT(g9710)
--	g7768 = NOT(I12469)
--	g4439 = NOT(I7793)
--	g11657 = NOT(I17773)
--	g5117 = NOT(g4682)
--	g6553 = NOT(I10477)
--	g8714 = NOT(I14005)
--	g11068 = NOT(g10974)
--	I7858 = NOT(g3631)
--	I11477 = NOT(g6488)
--	g7594 = NOT(I12120)
--	g10487 = NOT(I16098)
--	g7972 = NOT(I12770)
--	g2175 = NOT(g44)
--	I11119 = NOT(g6461)
--	g9025 = NOT(I14412)
--	g2871 = NOT(I6013)
--	g10619 = NOT(I16292)
--	I12759 = NOT(g7702)
--	I7757 = NOT(g3767)
--	I16817 = NOT(g10912)
--	I9673 = NOT(g5182)
--	I14236 = NOT(g8802)
--	g7806 = NOT(I12583)
--	I10952 = NOT(g6556)
--	g3220 = NOT(I6398)
--	I8109 = NOT(g3622)
--	g2651 = NOT(g2007)
--	I6217 = NOT(g2302)
--	g4583 = NOT(g3880)
--	g6412 = NOT(I10322)
--	I17390 = NOT(g11430)
--	g10279 = NOT(g10158)
--	g7065 = NOT(I11272)
--	I7315 = NOT(g2891)
--	g6389 = NOT(I10289)
--	I7642 = NOT(g3440)
--	I9168 = NOT(g5040)
--	g6706 = NOT(I10685)
--	I9669 = NOT(g5426)
--	g7887 = NOT(g7693)
--	g7122 = NOT(I11357)
--	I15792 = NOT(g10279)
--	I9368 = NOT(g5288)
--	g7322 = NOT(I11614)
--	g4919 = NOT(I8290)
--	I10063 = NOT(g5766)
--	g6990 = NOT(I11132)
--	I7447 = NOT(g3694)
--	g10278 = NOT(g10182)
--	g3977 = NOT(I7112)
--	I6861 = NOT(g2942)
--	g6888 = NOT(I10984)
--	I16656 = NOT(g10791)
--	I9531 = NOT(g5004)
--	g6171 = NOT(g5446)
--	g2184 = NOT(g1806)
--	I16295 = NOT(g10552)
--	I9458 = NOT(g5091)
--	g3161 = NOT(I6367)
--	I11704 = NOT(g7008)
--	I12849 = NOT(g7632)
--	I6055 = NOT(g2569)
--	I17522 = NOT(g11485)
--	g2339 = NOT(I5399)
--	g7033 = NOT(I11188)
--	g10039 = NOT(I15244)
--	I10873 = NOT(g6331)
--	g6956 = NOT(I11106)
--	g5597 = NOT(I9023)
--	I14873 = NOT(g9525)
--	I7654 = NOT(g3728)
--	I13809 = NOT(g8480)
--	I6133 = NOT(g2253)
--	g3051 = NOT(g2135)
--	g2838 = NOT(g2165)
--	g8076 = NOT(I12930)
--	g2024 = NOT(g1718)
--	I15458 = NOT(g10069)
--	I13466 = NOT(g8160)
--	I9505 = NOT(g5088)
--	g6281 = NOT(I10102)
--	g8476 = NOT(I13674)
--	g3327 = NOT(I6498)
--	g2424 = NOT(g1690)
--	I8449 = NOT(g4469)
--	I12652 = NOT(g7458)
--	g9766 = NOT(g9432)
--	g2809 = NOT(I5909)
--	g5784 = NOT(I9380)
--	g4004 = NOT(I7140)
--	I9734 = NOT(g5257)
--	I13036 = NOT(g8053)
--	I5002 = NOT(g1173)
--	I8865 = NOT(g4518)
--	g7550 = NOT(g6974)
--	g6297 = NOT(I10150)
--	I11560 = NOT(g7037)
--	g10187 = NOT(I15539)
--	I6196 = NOT(g2462)
--	I5824 = NOT(g2502)
--	g7845 = NOT(I12634)
--	I10834 = NOT(g6715)
--	g8871 = NOT(I14185)
--	g8375 = NOT(I13475)
--	I15545 = NOT(g10075)
--	g3633 = NOT(I6802)
--	I15079 = NOT(g9745)
--	I8098 = NOT(g3583)
--	g2077 = NOT(g219)
--	g2231 = NOT(I5218)
--	g7195 = NOT(I11417)
--	g11545 = NOT(g11519)
--	g11079 = NOT(I16850)
--	g11444 = NOT(I17381)
--	g5937 = NOT(I9567)
--	g7395 = NOT(g6941)
--	I13642 = NOT(g8378)
--	g7337 = NOT(I11659)
--	g3103 = NOT(g2391)
--	I9074 = NOT(g4764)
--	g7913 = NOT(g7467)
--	I6538 = NOT(g2827)
--	g2523 = NOT(I5632)
--	I7272 = NOT(g3253)
--	g2643 = NOT(g1989)
--	I9992 = NOT(g5633)
--	g10143 = NOT(I15427)
--	g5668 = NOT(I9165)
--	g11078 = NOT(I16847)
--	g6338 = NOT(I10237)
--	I15598 = NOT(g10170)
--	I10021 = NOT(g5692)
--	g5840 = NOT(g5320)
--	g4970 = NOT(g4411)
--	g8500 = NOT(I13695)
--	I7612 = NOT(g3817)
--	g11598 = NOT(I17642)
--	I7017 = NOT(g3068)
--	g6109 = NOT(g5052)
--	I12406 = NOT(g7464)
--	g6309 = NOT(I10186)
--	g11086 = NOT(I16867)
--	g7807 = NOT(I12586)
--	I7417 = NOT(g4160)
--	g3732 = NOT(I6914)
--	I17252 = NOT(g11343)
--	g10169 = NOT(I15503)
--	I7935 = NOT(g3440)
--	I9080 = NOT(g4775)
--	g8184 = NOT(I13105)
--	g10884 = NOT(g10809)
--	g6808 = NOT(I10834)
--	I15817 = NOT(g10199)
--	I9863 = NOT(g5557)
--	g8139 = NOT(g8025)
--	I16289 = NOT(g10541)
--	g8339 = NOT(I13397)
--	g2742 = NOT(I5798)
--	g3944 = NOT(g2920)
--	g10168 = NOT(I15500)
--	I10607 = NOT(g5763)
--	g6707 = NOT(g5949)
--	I13630 = NOT(g8334)
--	g2304 = NOT(I5348)
--	g11322 = NOT(I17121)
--	g9091 = NOT(g8892)
--	g4320 = NOT(g4013)
--	I15977 = NOT(g10411)
--	g11159 = NOT(g10950)
--	I10274 = NOT(g5811)
--	I11166 = NOT(g6480)
--	I11665 = NOT(g7038)
--	I16571 = NOT(g10819)
--	I13166 = NOT(g8009)
--	I7330 = NOT(g3761)
--	I8268 = NOT(g4674)
--	g8424 = NOT(I13586)
--	I5064 = NOT(g1690)
--	g8795 = NOT(I14112)
--	g10217 = NOT(I15589)
--	g7142 = NOT(I11383)
--	I6256 = NOT(g2462)
--	g4277 = NOT(g3688)
--	g6201 = NOT(I9938)
--	g7342 = NOT(I11674)
--	I11008 = NOT(g6795)
--	g6957 = NOT(I11109)
--	I15353 = NOT(g10007)
--	g2754 = NOT(I5830)
--	g4906 = NOT(I8275)
--	g7815 = NOT(I12610)
--	g11656 = NOT(I17770)
--	g4789 = NOT(g3337)
--	I7800 = NOT(g3791)
--	g10486 = NOT(I16095)
--	g11353 = NOT(I17176)
--	g8077 = NOT(I12933)
--	I15823 = NOT(g10201)
--	g6449 = NOT(g6172)
--	I13485 = NOT(g8194)
--	g2273 = NOT(g881)
--	g8477 = NOT(g8317)
--	g6575 = NOT(g5949)
--	g7692 = NOT(g7148)
--	I12613 = NOT(g7525)
--	g8523 = NOT(I13732)
--	I6381 = NOT(g2257)
--	g9767 = NOT(I14914)
--	g7097 = NOT(I11330)
--	I9688 = NOT(g5201)
--	g7726 = NOT(I12363)
--	I9857 = NOT(g5269)
--	I13454 = NOT(g8183)
--	g2613 = NOT(I5740)
--	g7497 = NOT(g7148)
--	g9535 = NOT(I14690)
--	g6715 = NOT(I10702)
--	g2044 = NOT(I4850)
--	g7354 = NOT(I11710)
--	g10580 = NOT(g10530)
--	I10153 = NOT(g5947)
--	g2444 = NOT(g876)
--	I5237 = NOT(g1107)
--	g5032 = NOT(I8403)
--	g2269 = NOT(I5308)
--	g10223 = NOT(I15595)
--	I7213 = NOT(g2635)
--	g9261 = NOT(g8892)
--	I6421 = NOT(g2346)
--	g4299 = NOT(g4144)
--	I14409 = NOT(g8938)
--	I12463 = NOT(g7579)
--	g3697 = NOT(I6856)
--	g8099 = NOT(g7990)
--	I8385 = NOT(g4238)
--	I14136 = NOT(g8775)
--	g8304 = NOT(I13280)
--	g3914 = NOT(g3015)
--	I9126 = NOT(g4891)
--	I13239 = NOT(g8266)
--	g10110 = NOT(I15344)
--	g11631 = NOT(I17707)
--	I9326 = NOT(g5320)
--	g2543 = NOT(I5662)
--	g6584 = NOT(I10538)
--	g11017 = NOT(I16742)
--	g6539 = NOT(I10461)
--	g6896 = NOT(I10996)
--	g5568 = NOT(I8985)
--	g10321 = NOT(I15759)
--	I5089 = NOT(g1854)
--	I5731 = NOT(g2089)
--	I11238 = NOT(g6543)
--	I17213 = NOT(g11290)
--	g7783 = NOT(I12514)
--	g10179 = NOT(g10041)
--	g10531 = NOT(g10471)
--	g7979 = NOT(I12783)
--	g3413 = NOT(g2896)
--	g5912 = NOT(I9544)
--	g7312 = NOT(I11584)
--	I7166 = NOT(g2620)
--	I5966 = NOT(g2541)
--	g10178 = NOT(I15526)
--	I7366 = NOT(g4012)
--	g4738 = NOT(g3440)
--	I13941 = NOT(g8488)
--	I13382 = NOT(g8134)
--	g6268 = NOT(I10063)
--	I11519 = NOT(g6591)
--	I11176 = NOT(g6501)
--	g10186 = NOT(I15536)
--	g7001 = NOT(I11140)
--	g8273 = NOT(I13191)
--	g10676 = NOT(g10570)
--	g6419 = NOT(I10331)
--	I10891 = NOT(g6334)
--	I13185 = NOT(g8192)
--	g11289 = NOT(I17070)
--	I7456 = NOT(g3716)
--	g1993 = NOT(g786)
--	g3820 = NOT(I7048)
--	g7676 = NOT(I12303)
--	g4140 = NOT(I7284)
--	g6052 = NOT(g5426)
--	g11309 = NOT(I17096)
--	g4078 = NOT(I7205)
--	I12514 = NOT(g7735)
--	g8613 = NOT(g8484)
--	I16525 = NOT(g10719)
--	I7348 = NOT(g4056)
--	g6452 = NOT(I10384)
--	I9383 = NOT(g5296)
--	I9608 = NOT(g5127)
--	I15308 = NOT(g10019)
--	g7329 = NOT(I11635)
--	g4478 = NOT(g3820)
--	g7761 = NOT(I12448)
--	g2014 = NOT(g1104)
--	g4907 = NOT(I8278)
--	g8444 = NOT(I13630)
--	g2885 = NOT(I6043)
--	I9779 = NOT(g5391)
--	g2946 = NOT(I6133)
--	g4435 = NOT(g3914)
--	I9023 = NOT(g4727)
--	g8983 = NOT(I14370)
--	g4082 = NOT(I7213)
--	I12421 = NOT(g7634)
--	I8406 = NOT(g4274)
--	I5254 = NOT(g1700)
--	I14109 = NOT(g8765)
--	g8572 = NOT(I13809)
--	g7727 = NOT(I12366)
--	I7964 = NOT(g3433)
--	g2903 = NOT(g2166)
--	I7260 = NOT(g2844)
--	I14537 = NOT(g9308)
--	I10108 = NOT(g5743)
--	g6086 = NOT(I9737)
--	g8712 = NOT(g8680)
--	g11495 = NOT(I17500)
--	I12012 = NOT(g6916)
--	I9588 = NOT(g5114)
--	g7746 = NOT(I12403)
--	I8487 = NOT(g4526)
--	I5438 = NOT(g18)
--	g3775 = NOT(I7002)
--	g7221 = NOT(I11459)
--	I17350 = NOT(g11377)
--	I14303 = NOT(g8811)
--	g6385 = NOT(g6119)
--	g6881 = NOT(I10971)
--	I12541 = NOT(g7662)
--	g7703 = NOT(g7085)
--	I9665 = NOT(g5174)
--	I15752 = NOT(g10264)
--	g4915 = NOT(g4413)
--	g2178 = NOT(g45)
--	g2436 = NOT(I5525)
--	I15374 = NOT(g10007)
--	g9028 = NOT(I14421)
--	g8729 = NOT(g8595)
--	g8961 = NOT(I14330)
--	I4900 = NOT(g583)
--	I11501 = NOT(g6581)
--	I16610 = NOT(g10792)
--	g9671 = NOT(I14802)
--	I17152 = NOT(g11308)
--	g3060 = NOT(g2135)
--	I13729 = NOT(g8290)
--	I13577 = NOT(g8330)
--	I10381 = NOT(g5847)
--	g4214 = NOT(I7459)
--	I16255 = NOT(g10554)
--	I14982 = NOT(g9672)
--	g6425 = NOT(g6141)
--	I11728 = NOT(g7010)
--	g11643 = NOT(I17733)
--	g2135 = NOT(I5064)
--	I16679 = NOT(g10784)
--	g2335 = NOT(I5391)
--	g5683 = NOT(I9202)
--	I13439 = NOT(g8187)
--	I9346 = NOT(g5281)
--	I7118 = NOT(g2979)
--	g4310 = NOT(I7577)
--	g2382 = NOT(g599)
--	I7318 = NOT(g3266)
--	I12829 = NOT(g7680)
--	I16124 = NOT(g10396)
--	g10909 = NOT(I16679)
--	I12535 = NOT(g7656)
--	g5778 = NOT(I9368)
--	I10174 = NOT(g5994)
--	I15669 = NOT(g10194)
--	g10543 = NOT(I16196)
--	g3784 = NOT(g2586)
--	I17413 = NOT(g11425)
--	g5894 = NOT(g5361)
--	g9826 = NOT(I14979)
--	g10117 = NOT(I15359)
--	g8660 = NOT(I13945)
--	g8946 = NOT(I14295)
--	g10908 = NOT(I16676)
--	g2916 = NOT(I6097)
--	I7843 = NOT(g3440)
--	g2022 = NOT(g1346)
--	g5735 = NOT(I9293)
--	I15392 = NOT(g10104)
--	g7677 = NOT(g7148)
--	g2749 = NOT(I5815)
--	g3995 = NOT(g3121)
--	g3937 = NOT(I7086)
--	I10840 = NOT(g6719)
--	g9741 = NOT(I14888)
--	g4002 = NOT(g3121)
--	I7393 = NOT(g4096)
--	I16938 = NOT(g11086)
--	I6531 = NOT(g3186)
--	I11348 = NOT(g6695)
--	I12344 = NOT(g7062)
--	I13083 = NOT(g7921)
--	g3479 = NOT(g2655)
--	g11195 = NOT(g11112)
--	g11489 = NOT(I17482)
--	g6131 = NOT(g5548)
--	g5661 = NOT(I9144)
--	g10747 = NOT(I16432)
--	I15559 = NOT(g10094)
--	g5075 = NOT(g4439)
--	g8513 = NOT(I13708)
--	I15488 = NOT(g10116)
--	I15424 = NOT(g10080)
--	g6406 = NOT(I10314)
--	g10242 = NOT(I15632)
--	I8007 = NOT(g3829)
--	g5475 = NOT(I8892)
--	g4762 = NOT(I8116)
--	g2798 = NOT(g2449)
--	g5949 = NOT(I9591)
--	g7349 = NOT(I11695)
--	I10192 = NOT(g6115)
--	g11424 = NOT(I17327)
--	I9240 = NOT(g5069)
--	g6635 = NOT(I10592)
--	I11566 = NOT(g6820)
--	g11016 = NOT(I16739)
--	g9108 = NOT(I14449)
--	g3390 = NOT(g3161)
--	g9308 = NOT(I14499)
--	g8036 = NOT(I12878)
--	g2560 = NOT(I5684)
--	g5627 = NOT(g4840)
--	g8436 = NOT(I13606)
--	g8178 = NOT(I13083)
--	g6801 = NOT(I10813)
--	g6305 = NOT(I10174)
--	I6856 = NOT(g3318)
--	g4590 = NOT(I7999)
--	g7848 = NOT(I12641)
--	g5292 = NOT(g4445)
--	I10663 = NOT(g6040)
--	g8378 = NOT(I13482)
--	g9883 = NOT(I15060)
--	I9043 = NOT(g4786)
--	g3501 = NOT(g3077)
--	I14522 = NOT(g9108)
--	I8535 = NOT(g4340)
--	I9443 = NOT(g5557)
--	g7747 = NOT(I12406)
--	g5998 = NOT(I9620)
--	g5646 = NOT(I9099)
--	g10974 = NOT(I16723)
--	g8335 = NOT(I13385)
--	g2873 = NOT(I6019)
--	g6748 = NOT(I10753)
--	g2632 = NOT(g2002)
--	I6074 = NOT(g2228)
--	g2095 = NOT(g143)
--	I11653 = NOT(g6954)
--	g2037 = NOT(g1771)
--	g8182 = NOT(I13099)
--	I4886 = NOT(g257)
--	g4222 = NOT(g3638)
--	g5603 = NOT(I9029)
--	I6474 = NOT(g2297)
--	I7625 = NOT(g4164)
--	g5039 = NOT(I8418)
--	I4951 = NOT(g262)
--	g10293 = NOT(I15701)
--	g2653 = NOT(g2011)
--	g2208 = NOT(g84)
--	g2302 = NOT(g29)
--	I12029 = NOT(g6922)
--	g5850 = NOT(g5320)
--	g6226 = NOT(I9973)
--	I10553 = NOT(g6192)
--	g3704 = NOT(I6861)
--	g8805 = NOT(I14136)
--	g10265 = NOT(g10143)
--	g2579 = NOT(g1969)
--	I5837 = NOT(g2507)
--	I7938 = NOT(g3406)
--	I9147 = NOT(g5011)
--	I13636 = NOT(g8357)
--	g8422 = NOT(I13580)
--	I10949 = NOT(g6747)
--	I17302 = NOT(g11391)
--	g4899 = NOT(I8262)
--	I11333 = NOT(g6670)
--	I13415 = NOT(g8144)
--	g4464 = NOT(I7829)
--	g2719 = NOT(g2043)
--	g9448 = NOT(g9091)
--	I7909 = NOT(g3387)
--	I6080 = NOT(g2108)
--	I14326 = NOT(g8818)
--	g4785 = NOT(g3337)
--	g11042 = NOT(I16787)
--	g10391 = NOT(g10313)
--	I6480 = NOT(g2462)
--	g5702 = NOT(I9243)
--	g6445 = NOT(I10367)
--	g2752 = NOT(I5824)
--	I14040 = NOT(g8649)
--	I14948 = NOT(g9555)
--	g9827 = NOT(I14982)
--	g6091 = NOT(I9744)
--	I10702 = NOT(g6071)
--	g3810 = NOT(g3228)
--	g3363 = NOT(I6549)
--	I10904 = NOT(g6558)
--	g8798 = NOT(I14119)
--	g7119 = NOT(I11354)
--	g7319 = NOT(I11605)
--	g3432 = NOT(g3144)
--	I6569 = NOT(g3186)
--	g10579 = NOT(g10528)
--	g4563 = NOT(g3946)
--	g9774 = NOT(g9474)
--	I7606 = NOT(g4166)
--	g8560 = NOT(I13773)
--	I14252 = NOT(g8783)
--	g6169 = NOT(I9896)
--	I15383 = NOT(g10107)
--	I16277 = NOT(g10536)
--	g6283 = NOT(I10108)
--	g7352 = NOT(I11704)
--	g2042 = NOT(g1796)
--	g4295 = NOT(I7556)
--	g10578 = NOT(g10527)
--	I9013 = NOT(g4767)
--	g4237 = NOT(g4013)
--	g6407 = NOT(I10317)
--	I14564 = NOT(g9026)
--	g6920 = NOT(I11034)
--	g6578 = NOT(I10526)
--	g6868 = NOT(I10946)
--	g5616 = NOT(I9046)
--	I16595 = NOT(g10783)
--	g8873 = NOT(I14191)
--	g8632 = NOT(I13915)
--	g8095 = NOT(g7942)
--	g2164 = NOT(I5095)
--	g6718 = NOT(g5949)
--	g2364 = NOT(g611)
--	g2233 = NOT(I5224)
--	g9780 = NOT(g9474)
--	g4194 = NOT(I7399)
--	I16623 = NOT(g10858)
--	g8437 = NOT(I13609)
--	I10183 = NOT(g6108)
--	I7586 = NOT(g4127)
--	g11065 = NOT(g10974)
--	g4394 = NOT(I7729)
--	I5192 = NOT(g55)
--	I6976 = NOT(g2884)
--	g2054 = NOT(g1864)
--	g6582 = NOT(g5949)
--	I13609 = NOT(g8312)
--	I14397 = NOT(g8888)
--	g7386 = NOT(I11767)
--	g4731 = NOT(I8085)
--	I11312 = NOT(g6488)
--	g5647 = NOT(I9102)
--	g2454 = NOT(I5549)
--	g8579 = NOT(I13822)
--	g8869 = NOT(I14179)
--	g7975 = NOT(I12773)
--	I13200 = NOT(g8251)
--	g6261 = NOT(I10042)
--	I11608 = NOT(g6903)
--	g2296 = NOT(I5332)
--	I11115 = NOT(g6462)
--	I12604 = NOT(g7630)
--	g10116 = NOT(I15356)
--	I9117 = NOT(g5615)
--	g6793 = NOT(I10795)
--	g8719 = NOT(g8579)
--	g4557 = NOT(g3946)
--	I9317 = NOT(g5576)
--	g2725 = NOT(g2018)
--	g1974 = NOT(g627)
--	I14509 = NOT(g8926)
--	g5546 = NOT(I8973)
--	g7026 = NOT(I11173)
--	I5854 = NOT(g2523)
--	I8388 = NOT(g4239)
--	g4966 = NOT(I8340)
--	I12770 = NOT(g7638)
--	I14933 = NOT(g9454)
--	g7426 = NOT(I11814)
--	g9994 = NOT(I15196)
--	g9290 = NOT(I14494)
--	I11921 = NOT(g6904)
--	I17662 = NOT(g11602)
--	I12981 = NOT(g8041)
--	g8752 = NOT(g8635)
--	g6227 = NOT(g5446)
--	g10041 = NOT(I15250)
--	g5503 = NOT(g4515)
--	I7710 = NOT(g3749)
--	g7614 = NOT(I12190)
--	g10275 = NOT(I15669)
--	g4242 = NOT(g3664)
--	g10493 = NOT(I16114)
--	g7325 = NOT(I11623)
--	I17249 = NOT(g11342)
--	g4948 = NOT(I8315)
--	I7691 = NOT(g3363)
--	g9816 = NOT(g9490)
--	I17482 = NOT(g11479)
--	g10465 = NOT(I15986)
--	g1980 = NOT(g646)
--	I8247 = NOT(g4615)
--	g7984 = NOT(I12796)
--	g2012 = NOT(g981)
--	g11160 = NOT(g10950)
--	g8442 = NOT(I13624)
--	I17710 = NOT(g11620)
--	g6203 = NOT(g5446)
--	I17552 = NOT(g11502)
--	I16853 = NOT(g10907)
--	I9581 = NOT(g5111)
--	g10035 = NOT(I15241)
--	g5120 = NOT(I8520)
--	I5031 = NOT(g928)
--	g5320 = NOT(g4418)
--	g4254 = NOT(g4013)
--	I16589 = NOT(g10820)
--	I11674 = NOT(g7051)
--	g10806 = NOT(I16518)
--	g7544 = NOT(I11964)
--	g8164 = NOT(g7872)
--	I13674 = NOT(g8304)
--	I15470 = NOT(g10111)
--	I5812 = NOT(g2090)
--	g8233 = NOT(g7872)
--	g11617 = NOT(I17669)
--	I6183 = NOT(g2131)
--	g11470 = NOT(I17447)
--	I7659 = NOT(g3731)
--	g10142 = NOT(I15424)
--	g2888 = NOT(I6046)
--	I6924 = NOT(g2843)
--	g7636 = NOT(I12248)
--	I6220 = NOT(g883)
--	I4891 = NOT(g582)
--	g2171 = NOT(I5116)
--	g4438 = NOT(I7790)
--	I14452 = NOT(g8922)
--	g4773 = NOT(I8133)
--	g7306 = NOT(I11566)
--	I13732 = NOT(g8291)
--	g8296 = NOT(I13242)
--	g2956 = NOT(I6159)
--	I15075 = NOT(g9761)
--	g8725 = NOT(g8589)
--	g7790 = NOT(I12535)
--	g9263 = NOT(g8892)
--	g3683 = NOT(I6844)
--	g11075 = NOT(g10937)
--	I5765 = NOT(g2004)
--	I15595 = NOT(g10165)
--	I15467 = NOT(g10079)
--	I15494 = NOT(g10117)
--	I17356 = NOT(g11384)
--	g8532 = NOT(I13741)
--	I8308 = NOT(g4443)
--	g7187 = NOT(I11405)
--	I7311 = NOT(g2803)
--	g4769 = NOT(g3586)
--	g5987 = NOT(I9605)
--	I11692 = NOT(g7048)
--	g7387 = NOT(I11770)
--	g11467 = NOT(I17438)
--	I9995 = NOT(g5536)
--	I12832 = NOT(g7681)
--	I4859 = NOT(g578)
--	I10051 = NOT(g5702)
--	I10072 = NOT(g5719)
--	g4212 = NOT(I7453)
--	I9479 = NOT(g4954)
--	g6689 = NOT(g5830)
--	g10130 = NOT(I15392)
--	g7756 = NOT(I12433)
--	g2297 = NOT(g865)
--	g11623 = NOT(I17687)
--	g6388 = NOT(I10286)
--	g10193 = NOT(g10057)
--	I16616 = NOT(g10796)
--	g11037 = NOT(I16772)
--	I10592 = NOT(g5865)
--	g5299 = NOT(g4393)
--	I10756 = NOT(g5810)
--	I15782 = NOT(g10259)
--	g7622 = NOT(g7067)
--	g3735 = NOT(I6921)
--	g7027 = NOT(I11176)
--	g7427 = NOT(I11817)
--	I17182 = NOT(g11309)
--	g10165 = NOT(I15491)
--	I13400 = NOT(g8236)
--	g10523 = NOT(g10456)
--	I17672 = NOT(g11605)
--	g3782 = NOT(I7006)
--	I13013 = NOT(g8048)
--	g5892 = NOT(I9519)
--	I11214 = NOT(g6528)
--	g7904 = NOT(I12690)
--	g11419 = NOT(I17312)
--	g2745 = NOT(I5809)
--	g2639 = NOT(I5754)
--	g6030 = NOT(I9639)
--	g2338 = NOT(g1909)
--	g11352 = NOT(I17173)
--	I15418 = NOT(g10083)
--	I5073 = NOT(g34)
--	I13329 = NOT(g8116)
--	I11207 = NOT(g6524)
--	g7446 = NOT(g7148)
--	g3475 = NOT(g3056)
--	I6999 = NOT(g2905)
--	g11155 = NOT(g10950)
--	I7284 = NOT(g3255)
--	I15266 = NOT(g10001)
--	g8990 = NOT(I14391)
--	I9156 = NOT(g5032)
--	I12099 = NOT(g7258)
--	I11005 = NOT(g6386)
--	I12388 = NOT(g7219)
--	I17331 = NOT(g11357)
--	I13005 = NOT(g8046)
--	g8888 = NOT(I14232)
--	g7403 = NOT(I11783)
--	g3627 = NOT(I6784)
--	g4822 = NOT(g3706)
--	g8029 = NOT(I12871)
--	g6564 = NOT(g5784)
--	I16808 = NOT(g10906)
--	g8171 = NOT(I13068)
--	g7345 = NOT(I11683)
--	I17513 = NOT(g11482)
--	I8711 = NOT(g4530)
--	g2808 = NOT(g2156)
--	g3292 = NOT(g2373)
--	I10846 = NOT(g6729)
--	g8787 = NOT(I14094)
--	I12251 = NOT(g7076)
--	g7763 = NOT(I12454)
--	I16101 = NOT(g10381)
--	g8956 = NOT(I14319)
--	g2707 = NOT(g2041)
--	I8827 = NOT(g4477)
--	g10437 = NOT(g10333)
--	I8133 = NOT(g3632)
--	g2759 = NOT(I5843)
--	I8333 = NOT(g4456)
--	I7420 = NOT(g4167)
--	g7637 = NOT(I12251)
--	I15589 = NOT(g10161)
--	g5078 = NOT(g4372)
--	g3039 = NOT(g2310)
--	g2201 = NOT(g102)
--	g3439 = NOT(g3144)
--	g7107 = NOT(I11342)
--	I7559 = NOT(g4116)
--	g7307 = NOT(I11569)
--	I12032 = NOT(g6923)
--	g8297 = NOT(I13245)
--	g10347 = NOT(I15807)
--	g5035 = NOT(I8410)
--	I6944 = NOT(g2859)
--	I8396 = NOT(g4255)
--	g10253 = NOT(g10138)
--	I6240 = NOT(g878)
--	I7931 = NOT(g3624)
--	g7359 = NOT(I11725)
--	g6108 = NOT(I9779)
--	g6308 = NOT(I10183)
--	I9810 = NOT(g5576)
--	g5082 = NOT(g4840)
--	g2449 = NOT(g790)
--	I9032 = NOT(g4732)
--	I11100 = NOT(g6442)
--	g5482 = NOT(I8903)
--	I14405 = NOT(g8937)
--	g10600 = NOT(I16277)
--	g11401 = NOT(I17246)
--	g10781 = NOT(I16475)
--	I4783 = NOT(g873)
--	I6043 = NOT(g2267)
--	I9053 = NOT(g4752)
--	g8684 = NOT(I13969)
--	g3583 = NOT(I6742)
--	g4895 = NOT(I8250)
--	g5876 = NOT(g5361)
--	g8138 = NOT(I13013)
--	I6443 = NOT(g2363)
--	I11235 = NOT(g6538)
--	g8338 = NOT(I13394)
--	g10236 = NOT(g10190)
--	g7757 = NOT(I12436)
--	g2604 = NOT(I5713)
--	g4062 = NOT(I7185)
--	g2098 = NOT(I4938)
--	I11683 = NOT(g7069)
--	g5656 = NOT(I9129)
--	g7416 = NOT(I11800)
--	g4620 = NOT(I8031)
--	g10351 = NOT(I15817)
--	g4462 = NOT(I7825)
--	I15864 = NOT(g10339)
--	I5399 = NOT(g895)
--	g6589 = NOT(I10549)
--	I12871 = NOT(g7638)
--	g10175 = NOT(I15517)
--	g10821 = NOT(I16531)
--	I7630 = NOT(g3524)
--	I15749 = NOT(g10263)
--	g2833 = NOT(I5949)
--	I6034 = NOT(g2210)
--	g7522 = NOT(I11904)
--	I8418 = NOT(g4794)
--	g7811 = NOT(I12598)
--	g7315 = NOT(I11593)
--	g11616 = NOT(I17666)
--	I17149 = NOT(g11306)
--	I6565 = NOT(g2614)
--	g7047 = NOT(I11222)
--	I7300 = NOT(g2883)
--	g11313 = NOT(I17104)
--	I12360 = NOT(g7183)
--	I8290 = NOT(g4778)
--	g10063 = NOT(I15287)
--	I17387 = NOT(g11438)
--	g8707 = NOT(g8671)
--	g6165 = NOT(g5446)
--	g10264 = NOT(g10128)
--	g6571 = NOT(I10503)
--	g6365 = NOT(I10274)
--	g6861 = NOT(I10941)
--	g5214 = NOT(g4640)
--	g10137 = NOT(I15409)
--	g6048 = NOT(I9673)
--	I11515 = NOT(g6589)
--	g9772 = NOT(g9432)
--	I11882 = NOT(g6895)
--	I5510 = NOT(g588)
--	g2539 = NOT(I5652)
--	g2896 = NOT(g2356)
--	I6347 = NOT(g2462)
--	I15704 = NOT(g10238)
--	I5245 = NOT(g925)
--	g6448 = NOT(I10374)
--	g9531 = NOT(I14678)
--	I15305 = NOT(g10001)
--	g6711 = NOT(g5949)
--	g6055 = NOT(I9688)
--	I12162 = NOT(g7146)
--	I17104 = NOT(g11223)
--	g10873 = NOT(I16589)
--	g11053 = NOT(g10950)
--	I8256 = NOT(g4711)
--	g9890 = NOT(I15075)
--	I10282 = NOT(g6163)
--	g3404 = NOT(g3121)
--	g6133 = NOT(I9836)
--	g11466 = NOT(I17435)
--	g5663 = NOT(I9150)
--	I10302 = NOT(g6179)
--	I6914 = NOT(g2828)
--	g9505 = NOT(g9052)
--	g2162 = NOT(I5089)
--	I7973 = NOT(g3437)
--	I15036 = NOT(g9721)
--	g2268 = NOT(g654)
--	g8449 = NOT(I13645)
--	g4192 = NOT(I7393)
--	I10105 = NOT(g5736)
--	g4298 = NOT(g4130)
--	g3764 = NOT(I6971)
--	I12451 = NOT(g7538)
--	g6846 = NOT(I10910)
--	g11036 = NOT(I16769)
--	I12472 = NOT(g7539)
--	g8575 = NOT(I13816)
--	g3546 = NOT(g3307)
--	I14105 = NOT(g8776)
--	g4485 = NOT(g3546)
--	I6013 = NOT(g2200)
--	g5402 = NOT(I8842)
--	g6196 = NOT(g5446)
--	g7880 = NOT(g7479)
--	g6396 = NOT(I10296)
--	g7595 = NOT(I12123)
--	g6803 = NOT(I10819)
--	g7537 = NOT(I11947)
--	g5236 = NOT(g4361)
--	I17368 = NOT(g11423)
--	g8604 = NOT(g8479)
--	g10208 = NOT(I15580)
--	I16239 = NOT(g10525)
--	g11642 = NOT(I17730)
--	g8498 = NOT(g8353)
--	I11584 = NOT(g6827)
--	g1972 = NOT(g461)
--	I8421 = NOT(g4309)
--	g9474 = NOT(g9331)
--	g7272 = NOT(I11519)
--	I13206 = NOT(g8197)
--	g10542 = NOT(I16193)
--	g6509 = NOT(I10427)
--	g11064 = NOT(g10974)
--	I15733 = NOT(g10257)
--	g7612 = NOT(I12186)
--	g7243 = NOT(I11483)
--	g2086 = NOT(I4906)
--	I11759 = NOT(g7244)
--	I11725 = NOT(g7040)
--	I12776 = NOT(g7586)
--	g5657 = NOT(I9132)
--	g10913 = NOT(I16691)
--	I16941 = NOT(g11076)
--	g2728 = NOT(g2025)
--	I13114 = NOT(g7930)
--	g6418 = NOT(g6137)
--	I11082 = NOT(g6749)
--	g7982 = NOT(I12790)
--	g4520 = NOT(I7923)
--	g5222 = NOT(g4640)
--	I17228 = NOT(g11300)
--	g11630 = NOT(I17704)
--	g2185 = NOT(g46)
--	g4219 = NOT(g3635)
--	g6290 = NOT(I10129)
--	I7151 = NOT(g2642)
--	g2881 = NOT(I6031)
--	I7351 = NOT(g4061)
--	I16518 = NOT(g10718)
--	I6601 = NOT(g3186)
--	I7648 = NOT(g3727)
--	I12825 = NOT(g7696)
--	g10320 = NOT(I15756)
--	g10905 = NOT(I16667)
--	g7629 = NOT(I12229)
--	I15665 = NOT(g10193)
--	g7328 = NOT(I11632)
--	g2070 = NOT(g213)
--	g10530 = NOT(g10466)
--	g3906 = NOT(g3015)
--	I17716 = NOT(g11622)
--	g7330 = NOT(I11638)
--	g10593 = NOT(I16264)
--	I4866 = NOT(g579)
--	g8362 = NOT(I13466)
--	I13744 = NOT(g8297)
--	g2025 = NOT(g1696)
--	I11345 = NOT(g6692)
--	g10346 = NOT(I15804)
--	I8631 = NOT(g4425)
--	g5899 = NOT(g5361)
--	g8419 = NOT(I13571)
--	g4958 = NOT(I8328)
--	g6256 = NOT(I10027)
--	g4176 = NOT(I7345)
--	g6816 = NOT(I10858)
--	g10122 = NOT(I15374)
--	g4376 = NOT(I7691)
--	g4005 = NOT(I7143)
--	g10464 = NOT(I15983)
--	I10027 = NOT(g5751)
--	I15476 = NOT(g10114)
--	I15485 = NOT(g10092)
--	g7800 = NOT(I12565)
--	g10034 = NOT(I15238)
--	g6181 = NOT(g5426)
--	I11804 = NOT(g7190)
--	I14249 = NOT(g8804)
--	g11454 = NOT(I17419)
--	g6847 = NOT(g6482)
--	g10292 = NOT(I15698)
--	I9475 = NOT(g5445)
--	I10248 = NOT(g6125)
--	g6685 = NOT(I10648)
--	g6197 = NOT(I9930)
--	g6700 = NOT(g5949)
--	I17112 = NOT(g11227)
--	I10710 = NOT(g6088)
--	g6397 = NOT(I10299)
--	I10003 = NOT(g4908)
--	g7213 = NOT(I11447)
--	I10204 = NOT(g6031)
--	I14552 = NOT(g9264)
--	I5336 = NOT(g1700)
--	g2131 = NOT(I5060)
--	g8486 = NOT(g8348)
--	I6784 = NOT(g2742)
--	g2006 = NOT(g932)
--	g2331 = NOT(g658)
--	I16577 = NOT(g10825)
--	g4733 = NOT(I8089)
--	g2406 = NOT(g1365)
--	g5844 = NOT(I9461)
--	I13332 = NOT(g8206)
--	g6263 = NOT(I10048)
--	g4270 = NOT(g4013)
--	I11135 = NOT(g6679)
--	I7372 = NOT(g4057)
--	g10136 = NOT(I15406)
--	g2635 = NOT(g2003)
--	I16439 = NOT(g10702)
--	I17742 = NOT(g11636)
--	I12318 = NOT(g6862)
--	g11074 = NOT(g10901)
--	g6950 = NOT(I11094)
--	g11239 = NOT(g11112)
--	I10081 = NOT(g5735)
--	I17096 = NOT(g11219)
--	g4225 = NOT(I7478)
--	I15238 = NOT(g9974)
--	g2087 = NOT(g225)
--	g11594 = NOT(I17636)
--	g3945 = NOT(I7096)
--	I7143 = NOT(g2614)
--	I5943 = NOT(g2233)
--	g2801 = NOT(g2117)
--	g5089 = NOT(g4840)
--	I13406 = NOT(g8179)
--	I9084 = NOT(g4886)
--	g3738 = NOT(g3062)
--	I13962 = NOT(g8451)
--	I14786 = NOT(g9266)
--	g7512 = NOT(g7148)
--	g8025 = NOT(I12867)
--	g9760 = NOT(g9454)
--	I6294 = NOT(g2238)
--	I17681 = NOT(g11608)
--	g8425 = NOT(I13589)
--	g3709 = NOT(I6870)
--	g4124 = NOT(I7269)
--	g4324 = NOT(g4144)
--	g2748 = NOT(I5812)
--	g6562 = NOT(g5774)
--	g7366 = NOT(I11746)
--	g10164 = NOT(I15488)
--	I11833 = NOT(g7077)
--	I11049 = NOT(g6635)
--	I15675 = NOT(g10133)
--	g4469 = NOT(I7840)
--	g5705 = NOT(I9248)
--	g5471 = NOT(g4370)
--	g2755 = NOT(I5833)
--	g11185 = NOT(I16956)
--	g7056 = NOT(I11249)
--	I17730 = NOT(g11638)
--	g3907 = NOT(I7076)
--	g10891 = NOT(I16635)
--	g2226 = NOT(g86)
--	I6501 = NOT(g2578)
--	I10090 = NOT(g5767)
--	g6723 = NOT(I10716)
--	I13048 = NOT(g8059)
--	g6257 = NOT(I10030)
--	I14090 = NOT(g8771)
--	g11518 = NOT(I17563)
--	g4177 = NOT(I7348)
--	I6156 = NOT(g2119)
--	g6101 = NOT(I9762)
--	g7148 = NOT(I11397)
--	g6817 = NOT(I10861)
--	g7649 = NOT(I12258)
--	g5948 = NOT(I9588)
--	g6301 = NOT(I10162)
--	g7348 = NOT(I11692)
--	I6356 = NOT(g2459)
--	g4377 = NOT(I7694)
--	g4206 = NOT(I7435)
--	I10651 = NOT(g6035)
--	g3517 = NOT(I6702)
--	g10575 = NOT(g10523)
--	I14182 = NOT(g8788)
--	I14672 = NOT(g9261)
--	g7355 = NOT(I11713)
--	g2045 = NOT(g1811)
--	g7851 = NOT(g7479)
--	I17549 = NOT(g11501)
--	g3876 = NOT(I7061)
--	g8131 = NOT(g8020)
--	g10327 = NOT(I15771)
--	g8331 = NOT(I13373)
--	g2173 = NOT(I5120)
--	I12120 = NOT(g7106)
--	g2373 = NOT(g471)
--	g4287 = NOT(I7546)
--	I9276 = NOT(g5241)
--	g10537 = NOT(I16178)
--	I10331 = NOT(g6198)
--	g7964 = NOT(g7651)
--	g8635 = NOT(I13918)
--	g6751 = NOT(I10762)
--	I12562 = NOT(g7377)
--	I8011 = NOT(g3820)
--	I11947 = NOT(g6905)
--	g8105 = NOT(g7992)
--	g2169 = NOT(g42)
--	I5395 = NOT(g892)
--	I14449 = NOT(g8973)
--	g10283 = NOT(g10166)
--	g2369 = NOT(g617)
--	I5913 = NOT(g2169)
--	I11106 = NOT(g6667)
--	g8487 = NOT(g8350)
--	g2602 = NOT(I5707)
--	I11605 = NOT(g6834)
--	g4199 = NOT(I7414)
--	g6585 = NOT(I10541)
--	g2007 = NOT(g936)
--	g5773 = NOT(I9359)
--	g10492 = NOT(I16111)
--	g4399 = NOT(g3638)
--	g7463 = NOT(g6921)
--	g2407 = NOT(g197)
--	I6163 = NOT(g2547)
--	g2920 = NOT(g2462)
--	I14961 = NOT(g9769)
--	g2578 = NOT(g1962)
--	g2868 = NOT(I6010)
--	g3214 = NOT(I6391)
--	g4781 = NOT(I8147)
--	g6041 = NOT(I9658)
--	I6363 = NOT(g2459)
--	I7202 = NOT(g2647)
--	I15729 = NOT(g10254)
--	I13812 = NOT(g8519)
--	I9647 = NOT(g5148)
--	g4898 = NOT(I8259)
--	g6441 = NOT(g6151)
--	I13463 = NOT(g8156)
--	g9451 = NOT(I14642)
--	g4900 = NOT(I8265)
--	I6432 = NOT(g2350)
--	g11501 = NOT(I17522)
--	g3110 = NOT(g2482)
--	g11577 = NOT(I17613)
--	g7279 = NOT(g6382)
--	g5836 = NOT(g5320)
--	g4510 = NOT(I7909)
--	g11439 = NOT(I17368)
--	g3663 = NOT(I6832)
--	I12427 = NOT(g7636)
--	g10091 = NOT(I15320)
--	g9346 = NOT(I14543)
--	I12366 = NOT(g7134)
--	g2261 = NOT(g1713)
--	g7619 = NOT(I12205)
--	g7318 = NOT(I11602)
--	g2793 = NOT(g2276)
--	g4291 = NOT(g4013)
--	g7872 = NOT(I12655)
--	g11438 = NOT(I17365)
--	g10174 = NOT(I15514)
--	g10796 = NOT(I16500)
--	I16664 = NOT(g10795)
--	g9103 = NOT(g8892)
--	I8080 = NOT(g3538)
--	g2015 = NOT(g1107)
--	g6368 = NOT(g5987)
--	g8445 = NOT(I13633)
--	I7776 = NOT(g3773)
--	g7057 = NOT(I11252)
--	g2227 = NOT(g95)
--	g4344 = NOT(g3946)
--	I5142 = NOT(g639)
--	I7593 = NOT(g4142)
--	I5248 = NOT(g1110)
--	g7989 = NOT(I12805)
--	I9224 = NOT(g5063)
--	I15284 = NOT(g10034)
--	g3762 = NOT(I6965)
--	I12403 = NOT(g7611)
--	I12547 = NOT(g7673)
--	g4207 = NOT(I7438)
--	g11083 = NOT(g10913)
--	g11348 = NOT(g11276)
--	g10390 = NOT(g10309)
--	I16484 = NOT(g10770)
--	g9732 = NOT(I14873)
--	I5815 = NOT(g1994)
--	I9120 = NOT(g5218)
--	g11284 = NOT(g11208)
--	I9320 = NOT(g5013)
--	g2246 = NOT(g1810)
--	g5822 = NOT(g5320)
--	g4819 = NOT(g3354)
--	g3877 = NOT(I7064)
--	g9508 = NOT(g9271)
--	I12226 = NOT(g7066)
--	g8007 = NOT(I12843)
--	I7264 = NOT(g3252)
--	g11622 = NOT(I17684)
--	g2203 = NOT(g677)
--	g7686 = NOT(g7148)
--	g10192 = NOT(I15554)
--	I10620 = NOT(g5884)
--	I5497 = NOT(g587)
--	I6929 = NOT(g2846)
--	I12481 = NOT(g7570)
--	I13421 = NOT(g8200)
--	I16200 = NOT(g10494)
--	g8868 = NOT(I14176)
--	I5960 = NOT(g2239)
--	I7360 = NOT(g4081)
--	I14097 = NOT(g8773)
--	I9617 = NOT(g5405)
--	g6856 = NOT(I10924)
--	g6411 = NOT(g6135)
--	g6734 = NOT(I10733)
--	I9789 = NOT(g5401)
--	I10343 = NOT(g6003)
--	g8535 = NOT(I13744)
--	I7450 = NOT(g3704)
--	I10971 = NOT(g6344)
--	g7321 = NOT(I11611)
--	g8582 = NOT(I13825)
--	g7670 = NOT(I12289)
--	I17261 = NOT(g11346)
--	g4215 = NOT(I7462)
--	I7996 = NOT(g3462)
--	g11653 = NOT(I17761)
--	g2502 = NOT(I5579)
--	g4886 = NOT(I8231)
--	g4951 = NOT(I8320)
--	I16799 = NOT(g11017)
--	g7232 = NOT(I11472)
--	I12490 = NOT(g7637)
--	g10553 = NOT(I16220)
--	g8015 = NOT(I12857)
--	I15415 = NOT(g10075)
--	g5895 = NOT(g5361)
--	g7938 = NOT(g7403)
--	I8126 = NOT(g3662)
--	g7813 = NOT(I12604)
--	I5979 = NOT(g2543)
--	g4314 = NOT(g4013)
--	I5218 = NOT(g1104)
--	g5062 = NOT(g4840)
--	I13788 = NOT(g8517)
--	g9347 = NOT(I14546)
--	I12376 = NOT(g7195)
--	g10326 = NOT(I15768)
--	g5620 = NOT(g4417)
--	g7909 = NOT(g7664)
--	g2689 = NOT(g2038)
--	I12103 = NOT(g6859)
--	I11829 = NOT(g7213)
--	g6863 = NOT(g6740)
--	I16184 = NOT(g10484)
--	I16805 = NOT(g10904)
--	g10536 = NOT(I16175)
--	g8664 = NOT(I13949)
--	g10040 = NOT(I15247)
--	I10412 = NOT(g5821)
--	I12354 = NOT(g7143)
--	g2216 = NOT(g41)
--	g9533 = NOT(I14684)
--	g6713 = NOT(I10698)
--	I14412 = NOT(g8939)
--	g7519 = NOT(g6956)
--	I13828 = NOT(g8488)
--	g10904 = NOT(I16664)
--	g2028 = NOT(g1703)
--	I14133 = NOT(g8772)
--	g10252 = NOT(g10137)
--	g8721 = NOT(g8582)
--	g6569 = NOT(I10499)
--	g10621 = NOT(I16298)
--	g7606 = NOT(I12168)
--	I6894 = NOT(g2813)
--	I13344 = NOT(g8121)
--	I10228 = NOT(g6113)
--	g2247 = NOT(I5258)
--	I14228 = NOT(g8797)
--	g4336 = NOT(g4130)
--	g3394 = NOT(I6598)
--	I5830 = NOT(g2067)
--	g2564 = NOT(g1814)
--	g7687 = NOT(I12318)
--	g4768 = NOT(I8126)
--	g11576 = NOT(I17610)
--	I10716 = NOT(g6093)
--	I13682 = NOT(g8310)
--	g3731 = NOT(I6911)
--	I15554 = NOT(g10088)
--	g2826 = NOT(g2163)
--	I6661 = NOT(g2752)
--	g6688 = NOT(I10655)
--	I11173 = NOT(g6500)
--	g10183 = NOT(g10042)
--	g6857 = NOT(I10927)
--	g5192 = NOT(g4640)
--	g5085 = NOT(g4377)
--	I5221 = NOT(g1407)
--	g9820 = NOT(I14961)
--	g4943 = NOT(I8311)
--	I12190 = NOT(g7268)
--	I7674 = NOT(g3352)
--	g11200 = NOT(g11112)
--	g10062 = NOT(I15284)
--	g3705 = NOT(g3113)
--	I16214 = NOT(g10500)
--	I17271 = NOT(g11388)
--	I12520 = NOT(g7415)
--	g2638 = NOT(I5751)
--	g4065 = NOT(g2794)
--	I8161 = NOT(g3637)
--	g4887 = NOT(I8234)
--	g4228 = NOT(g3914)
--	g4322 = NOT(I7593)
--	g7570 = NOT(I12032)
--	g2108 = NOT(I4992)
--	g5941 = NOT(I9571)
--	I14379 = NOT(g8961)
--	g2609 = NOT(I5728)
--	g4934 = NOT(g4243)
--	g7341 = NOT(I11671)
--	I11029 = NOT(g6485)
--	g10851 = NOT(I16553)
--	g10872 = NOT(I16586)
--	g11052 = NOT(I16817)
--	I5932 = NOT(g2539)
--	I10958 = NOT(g6559)
--	g6400 = NOT(I10308)
--	I14112 = NOT(g8777)
--	I10378 = NOT(g6244)
--	g7525 = NOT(I11921)
--	I7680 = NOT(g3736)
--	I14958 = NOT(g9767)
--	g2883 = NOT(I6037)
--	g8671 = NOT(I13956)
--	I6484 = NOT(g2073)
--	I6439 = NOT(g2352)
--	I9915 = NOT(g5304)
--	g3254 = NOT(g2322)
--	g9775 = NOT(g9474)
--	I17736 = NOT(g11640)
--	I15798 = NOT(g10281)
--	g3814 = NOT(g3228)
--	g5708 = NOT(I9253)
--	I10096 = NOT(g5794)
--	g2217 = NOT(I5192)
--	g2758 = NOT(I5840)
--	g5520 = NOT(I8943)
--	I14944 = NOT(g9454)
--	I17198 = NOT(g11319)
--	I15184 = NOT(g9974)
--	g4096 = NOT(I7236)
--	g8564 = NOT(I13785)
--	g3038 = NOT(g1982)
--	g4496 = NOT(I7889)
--	I8303 = NOT(g4784)
--	g11184 = NOT(I16953)
--	g5252 = NOT(g4640)
--	g7607 = NOT(I12171)
--	I17528 = NOT(g11487)
--	I6702 = NOT(g2801)
--	g3773 = NOT(I6996)
--	g5812 = NOT(g5320)
--	g3009 = NOT(g2135)
--	I14681 = NOT(g9110)
--	g2165 = NOT(I5098)
--	g6183 = NOT(g5320)
--	g2571 = NOT(g1822)
--	g7659 = NOT(I12274)
--	g2861 = NOT(I6001)
--	g7358 = NOT(I11722)
--	g4195 = NOT(I7402)
--	g5176 = NOT(g4682)
--	g6220 = NOT(g5446)
--	I5716 = NOT(g2068)
--	g10574 = NOT(I16239)
--	I17764 = NOT(g11651)
--	I5149 = NOT(g1453)
--	g4395 = NOT(I7732)
--	g10047 = NOT(I15266)
--	g4337 = NOT(g4144)
--	g4913 = NOT(I8285)
--	I17365 = NOT(g11380)
--	I14802 = NOT(g9666)
--	g10205 = NOT(g10176)
--	g2055 = NOT(g1950)
--	g3769 = NOT(I6982)
--	g10912 = NOT(I16688)
--	g10311 = NOT(g10242)
--	g2455 = NOT(g826)
--	g9739 = NOT(I14884)
--	g2827 = NOT(g2164)
--	I6952 = NOT(g2867)
--	I14793 = NOT(g9269)
--	g3212 = NOT(I6385)
--	I9402 = NOT(g5107)
--	I12339 = NOT(g7054)
--	I8240 = NOT(g4380)
--	g1975 = NOT(g622)
--	I5198 = NOT(g143)
--	I12296 = NOT(g7236)
--	g7311 = NOT(I11581)
--	g2774 = NOT(g2276)
--	I6616 = NOT(g3186)
--	g3967 = NOT(g3247)
--	I17161 = NOT(g11314)
--	g6588 = NOT(I10546)
--	I4935 = NOT(g585)
--	I12644 = NOT(g7729)
--	g2846 = NOT(I5970)
--	I9762 = NOT(g5276)
--	I10549 = NOT(g6184)
--	g9079 = NOT(g8892)
--	I13648 = NOT(g8376)
--	g10051 = NOT(I15272)
--	I14690 = NOT(g9150)
--	g6161 = NOT(I9886)
--	I14549 = NOT(g9262)
--	g7615 = NOT(I12193)
--	g6361 = NOT(g5867)
--	g2196 = NOT(g91)
--	g4266 = NOT(g3688)
--	I7600 = NOT(g4159)
--	g9668 = NOT(g9490)
--	g2396 = NOT(g1389)
--	g10592 = NOT(I16261)
--	I15400 = NOT(g10069)
--	g2803 = NOT(g2154)
--	g5733 = NOT(I9287)
--	I17225 = NOT(g11298)
--	g11400 = NOT(I17243)
--	g6051 = NOT(I9680)
--	I11770 = NOT(g7202)
--	g5270 = NOT(g4367)
--	g7374 = NOT(I11752)
--	I11563 = NOT(g6819)
--	I8116 = NOT(g3627)
--	g6127 = NOT(I9826)
--	g6451 = NOT(I10381)
--	g8758 = NOT(I14055)
--	g8066 = NOT(I12916)
--	g8589 = NOT(I13834)
--	I15329 = NOT(g9995)
--	g7985 = NOT(I12799)
--	I17258 = NOT(g11345)
--	g4142 = NOT(I7288)
--	g2509 = NOT(I5588)
--	I16407 = NOT(g10696)
--	I15539 = NOT(g10069)
--	I6546 = NOT(g2987)
--	g5073 = NOT(g4840)
--	g10350 = NOT(I15814)
--	g11207 = NOT(I16982)
--	g1984 = NOT(g758)
--	I10317 = NOT(g6003)
--	g7284 = NOT(I11528)
--	g11539 = NOT(g11519)
--	g6146 = NOT(I9863)
--	g10820 = NOT(I16528)
--	g4081 = NOT(I7210)
--	g7545 = NOT(I11967)
--	g9356 = NOT(I14573)
--	g8571 = NOT(I13806)
--	I8147 = NOT(g3633)
--	g2662 = NOT(g2014)
--	g5124 = NOT(g4596)
--	g2018 = NOT(g1336)
--	g5980 = NOT(I9594)
--	g2067 = NOT(g108)
--	g7380 = NOT(g7279)
--	g8448 = NOT(I13642)
--	g6103 = NOT(I9766)
--	I10129 = NOT(g5688)
--	I9930 = NOT(g5317)
--	I11767 = NOT(g7201)
--	I11794 = NOT(g7188)
--	g8711 = NOT(g8677)
--	g7591 = NOT(I12103)
--	g6303 = NOT(I10168)
--	g2418 = NOT(I5497)
--	I11845 = NOT(g6869)
--	g5069 = NOT(g4368)
--	I13794 = NOT(g8472)
--	I10057 = NOT(g5741)
--	g4726 = NOT(g3546)
--	g2994 = NOT(g2057)
--	g5469 = NOT(I8880)
--	g7853 = NOT(I12652)
--	g4354 = NOT(I7639)
--	I5258 = NOT(g67)
--	g7020 = NOT(I11159)
--	I5818 = NOT(g2098)
--	g8133 = NOT(I13002)
--	g8333 = NOT(I13379)
--	g7420 = NOT(I11804)
--	I15241 = NOT(g10013)
--	I11898 = NOT(g6896)
--	g5177 = NOT(g4596)
--	g6732 = NOT(I10729)
--	I12867 = NOT(g7638)
--	I17657 = NOT(g11598)
--	I13633 = NOT(g8346)
--	g11241 = NOT(g11112)
--	I16206 = NOT(g10453)
--	I10299 = NOT(g6243)
--	g2256 = NOT(I5279)
--	I11191 = NOT(g6514)
--	I11719 = NOT(g7029)
--	g7559 = NOT(I12009)
--	I14323 = NOT(g8817)
--	g10691 = NOT(I16360)
--	g7794 = NOT(I12547)
--	I7076 = NOT(g2985)
--	I13191 = NOT(g8132)
--	I14299 = NOT(g8810)
--	I7889 = NOT(g3373)
--	g8196 = NOT(I13125)
--	g6944 = NOT(I11082)
--	g8803 = NOT(I14130)
--	I6277 = NOT(g1206)
--	g6072 = NOT(g4977)
--	I15771 = NOT(g10250)
--	I9237 = NOT(g5205)
--	I17337 = NOT(g11363)
--	g2181 = NOT(I5142)
--	g8538 = NOT(I13747)
--	g2381 = NOT(g1368)
--	g9432 = NOT(g9313)
--	I15235 = NOT(g9968)
--	I6789 = NOT(g2748)
--	I16114 = NOT(g10387)
--	g4783 = NOT(g3829)
--	g6043 = NOT(I9662)
--	I12910 = NOT(g7922)
--	I7375 = NOT(g4062)
--	g2847 = NOT(I5973)
--	g8780 = NOT(I14077)
--	g6443 = NOT(g6157)
--	I12202 = NOT(g6983)
--	g8509 = NOT(g8366)
--	g9453 = NOT(g9100)
--	g4112 = NOT(g2994)
--	g7905 = NOT(g7450)
--	g2197 = NOT(g101)
--	I7651 = NOT(g3332)
--	g4312 = NOT(g4144)
--	I8820 = NOT(g4473)
--	I11440 = NOT(g6577)
--	g10929 = NOT(g10827)
--	I12496 = NOT(g7724)
--	g2021 = NOT(g1341)
--	I9194 = NOT(g5236)
--	g7628 = NOT(I12226)
--	I9394 = NOT(g5195)
--	g6116 = NOT(I9801)
--	g2421 = NOT(g1374)
--	g7630 = NOT(I12232)
--	g4001 = NOT(g3200)
--	I12978 = NOT(g8040)
--	I14232 = NOT(g8800)
--	g10928 = NOT(g10827)
--	g8067 = NOT(I12919)
--	I9731 = NOT(g5255)
--	g5898 = NOT(g5361)
--	g8418 = NOT(I13568)
--	g6434 = NOT(I10352)
--	g4676 = NOT(g3354)
--	g5900 = NOT(I9531)
--	g6565 = NOT(g5790)
--	I5821 = NOT(g2101)
--	I6299 = NOT(g2242)
--	I11926 = NOT(g6900)
--	g8290 = NOT(I13224)
--	I12986 = NOT(g8042)
--	g4129 = NOT(I7280)
--	g5797 = NOT(I9399)
--	g4329 = NOT(g4144)
--	I14697 = NOT(g9260)
--	g4761 = NOT(g3440)
--	g11515 = NOT(g11490)
--	I7384 = NOT(g4082)
--	I13612 = NOT(g8325)
--	g5245 = NOT(g4369)
--	I7339 = NOT(g4004)
--	I13099 = NOT(g7927)
--	I12384 = NOT(g7212)
--	g8093 = NOT(I12948)
--	I13388 = NOT(g8230)
--	g6681 = NOT(g5830)
--	I11701 = NOT(g7065)
--	I11534 = NOT(g6917)
--	g10787 = NOT(I16487)
--	g5291 = NOT(g4384)
--	g3392 = NOT(g3121)
--	I11272 = NOT(g6546)
--	g10282 = NOT(g10164)
--	g7750 = NOT(I12415)
--	g3485 = NOT(g2662)
--	g2562 = NOT(g1383)
--	g6697 = NOT(g5949)
--	g5144 = NOT(g4682)
--	g4592 = NOT(g3829)
--	g6914 = NOT(I11024)
--	I17444 = NOT(g11446)
--	g5344 = NOT(I8811)
--	g6210 = NOT(g5205)
--	I12150 = NOT(g7074)
--	g4746 = NOT(I8098)
--	g8181 = NOT(I13096)
--	g10827 = NOT(I16543)
--	g6596 = NOT(I10566)
--	I6738 = NOT(g3113)
--	g4221 = NOT(g3914)
--	g8381 = NOT(I13489)
--	g2101 = NOT(I4951)
--	g2817 = NOT(I5919)
--	g3941 = NOT(g3015)
--	g7040 = NOT(I11207)
--	g6413 = NOT(I10325)
--	I10831 = NOT(g6710)
--	g7440 = NOT(I11836)
--	g8197 = NOT(I13128)
--	g8700 = NOT(g8574)
--	I10445 = NOT(g5770)
--	I7523 = NOT(g4095)
--	I11140 = NOT(g6448)
--	I12196 = NOT(g7272)
--	g2605 = NOT(I5716)
--	g11441 = NOT(I17374)
--	I9150 = NOT(g5012)
--	I10499 = NOT(g6149)
--	g8421 = NOT(I13577)
--	g7123 = NOT(I11360)
--	g5088 = NOT(I8456)
--	g11206 = NOT(I16979)
--	g7323 = NOT(I11617)
--	I14499 = NOT(g8889)
--	I6907 = NOT(g2994)
--	I12526 = NOT(g7648)
--	g10803 = NOT(g10708)
--	I7205 = NOT(g2632)
--	I9773 = NOT(g4934)
--	I15759 = NOT(g10267)
--	I11061 = NOT(g6641)
--	I15725 = NOT(g10251)
--	g5701 = NOT(I9240)
--	g3708 = NOT(I6867)
--	g4953 = NOT(I8324)
--	g2751 = NOT(I5821)
--	g3520 = NOT(g2779)
--	g8950 = NOT(I14303)
--	I16500 = NOT(g10711)
--	g3219 = NOT(I6395)
--	I6517 = NOT(g3271)
--	I6690 = NOT(g2743)
--	I9409 = NOT(g5013)
--	I15114 = NOT(g9875)
--	I5427 = NOT(g913)
--	g4468 = NOT(I7837)
--	I15082 = NOT(g9719)
--	g6117 = NOT(I9804)
--	I14989 = NOT(g9813)
--	I17158 = NOT(g11312)
--	g3252 = NOT(I6414)
--	g10881 = NOT(I16613)
--	I7104 = NOT(g3186)
--	g11435 = NOT(I17356)
--	I6876 = NOT(g2956)
--	I9769 = NOT(g5287)
--	g11082 = NOT(I16859)
--	g3812 = NOT(g3228)
--	I7099 = NOT(g3228)
--	I12457 = NOT(g7559)
--	I10924 = NOT(g6736)
--	g5886 = NOT(g5361)
--	g11107 = NOT(g10974)
--	I9836 = NOT(g5405)
--	I14080 = NOT(g8714)
--	g7351 = NOT(I11701)
--	g2041 = NOT(g1791)
--	g7648 = NOT(I12255)
--	g7530 = NOT(I11926)
--	I11360 = NOT(g6351)
--	g8562 = NOT(I13779)
--	I15744 = NOT(g10261)
--	I13360 = NOT(g8126)
--	I17353 = NOT(g11381)
--	g3405 = NOT(g3144)
--	g5114 = NOT(I8506)
--	I5403 = NOT(g636)
--	g9778 = NOT(g9474)
--	g5314 = NOT(g4387)
--	I11447 = NOT(g6431)
--	g11345 = NOT(I17158)
--	g9894 = NOT(I15085)
--	g8723 = NOT(g8585)
--	g4716 = NOT(g3546)
--	I11162 = NOT(g6479)
--	I16613 = NOT(g10794)
--	g11399 = NOT(I17240)
--	g3765 = NOT(g3120)
--	I10753 = NOT(g5814)
--	I10461 = NOT(g5849)
--	I5391 = NOT(g1101)
--	g3911 = NOT(g3015)
--	I9229 = NOT(g4954)
--	g7010 = NOT(I11155)
--	g6581 = NOT(I10531)
--	g10890 = NOT(I16632)
--	g5650 = NOT(I9111)
--	g7410 = NOT(I11790)
--	g9782 = NOT(I14933)
--	g11398 = NOT(I17237)
--	I15804 = NOT(g10283)
--	I16947 = NOT(g11080)
--	I5695 = NOT(g575)
--	g10249 = NOT(g10135)
--	g2168 = NOT(I5111)
--	g2669 = NOT(g2015)
--	g6060 = NOT(I9695)
--	I16273 = NOT(g10559)
--	g2368 = NOT(I5445)
--	I11629 = NOT(g6914)
--	g11652 = NOT(I17758)
--	I9822 = NOT(g5219)
--	g9661 = NOT(I14786)
--	g4198 = NOT(I7411)
--	g4747 = NOT(g3586)
--	I11472 = NOT(g6488)
--	I10736 = NOT(g6104)
--	g4398 = NOT(g3914)
--	I13451 = NOT(g8152)
--	g3733 = NOT(I6917)
--	I7444 = NOT(g3683)
--	g10248 = NOT(g10134)
--	g2772 = NOT(g2508)
--	I7269 = NOT(g2851)
--	I15263 = NOT(g9995)
--	I10198 = NOT(g6118)
--	I12300 = NOT(g7240)
--	g10552 = NOT(I16217)
--	g8751 = NOT(g8632)
--	I15332 = NOT(g10001)
--	g10204 = NOT(g10174)
--	g2743 = NOT(I5801)
--	g4241 = NOT(g3664)
--	g2890 = NOT(I6052)
--	g5768 = NOT(I9352)
--	I10843 = NOT(g6723)
--	g8585 = NOT(I13828)
--	I5858 = NOT(g2529)
--	g5594 = NOT(I9016)
--	I14528 = NOT(g9270)
--	g3473 = NOT(I6676)
--	g7278 = NOT(I11524)
--	I14330 = NOT(g8819)
--	g9526 = NOT(g9256)
--	I4938 = NOT(g261)
--	I8250 = NOT(g4589)
--	I11071 = NOT(g6656)
--	I15406 = NOT(g10065)
--	I15962 = NOT(g10405)
--	g2011 = NOT(g976)
--	g6995 = NOT(g6482)
--	g7618 = NOT(I12202)
--	g3980 = NOT(g3121)
--	g8441 = NOT(I13621)
--	g11406 = NOT(I17261)
--	g5943 = NOT(I9581)
--	g7343 = NOT(I11677)
--	g2411 = NOT(I5494)
--	I10132 = NOT(g5696)
--	g10786 = NOT(I16484)
--	g3069 = NOT(I6277)
--	I13776 = NOT(g8513)
--	I13785 = NOT(g8516)
--	g1982 = NOT(g736)
--	g4524 = NOT(g3946)
--	g6294 = NOT(I10141)
--	I15500 = NOT(g10051)
--	I5251 = NOT(g1424)
--	I6590 = NOT(g3186)
--	g3540 = NOT(g3307)
--	I7729 = NOT(g3757)
--	g5887 = NOT(I9510)
--	g10356 = NOT(I15832)
--	I5047 = NOT(g1185)
--	g5122 = NOT(g4682)
--	g11500 = NOT(I17519)
--	g6190 = NOT(g5426)
--	g2074 = NOT(g1377)
--	g4319 = NOT(g4144)
--	g7693 = NOT(I12326)
--	g11049 = NOT(I16808)
--	I11950 = NOT(g6906)
--	I16514 = NOT(g10717)
--	g10826 = NOT(I16540)
--	I9062 = NOT(g4759)
--	g7334 = NOT(I11650)
--	g10380 = NOT(I15864)
--	g3206 = NOT(g2055)
--	I13825 = NOT(g8488)
--	I13370 = NOT(g8128)
--	I9620 = NOT(g5189)
--	g4258 = NOT(I7509)
--	I16507 = NOT(g10712)
--	g4352 = NOT(I7633)
--	I11858 = NOT(g6888)
--	g11048 = NOT(I16805)
--	g4577 = NOT(I7984)
--	g4867 = NOT(I8204)
--	I14709 = NOT(g9267)
--	g5033 = NOT(I8406)
--	g10233 = NOT(g10187)
--	g6156 = NOT(g5426)
--	g4717 = NOT(g3829)
--	I7014 = NOT(g2919)
--	I12511 = NOT(g7733)
--	g10182 = NOT(I15530)
--	g7555 = NOT(I11989)
--	g7804 = NOT(I12577)
--	I7414 = NOT(g4156)
--	I10087 = NOT(g5753)
--	g9919 = NOT(I15114)
--	g2080 = NOT(I4894)
--	I7946 = NOT(g3417)
--	I10258 = NOT(g6134)
--	I14087 = NOT(g8770)
--	g7792 = NOT(I12541)
--	g2480 = NOT(I5561)
--	I11367 = NOT(g6392)
--	I11394 = NOT(g6621)
--	g5096 = NOT(g4840)
--	g6942 = NOT(I11076)
--	g8890 = NOT(I14236)
--	g2713 = NOT(g2042)
--	I13367 = NOT(g8221)
--	I13394 = NOT(g8137)
--	g4211 = NOT(I7450)
--	g4186 = NOT(I7375)
--	g6704 = NOT(g5949)
--	I17687 = NOT(g11610)
--	g4386 = NOT(I7713)
--	g10932 = NOT(g10827)
--	I8929 = NOT(g4582)
--	g5845 = NOT(g5320)
--	g4975 = NOT(I8351)
--	g2569 = NOT(I5695)
--	I7513 = NOT(g4144)
--	g8011 = NOT(I12853)
--	I17752 = NOT(g11645)
--	g5195 = NOT(g4453)
--	g5395 = NOT(I8831)
--	g5891 = NOT(g5361)
--	I9842 = NOT(g5405)
--	I17374 = NOT(g11411)
--	g7113 = NOT(I11348)
--	g11106 = NOT(g10974)
--	g7313 = NOT(I11587)
--	I11420 = NOT(g6417)
--	g4426 = NOT(g3914)
--	g10897 = NOT(g10827)
--	I12916 = NOT(g7849)
--	I10069 = NOT(g5787)
--	g6954 = NOT(I11100)
--	g6250 = NOT(I10009)
--	g4170 = NOT(g3328)
--	g6810 = NOT(I10840)
--	g4614 = NOT(g3829)
--	g9527 = NOT(I14668)
--	g4370 = NOT(I7671)
--	I12550 = NOT(g7675)
--	I7378 = NOT(g4067)
--	I10810 = NOT(g6539)
--	I11318 = NOT(g6488)
--	g4125 = NOT(I7272)
--	I15371 = NOT(g9990)
--	g6432 = NOT(g6146)
--	g7908 = NOT(g7454)
--	I13227 = NOT(g8264)
--	g6053 = NOT(I9684)
--	I14955 = NOT(g9765)
--	I17669 = NOT(g11604)
--	g8992 = NOT(I14397)
--	g9764 = NOT(g9432)
--	I16920 = NOT(g11084)
--	g11033 = NOT(I16760)
--	g3291 = NOT(g2161)
--	I12307 = NOT(g7245)
--	I5935 = NOT(g2174)
--	I6844 = NOT(g2915)
--	g6453 = NOT(g5817)
--	I9854 = NOT(g5557)
--	I14970 = NOT(g9732)
--	g4280 = NOT(g4013)
--	I7182 = NOT(g2645)
--	I7288 = NOT(g2873)
--	g4939 = NOT(I8303)
--	I11540 = NOT(g6877)
--	I5982 = NOT(g2510)
--	g3144 = NOT(g2462)
--	I11058 = NOT(g6641)
--	I15795 = NOT(g10280)
--	g3344 = NOT(I6528)
--	I16121 = NOT(g10396)
--	g6568 = NOT(g5797)
--	I10171 = NOT(g5992)
--	g4083 = NOT(I7216)
--	g8080 = NOT(I12942)
--	I4879 = NOT(g256)
--	g4544 = NOT(g3880)
--	g3207 = NOT(g2439)
--	g8573 = NOT(I13812)
--	I7916 = NOT(g3664)
--	I7022 = NOT(g2941)
--	I13203 = NOT(g8196)
--	g8480 = NOT(I13682)
--	g7776 = NOT(I12493)
--	g2000 = NOT(g810)
--	I7749 = NOT(g3764)
--	I6557 = NOT(g3086)
--	g8713 = NOT(g8684)
--	I17525 = NOT(g11486)
--	g2126 = NOT(g12)
--	g4636 = NOT(I8036)
--	I15514 = NOT(g10122)
--	I17424 = NOT(g11424)
--	g3694 = NOT(I6851)
--	g6157 = NOT(I9880)
--	I6071 = NOT(g2269)
--	I14967 = NOT(g9763)
--	I12773 = NOT(g7581)
--	I16682 = NOT(g10799)
--	I17558 = NOT(g11504)
--	I15507 = NOT(g10047)
--	g5081 = NOT(I8449)
--	I12942 = NOT(g7982)
--	g3088 = NOT(I6294)
--	g5815 = NOT(I9421)
--	g8569 = NOT(I13800)
--	g4306 = NOT(g3586)
--	g7965 = NOT(I12759)
--	I12268 = NOT(g7107)
--	g5481 = NOT(I8900)
--	g11507 = NOT(I17540)
--	I12156 = NOT(g6878)
--	g4790 = NOT(g3337)
--	I12655 = NOT(g7402)
--	g5692 = NOT(I9221)
--	I15421 = NOT(g10083)
--	g1964 = NOT(g114)
--	g10387 = NOT(g10357)
--	g97 = NOT(I4780)
--	g7264 = NOT(I11501)
--	I12180 = NOT(g7263)
--	g10620 = NOT(I16295)
--	g4187 = NOT(I7378)
--	g4061 = NOT(I7182)
--	g10148 = NOT(g10121)
--	g11421 = NOT(I17318)
--	g4387 = NOT(I7716)
--	g4461 = NOT(g3829)
--	I6955 = NOT(g2871)
--	g7360 = NOT(I11728)
--	g11163 = NOT(I16920)
--	g10104 = NOT(I15338)
--	I11146 = NOT(g6439)
--	g4756 = NOT(g3440)
--	I17713 = NOT(g11621)
--	I13738 = NOT(g8295)
--	I13645 = NOT(g8379)
--	g8688 = NOT(g8507)
--	I12335 = NOT(g7133)
--	g7521 = NOT(I11901)
--	g10343 = NOT(I15795)
--	I14010 = NOT(g8642)
--	I14918 = NOT(g9535)
--	g8976 = NOT(I14349)
--	g2608 = NOT(I5725)
--	I9829 = NOT(g5013)
--	I16760 = NOT(g10888)
--	g2220 = NOT(g104)
--	g4427 = NOT(g3638)
--	I12930 = NOT(g7896)
--	g7450 = NOT(g7148)
--	I12993 = NOT(g8044)
--	I15473 = NOT(g10087)
--	I13290 = NOT(g8254)
--	g2779 = NOT(g1974)
--	I6150 = NOT(g2122)
--	g9987 = NOT(I15187)
--	g11541 = NOT(g11519)
--	I17610 = NOT(g11549)
--	I11698 = NOT(g7057)
--	g4200 = NOT(I7417)
--	g9771 = NOT(g9432)
--	I12694 = NOT(g7374)
--	I12838 = NOT(g7682)
--	g11473 = NOT(I17456)
--	g2023 = NOT(g1357)
--	I10078 = NOT(g5729)
--	I17255 = NOT(g11344)
--	g4514 = NOT(g3946)
--	I10598 = NOT(g5874)
--	g5783 = NOT(I9377)
--	g4003 = NOT(g3144)
--	g7724 = NOT(I12357)
--	I15359 = NOT(g10019)
--	I6409 = NOT(g2356)
--	g8126 = NOT(I12989)
--	I7719 = NOT(g3752)
--	g5112 = NOT(g4682)
--	g7379 = NOT(g6863)
--	g5218 = NOT(I8647)
--	g8326 = NOT(I13360)
--	I17188 = NOT(g11313)
--	I17124 = NOT(g11232)
--	g5267 = NOT(I8711)
--	I17678 = NOT(g11607)
--	I11427 = NOT(g6573)
--	I12487 = NOT(g7723)
--	I15829 = NOT(g10203)
--	I13427 = NOT(g8241)
--	g9892 = NOT(I15079)
--	I8039 = NOT(g3506)
--	I7752 = NOT(g3407)
--	g4763 = NOT(g3586)
--	I12502 = NOT(g7726)
--	g4191 = NOT(I7390)
--	I11632 = NOT(g6931)
--	g7878 = NOT(g7479)
--	g10850 = NOT(I16550)
--	g8760 = NOT(g8670)
--	g11434 = NOT(I17353)
--	g4391 = NOT(g3638)
--	g1989 = NOT(g770)
--	I10322 = NOT(g6193)
--	g7289 = NOT(I11543)
--	g7777 = NOT(I12496)
--	g7658 = NOT(I12271)
--	g5401 = NOT(I8839)
--	g3408 = NOT(g3108)
--	I10159 = NOT(g5936)
--	g10133 = NOT(g10064)
--	g5676 = NOT(I9185)
--	g2451 = NOT(g248)
--	I10901 = NOT(g6620)
--	g4637 = NOT(I8039)
--	I12279 = NOT(g7225)
--	I5348 = NOT(g746)
--	g3336 = NOT(I6523)
--	I15344 = NOT(g10025)
--	g6778 = NOT(g5987)
--	g7882 = NOT(g7479)
--	g3768 = NOT(I6979)
--	g10896 = NOT(I16650)
--	I13403 = NOT(g8236)
--	g11344 = NOT(I17155)
--	g4307 = NOT(g4013)
--	g4536 = NOT(g3880)
--	g10228 = NOT(I15604)
--	g4159 = NOT(I7300)
--	g2346 = NOT(I5414)
--	g4359 = NOT(g3880)
--	I12469 = NOT(g7531)
--	g6735 = NOT(I10736)
--	g8183 = NOT(I13102)
--	g8608 = NOT(g8482)
--	g8924 = NOT(I14249)
--	g5830 = NOT(I9446)
--	g7611 = NOT(I12183)
--	g8220 = NOT(g7826)
--	I12286 = NOT(g7231)
--	I14561 = NOT(g9025)
--	g5727 = NOT(I9273)
--	g2103 = NOT(I4961)
--	I8919 = NOT(g4576)
--	g3943 = NOT(g2779)
--	I9177 = NOT(g4904)
--	I7233 = NOT(g2817)
--	I10144 = NOT(g5689)
--	g9340 = NOT(I14525)
--	I14295 = NOT(g8806)
--	I9377 = NOT(g5576)
--	I17219 = NOT(g11292)
--	g7799 = NOT(I12562)
--	g4757 = NOT(I8109)
--	I16604 = NOT(g10786)
--	I7054 = NOT(g3093)
--	I11572 = NOT(g6822)
--	g8423 = NOT(I13583)
--	g6475 = NOT(g5987)
--	g4416 = NOT(g3638)
--	g7981 = NOT(g7624)
--	g6949 = NOT(I11091)
--	g3228 = NOT(I6409)
--	g8977 = NOT(I14352)
--	g2732 = NOT(I5792)
--	I9287 = NOT(g5576)
--	g9082 = NOT(g8892)
--	g10310 = NOT(I15736)
--	g8588 = NOT(I13831)
--	g7997 = NOT(g7697)
--	g2753 = NOT(I5827)
--	I12601 = NOT(g7629)
--	g6292 = NOT(I10135)
--	I11127 = NOT(g6452)
--	g4315 = NOT(g3863)
--	g4811 = NOT(g3661)
--	g2508 = NOT(g940)
--	g8361 = NOT(I13463)
--	g10379 = NOT(I15861)
--	I10966 = NOT(g6561)
--	g2240 = NOT(g88)
--	I8004 = NOT(g3967)
--	g2072 = NOT(I4876)
--	g3433 = NOT(I6648)
--	I6921 = NOT(g2839)
--	I5279 = NOT(g73)
--	g7332 = NOT(I11644)
--	g10050 = NOT(I15269)
--	I9199 = NOT(g4935)
--	g10378 = NOT(I15858)
--	I8647 = NOT(g4219)
--	I9399 = NOT(g5013)
--	g5624 = NOT(I9056)
--	g7680 = NOT(g7148)
--	g11506 = NOT(I17537)
--	g7353 = NOT(I11707)
--	g2043 = NOT(g1801)
--	g6084 = NOT(I9731)
--	g8327 = NOT(g8164)
--	I14364 = NOT(g8952)
--	g4874 = NOT(I8215)
--	g6039 = NOT(I9652)
--	g5068 = NOT(g4840)
--	I11956 = NOT(g6912)
--	g3096 = NOT(g2482)
--	I13956 = NOT(g8451)
--	I13376 = NOT(g8226)
--	I13385 = NOT(g8230)
--	I11103 = NOT(g6667)
--	g3496 = NOT(I6686)
--	g7744 = NOT(I12397)
--	I11889 = NOT(g6898)
--	I17470 = NOT(g11452)
--	g7802 = NOT(I12571)
--	I5652 = NOT(g554)
--	g8146 = NOT(g8033)
--	I5057 = NOT(g1961)
--	I11354 = NOT(g6553)
--	g2116 = NOT(I5020)
--	g8346 = NOT(I13418)
--	I5843 = NOT(g2509)
--	I13354 = NOT(g8214)
--	I8503 = NOT(g4445)
--	I5989 = NOT(g2252)
--	I9510 = NOT(g5421)
--	I11824 = NOT(g7246)
--	g2034 = NOT(g1766)
--	g5677 = NOT(I9188)
--	g8103 = NOT(g7994)
--	g3395 = NOT(I6601)
--	g2434 = NOT(g1362)
--	g3337 = NOT(g2745)
--	g3913 = NOT(g2920)
--	I10289 = NOT(g6003)
--	I17277 = NOT(g11390)
--	I12168 = NOT(g7256)
--	I11671 = NOT(g7047)
--	g9310 = NOT(I14503)
--	g6583 = NOT(I10535)
--	g6702 = NOT(g5949)
--	g4880 = NOT(g3638)
--	g5866 = NOT(g5361)
--	g8696 = NOT(g8656)
--	I5549 = NOT(g868)
--	I7029 = NOT(g2946)
--	I14309 = NOT(g8813)
--	g2347 = NOT(g1945)
--	I7429 = NOT(g3344)
--	g10802 = NOT(I16510)
--	g5149 = NOT(I8551)
--	I9144 = NOT(g5007)
--	I14224 = NOT(g8794)
--	g6919 = NOT(g6453)
--	I10308 = NOT(g6003)
--	I12363 = NOT(g7187)
--	I7956 = NOT(g3428)
--	g7901 = NOT(g7712)
--	g4272 = NOT(g3586)
--	I8320 = NOT(g4452)
--	g10730 = NOT(I16407)
--	I12478 = NOT(g7560)
--	I12015 = NOT(g6924)
--	g6276 = NOT(I10087)
--	g11649 = NOT(I17749)
--	g9824 = NOT(I14973)
--	g4243 = NOT(g3524)
--	g3266 = NOT(I6436)
--	I9259 = NOT(g5301)
--	g8240 = NOT(g7972)
--	g2914 = NOT(I6091)
--	g5198 = NOT(I8614)
--	g5747 = NOT(I9317)
--	I15491 = NOT(g10093)
--	g2210 = NOT(g103)
--	g4417 = NOT(I7757)
--	I10495 = NOT(g6144)
--	g8472 = NOT(I13666)
--	g6561 = NOT(g5773)
--	g11648 = NOT(I17746)
--	g4935 = NOT(g4420)
--	g9762 = NOT(I14903)
--	I17419 = NOT(g11421)
--	I12556 = NOT(g7678)
--	I15604 = NOT(g10148)
--	I10816 = NOT(g6406)
--	I9923 = NOT(g5308)
--	g2013 = NOT(g1101)
--	g8443 = NOT(I13627)
--	g7600 = NOT(I12150)
--	I12580 = NOT(g7540)
--	g7574 = NOT(g6995)
--	I6085 = NOT(g2234)
--	g10548 = NOT(I16209)
--	I17155 = NOT(g11310)
--	g3142 = NOT(I6360)
--	g5241 = NOT(g4386)
--	g6527 = NOT(I10445)
--	I12223 = NOT(g7049)
--	g4328 = NOT(g4130)
--	I14687 = NOT(g9258)
--	I17170 = NOT(g11294)
--	I14976 = NOT(g9670)
--	g8116 = NOT(I12971)
--	g3255 = NOT(I6421)
--	I7639 = NOT(g3722)
--	g8316 = NOT(I13332)
--	g3815 = NOT(g3228)
--	I11211 = NOT(g6527)
--	I10374 = NOT(g5852)
--	g6764 = NOT(g5987)
--	I7109 = NOT(g2970)
--	I5909 = NOT(g2207)
--	I16534 = NOT(g10747)
--	I10643 = NOT(g6026)
--	I11088 = NOT(g6434)
--	I11024 = NOT(g6399)
--	g9556 = NOT(I14701)
--	I16098 = NOT(g10369)
--	g10317 = NOT(I15749)
--	g8565 = NOT(I13788)
--	g2820 = NOT(I5926)
--	g3097 = NOT(g2482)
--	I9886 = NOT(g5286)
--	I6941 = NOT(g2858)
--	g3726 = NOT(I6898)
--	g7580 = NOT(I12056)
--	g6503 = NOT(I10421)
--	g5644 = NOT(I9093)
--	I5740 = NOT(g2341)
--	g6970 = NOT(I11122)
--	g8347 = NOT(I13421)
--	I15395 = NOT(g10058)
--	g2317 = NOT(g622)
--	I8892 = NOT(g4554)
--	g10129 = NOT(I15389)
--	g9930 = NOT(I15127)
--	I9114 = NOT(g5603)
--	g6925 = NOT(I11043)
--	I17194 = NOT(g11317)
--	I7707 = NOT(g3370)
--	g11395 = NOT(I17228)
--	g1962 = NOT(g27)
--	g10057 = NOT(I15278)
--	g2601 = NOT(I5704)
--	g10128 = NOT(I15386)
--	g5818 = NOT(g5320)
--	g8697 = NOT(g8660)
--	I6520 = NOT(g3186)
--	I14668 = NOT(g9309)
--	g4213 = NOT(I7456)
--	g11633 = NOT(I17713)
--	I11659 = NOT(g7097)
--	I12186 = NOT(g7264)
--	g6120 = NOT(I9813)
--	I10195 = NOT(g6116)
--	I6031 = NOT(g2209)
--	I12953 = NOT(g8024)
--	g10323 = NOT(I15763)
--	g11191 = NOT(g11112)
--	g2775 = NOT(I5862)
--	g7076 = NOT(I11303)
--	I6812 = NOT(g3290)
--	g3783 = NOT(I7009)
--	g7476 = NOT(g6933)
--	I6958 = NOT(g2872)
--	g5893 = NOT(g5106)
--	g6277 = NOT(I10090)
--	I14525 = NOT(g9109)
--	I14424 = NOT(g8945)
--	g3112 = NOT(g2482)
--	g3267 = NOT(I6439)
--	g10775 = NOT(I16461)
--	I16766 = NOT(g10892)
--	I12936 = NOT(g7983)
--	I15832 = NOT(g10206)
--	I8340 = NOT(g4804)
--	I11296 = NOT(g6525)
--	g2060 = NOT(g1380)
--	g6617 = NOT(g6019)
--	I14558 = NOT(g9024)
--	g6789 = NOT(I10789)
--	I17749 = NOT(g11644)
--	I11644 = NOT(g6970)
--	I17616 = NOT(g11561)
--	I16871 = NOT(g10973)
--	I11338 = NOT(g6680)
--	I13338 = NOT(g8210)
--	I9594 = NOT(g5083)
--	g4166 = NOT(I7315)
--	g11440 = NOT(I17371)
--	g4366 = NOT(I7659)
--	g5426 = NOT(I8869)
--	I15861 = NOT(g10339)
--	I16360 = NOT(g10590)
--	I6911 = NOT(g2825)
--	I13969 = NOT(g8451)
--	I7833 = NOT(g3585)
--	g7285 = NOT(I11531)
--	g3329 = NOT(I6504)
--	I15247 = NOT(g10032)
--	g11573 = NOT(g11561)
--	I5525 = NOT(g589)
--	I5710 = NOT(g2431)
--	g3761 = NOT(I6962)
--	g5614 = NOT(I9040)
--	I12762 = NOT(g7541)
--	I17704 = NOT(g11618)
--	g4056 = NOT(I7173)
--	g7500 = NOT(g6943)
--	I10713 = NOT(g6003)
--	g8317 = NOT(I13335)
--	I15389 = NOT(g10110)
--	g4456 = NOT(g3375)
--	I14713 = NOT(g9052)
--	g6299 = NOT(I10156)
--	g5821 = NOT(I9433)
--	g3828 = NOT(g2920)
--	g10697 = NOT(I16370)
--	g6547 = NOT(g5893)
--	I13197 = NOT(g8186)
--	g11389 = NOT(I17216)
--	g11045 = NOT(I16796)
--	I6733 = NOT(g3321)
--	I9065 = NOT(g4760)
--	I17466 = NOT(g11447)
--	g8601 = NOT(g8477)
--	g10261 = NOT(g10126)
--	g2937 = NOT(I6106)
--	g3727 = NOT(I6901)
--	g2079 = NOT(I4891)
--	g5984 = NOT(I9602)
--	I10610 = NOT(g5879)
--	g10880 = NOT(I16610)
--	I15701 = NOT(g10236)
--	g4355 = NOT(I7642)
--	g11388 = NOT(I17213)
--	g7339 = NOT(I11665)
--	g2479 = NOT(g26)
--	I10042 = NOT(g5723)
--	I15272 = NOT(g10019)
--	I16629 = NOT(g10860)
--	g2840 = NOT(I5960)
--	I10189 = NOT(g6112)
--	g7024 = NOT(I11169)
--	I16220 = NOT(g10502)
--	g2190 = NOT(I5149)
--	g4260 = NOT(I7513)
--	g2390 = NOT(I5475)
--	g7795 = NOT(I12550)
--	I9433 = NOT(g5069)
--	I17642 = NOT(g11579)
--	I10678 = NOT(g5777)
--	g7737 = NOT(I12388)
--	g7809 = NOT(I12592)
--	g3703 = NOT(g2920)
--	I14188 = NOT(g8792)
--	I14678 = NOT(g9265)
--	g5106 = NOT(I8490)
--	g4463 = NOT(g3829)
--	I9096 = NOT(g5568)
--	g2156 = NOT(I5073)
--	g7672 = NOT(I12293)
--	I14939 = NOT(g9454)
--	g2356 = NOT(I5438)
--	g7077 = NOT(I11306)
--	g6709 = NOT(g5949)
--	I17733 = NOT(g11639)
--	g9814 = NOT(g9490)
--	g5790 = NOT(I9388)
--	I9550 = NOT(g5030)
--	I10030 = NOT(g5685)
--	g7477 = NOT(I11869)
--	I10093 = NOT(g5779)
--	I9845 = NOT(g5405)
--	g3624 = NOT(I6767)
--	g6140 = NOT(I9851)
--	g6340 = NOT(I10243)
--	I5111 = NOT(g39)
--	I11581 = NOT(g6826)
--	I11450 = NOT(g6488)
--	I12568 = NOT(g7502)
--	g9350 = NOT(I14555)
--	g10499 = NOT(I16124)
--	I5311 = NOT(g98)
--	g3068 = NOT(g2303)
--	I13714 = NOT(g8351)
--	I11315 = NOT(g6644)
--	g8784 = NOT(I14087)
--	g2942 = NOT(I6121)
--	g8739 = NOT(g8640)
--	I12242 = NOT(g7089)
--	g4279 = NOT(I7536)
--	I11707 = NOT(g7009)
--	g7205 = NOT(I11433)
--	g9773 = NOT(g9474)
--	I7086 = NOT(g3142)
--	I13819 = NOT(g8488)
--	g11061 = NOT(g10974)
--	g10498 = NOT(I16121)
--	g9009 = NOT(I14405)
--	g6435 = NOT(I10355)
--	g4167 = NOT(I7318)
--	g5027 = NOT(I8396)
--	g6517 = NOT(I10434)
--	g6082 = NOT(I9727)
--	I12123 = NOT(g6861)
--	g4318 = NOT(g4130)
--	g4367 = NOT(I7662)
--	I16859 = NOT(g10911)
--	g4872 = NOT(I8211)
--	g7634 = NOT(I12242)
--	I5174 = NOT(g52)
--	I16950 = NOT(g11081)
--	g8079 = NOT(I12939)
--	I16370 = NOT(g10592)
--	g6482 = NOT(I10412)
--	I11055 = NOT(g6419)
--	g10056 = NOT(I15275)
--	I9807 = NOT(g5419)
--	g8479 = NOT(g8319)
--	I7185 = NOT(g2626)
--	I12751 = NOT(g7626)
--	g9769 = NOT(I14918)
--	g4057 = NOT(I7176)
--	g5904 = NOT(I9539)
--	g7304 = NOT(I11560)
--	g5200 = NOT(g4567)
--	g10080 = NOT(I15308)
--	g8294 = NOT(I13236)
--	I13978 = NOT(g8575)
--	g4457 = NOT(g3829)
--	g2163 = NOT(I5092)
--	I8877 = NOT(g4421)
--	g2363 = NOT(I5441)
--	I7070 = NOT(g3138)
--	g5446 = NOT(I8877)
--	I11590 = NOT(g6829)
--	I16172 = NOT(g10498)
--	g4193 = NOT(I7396)
--	g3716 = NOT(I6876)
--	g11360 = NOT(I17185)
--	g4393 = NOT(I7726)
--	I10837 = NOT(g6717)
--	g2432 = NOT(I5513)
--	I12293 = NOT(g7116)
--	g10271 = NOT(I15665)
--	I12638 = NOT(g7708)
--	g11447 = NOT(I17390)
--	I13741 = NOT(g8296)
--	I15162 = NOT(g9958)
--	g4549 = NOT(I7956)
--	I17555 = NOT(g11503)
--	I6898 = NOT(g2964)
--	I12265 = NOT(g7211)
--	g11162 = NOT(g10950)
--	g7754 = NOT(I12427)
--	g10461 = NOT(I15974)
--	g5191 = NOT(g4640)
--	g8156 = NOT(I13051)
--	I9248 = NOT(g4954)
--	g3747 = NOT(g3015)
--	I11094 = NOT(g6657)
--	g1973 = NOT(g466)
--	g5391 = NOT(I8827)
--	g8356 = NOT(I13448)
--	g10342 = NOT(I15792)
--	g3398 = NOT(g2896)
--	g6214 = NOT(g5446)
--	g7273 = NOT(g6365)
--	I5020 = NOT(g1176)
--	I6510 = NOT(g3267)
--	g9993 = NOT(I15193)
--	g10145 = NOT(I15437)
--	g10031 = NOT(I15229)
--	g6110 = NOT(I9783)
--	g5637 = NOT(I9074)
--	g6310 = NOT(I10189)
--	g11629 = NOT(I17701)
--	g9822 = NOT(I14967)
--	g10199 = NOT(g10172)
--	g11451 = NOT(I17410)
--	g11472 = NOT(I17453)
--	g7044 = NOT(I11217)
--	g10887 = NOT(I16623)
--	g2912 = NOT(I6085)
--	I13735 = NOT(g8293)
--	g1969 = NOT(g456)
--	g4121 = NOT(I7264)
--	g5107 = NOT(g4459)
--	g8704 = NOT(g8667)
--	g4321 = NOT(g3863)
--	g2157 = NOT(g1703)
--	g11628 = NOT(I17698)
--	g10198 = NOT(I15568)
--	I7131 = NOT(g2640)
--	I7006 = NOT(g2912)
--	g7983 = NOT(I12793)
--	I10201 = NOT(g5998)
--	g5223 = NOT(g4640)
--	I11695 = NOT(g7052)
--	g10528 = NOT(g10464)
--	g10696 = NOT(g10621)
--	g4232 = NOT(I7487)
--	I12835 = NOT(g7660)
--	I13695 = NOT(g8363)
--	g10330 = NOT(I15778)
--	g5858 = NOT(I9475)
--	g10393 = NOT(g10317)
--	I10075 = NOT(g5724)
--	I7766 = NOT(g3770)
--	g8954 = NOT(I14315)
--	I16540 = NOT(g10722)
--	g6236 = NOT(I9981)
--	I6694 = NOT(g2749)
--	g7543 = NOT(I11961)
--	I12586 = NOT(g7561)
--	g11071 = NOT(g10913)
--	g8363 = NOT(I13469)
--	I7487 = NOT(g3371)
--	I8237 = NOT(g4295)
--	g5416 = NOT(I8851)
--	I14494 = NOT(g8887)
--	g3119 = NOT(I6347)
--	g10132 = NOT(g10063)
--	I17519 = NOT(g11484)
--	g10869 = NOT(I16577)
--	I6088 = NOT(g2235)
--	I17176 = NOT(g11286)
--	I17185 = NOT(g11311)
--	I10623 = NOT(g6002)
--	I12442 = NOT(g7672)
--	I17675 = NOT(g11606)
--	I17092 = NOT(g11217)
--	I16203 = NOT(g10454)
--	g4519 = NOT(I7920)
--	g5251 = NOT(g4640)
--	g6590 = NOT(g5949)
--	g6877 = NOT(I10963)
--	I4777 = NOT(g18)
--	g10868 = NOT(I16574)
--	g5811 = NOT(I9415)
--	g5642 = NOT(I9087)
--	g3352 = NOT(I6538)
--	I9783 = NOT(g5395)
--	g2626 = NOT(g2000)
--	g7534 = NOT(I11942)
--	g7729 = NOT(I12372)
--	g7961 = NOT(g7664)
--	g5047 = NOT(g4354)
--	I13457 = NOT(g8184)
--	I10984 = NOT(g6757)
--	g9895 = NOT(I15088)
--	g6657 = NOT(I10620)
--	g10161 = NOT(I15479)
--	g4552 = NOT(g3880)
--	g4606 = NOT(g3829)
--	I15858 = NOT(g10336)
--	g8568 = NOT(I13797)
--	I8089 = NOT(g3545)
--	I10352 = NOT(g6216)
--	g6556 = NOT(g5747)
--	I14352 = NOT(g8946)
--	g7927 = NOT(g7500)
--	I10822 = NOT(g6584)
--	g5874 = NOT(I9491)
--	I9001 = NOT(g4762)
--	g10259 = NOT(g10141)
--	I14418 = NOT(g8941)
--	g10708 = NOT(I16387)
--	I16739 = NOT(g10856)
--	I12430 = NOT(g7649)
--	g3186 = NOT(I6373)
--	g5654 = NOT(I9123)
--	I12493 = NOT(g7650)
--	g10471 = NOT(g10378)
--	g7414 = NOT(I11794)
--	I9293 = NOT(g5486)
--	g3386 = NOT(g3144)
--	g10087 = NOT(I15314)
--	g8357 = NOT(I13451)
--	I9129 = NOT(g4892)
--	g7946 = NOT(g7416)
--	g10258 = NOT(g10198)
--	g3975 = NOT(g3121)
--	I7173 = NOT(g2644)
--	I9329 = NOT(g5504)
--	I5973 = NOT(g2247)
--	g4586 = NOT(g4089)
--	g11394 = NOT(I17225)
--	g6464 = NOT(I10398)
--	g7903 = NOT(g7446)
--	g2683 = NOT(g2037)
--	I11689 = NOT(g7044)
--	I6870 = NOT(g2852)
--	g3274 = NOT(I6454)
--	g3426 = NOT(g3121)
--	g5880 = NOT(g5361)
--	I12035 = NOT(g6930)
--	I13280 = NOT(g8250)
--	g2778 = NOT(g2276)
--	g10244 = NOT(g10131)
--	I9727 = NOT(g5250)
--	I7369 = NOT(g4051)
--	g3370 = NOT(I6560)
--	I10589 = NOT(g5763)
--	I13624 = NOT(g8320)
--	I14194 = NOT(g8798)
--	g11420 = NOT(I17315)
--	g6563 = NOT(g5783)
--	I7920 = NOT(g3440)
--	g5272 = NOT(I8724)
--	g11319 = NOT(I17116)
--	g7036 = NOT(g6420)
--	g9085 = NOT(g8892)
--	g10069 = NOT(I15296)
--	I7459 = NOT(g3720)
--	I9221 = NOT(g5236)
--	g4525 = NOT(g3880)
--	g7436 = NOT(g7227)
--	g8626 = NOT(g8498)
--	g6295 = NOT(I10144)
--	I12517 = NOT(g7737)
--	I13102 = NOT(g7928)
--	g6237 = NOT(I9984)
--	g11446 = NOT(I17387)
--	g10774 = NOT(I16458)
--	I17438 = NOT(g11444)
--	I10477 = NOT(g6049)
--	I16366 = NOT(g10591)
--	g5417 = NOT(I8854)
--	g2075 = NOT(I4883)
--	I14477 = NOT(g8943)
--	g10879 = NOT(I16607)
--	I16632 = NOT(g10861)
--	g11059 = NOT(g10974)
--	g6844 = NOT(I10904)
--	g7335 = NOT(I11653)
--	g2475 = NOT(g192)
--	I14119 = NOT(g8779)
--	g1988 = NOT(g766)
--	g3544 = NOT(g3164)
--	g2949 = NOT(I6150)
--	g7288 = NOT(I11540)
--	g11540 = NOT(g11519)
--	g5982 = NOT(I9598)
--	g10878 = NOT(I16604)
--	I7793 = NOT(g3783)
--	I10864 = NOT(g6634)
--	g3636 = NOT(I6815)
--	g5629 = NOT(I9065)
--	I9953 = NOT(g5484)
--	g6089 = NOT(g4977)
--	I12193 = NOT(g7270)
--	g10171 = NOT(I15507)
--	g6731 = NOT(g6001)
--	I9068 = NOT(g4768)
--	g7805 = NOT(I12580)
--	I5655 = NOT(g557)
--	g7916 = NOT(g7651)
--	g11203 = NOT(g11112)
--	g5542 = NOT(I8967)
--	g7022 = NOT(g6389)
--	g3306 = NOT(I6477)
--	g2998 = NOT(g2462)
--	g2646 = NOT(g1992)
--	g4158 = NOT(g3304)
--	g7422 = NOT(I11810)
--	g7749 = NOT(I12412)
--	I6065 = NOT(g2226)
--	g6557 = NOT(g5748)
--	I12165 = NOT(g6882)
--	I12523 = NOT(g7421)
--	g10792 = NOT(I16492)
--	g11044 = NOT(I16793)
--	g3790 = NOT(g3228)
--	I15281 = NOT(g10025)
--	g2084 = NOT(I4900)
--	g2603 = NOT(I5710)
--	I8967 = NOT(g4482)
--	g6705 = NOT(I10682)
--	g2039 = NOT(g1781)
--	I9677 = NOT(g5190)
--	g3387 = NOT(I6587)
--	I10305 = NOT(g6180)
--	g5800 = NOT(I9402)
--	I5410 = NOT(g901)
--	g3461 = NOT(I6671)
--	I15377 = NOT(g10104)
--	g6242 = NOT(I9995)
--	g2850 = NOT(I5976)
--	g9431 = NOT(g9085)
--	g7798 = NOT(I12559)
--	g11301 = NOT(I17084)
--	g10459 = NOT(I15968)
--	g9812 = NOT(g9490)
--	g3756 = NOT(g3015)
--	g4587 = NOT(g3829)
--	I12475 = NOT(g7545)
--	g11377 = NOT(I17202)
--	I9866 = NOT(g5274)
--	g6948 = NOT(I11088)
--	g3622 = NOT(I6757)
--	g9958 = NOT(I15157)
--	g7560 = NOT(I12012)
--	g4275 = NOT(g3664)
--	g4311 = NOT(g4130)
--	g10458 = NOT(I15965)
--	g8782 = NOT(I14083)
--	g3427 = NOT(g3144)
--	I15562 = NOT(g10098)
--	I9349 = NOT(g5515)
--	g6955 = NOT(I11103)
--	I10036 = NOT(g5701)
--	g4615 = NOT(I8024)
--	g5213 = NOT(g4640)
--	g11645 = NOT(I17739)
--	I10177 = NOT(g6103)
--	I10560 = NOT(g5887)
--	I11456 = NOT(g6440)
--	I14101 = NOT(g8774)
--	I9848 = NOT(g5557)
--	I15290 = NOT(g9984)
--	g6254 = NOT(I10021)
--	g8475 = NOT(g8314)
--	g4174 = NOT(I7339)
--	g6814 = NOT(I10852)
--	g9765 = NOT(I14910)
--	I17636 = NOT(g11577)
--	I15698 = NOT(g10235)
--	g10545 = NOT(I16200)
--	g2919 = NOT(I6102)
--	g7037 = NOT(I11198)
--	g10079 = NOT(I15305)
--	g10444 = NOT(g10325)
--	I9699 = NOT(g5426)
--	g6150 = NOT(I9869)
--	I14642 = NOT(g9088)
--	g7437 = NOT(I11829)
--	I16784 = NOT(g10895)
--	I5667 = NOT(g566)
--	I6395 = NOT(g2334)
--	I6891 = NOT(g2962)
--	g8292 = NOT(I13230)
--	g2952 = NOT(g2455)
--	I16956 = NOT(g11096)
--	g3345 = NOT(I6531)
--	I16376 = NOT(g10596)
--	I13314 = NOT(g8260)
--	g4284 = NOT(g3664)
--	g7579 = NOT(I12053)
--	g8526 = NOT(I13735)
--	g10598 = NOT(I16273)
--	g3763 = NOT(I6968)
--	I10733 = NOT(g6099)
--	g4545 = NOT(I7952)
--	I11076 = NOT(g6649)
--	I11085 = NOT(g6433)
--	g3391 = NOT(g2896)
--	g9733 = NOT(I14876)
--	I15427 = NOT(g10088)
--	I16095 = NOT(g10401)
--	g4180 = NOT(I7357)
--	g5490 = NOT(I8911)
--	g9270 = NOT(I14485)
--	g4380 = NOT(I7701)
--	g11427 = NOT(I17334)
--	g5166 = NOT(g4682)
--	I11596 = NOT(g6831)
--	g4591 = NOT(g3829)
--	I15632 = NOT(g10184)
--	g11366 = NOT(I17191)
--	g3637 = NOT(I6818)
--	I7216 = NOT(g2952)
--	g7752 = NOT(I12421)
--	g11632 = NOT(I17710)
--	g8484 = NOT(g8336)
--	I16181 = NOT(g10491)
--	I10630 = NOT(g5889)
--	g8439 = NOT(I13615)
--	g2004 = NOT(I4820)
--	I10693 = NOT(g6068)
--	g6836 = NOT(I10888)
--	I12372 = NOT(g7137)
--	g7917 = NOT(g7497)
--	g2986 = NOT(I6220)
--	g3307 = NOT(I6480)
--	g9473 = NOT(g9103)
--	I7671 = NOT(g3351)
--	g2647 = NOT(g1993)
--	g10159 = NOT(I15473)
--	g4420 = NOT(I7766)
--	g10125 = NOT(I15377)
--	g10532 = NOT(g10473)
--	g10901 = NOT(g10802)
--	I10009 = NOT(g5542)
--	g5649 = NOT(I9108)
--	g3359 = NOT(I6543)
--	I15403 = NOT(g10069)
--	g1965 = NOT(g119)
--	g4507 = NOT(g3546)
--	g5348 = NOT(I8815)
--	g6967 = NOT(I11119)
--	I5555 = NOT(g110)
--	I11269 = NOT(g6545)
--	g9980 = NOT(I15181)
--	g2764 = NOT(I5850)
--	I8462 = NOT(g4475)
--	g11403 = NOT(I17252)
--	g10158 = NOT(I15470)
--	g11547 = NOT(g11519)
--	g7042 = NOT(I11211)
--	I11773 = NOT(g7257)
--	g10783 = NOT(I16479)
--	g4794 = NOT(I8164)
--	I11942 = NOT(g6909)
--	I13773 = NOT(g8384)
--	I5792 = NOT(g2080)
--	g7442 = NOT(g7237)
--	g8702 = NOT(g8664)
--	I13341 = NOT(g8210)
--	I12790 = NOT(g7618)
--	g7786 = NOT(I12523)
--	g2503 = NOT(g1872)
--	g3757 = NOT(I6952)
--	I9352 = NOT(g4944)
--	I17312 = NOT(g11392)
--	g10353 = NOT(I15823)
--	g3416 = NOT(g3144)
--	g6993 = NOT(I11135)
--	I11180 = NOT(g6506)
--	I16190 = NOT(g10493)
--	I14485 = NOT(g8883)
--	g7364 = NOT(I11740)
--	I6815 = NOT(g2755)
--	I9717 = NOT(g5426)
--	I15551 = NOT(g10080)
--	I14555 = NOT(g9009)
--	g3522 = NOT(g3164)
--	g8952 = NOT(I14309)
--	g11572 = NOT(g11561)
--	I11734 = NOT(g7024)
--	g8276 = NOT(I13200)
--	g3811 = NOT(I7029)
--	g2224 = NOT(g695)
--	I6097 = NOT(g2391)
--	g5063 = NOT(g4363)
--	I10914 = NOT(g6728)
--	g7454 = NOT(g7148)
--	I6726 = NOT(g3306)
--	I14570 = NOT(g9028)
--	I9893 = NOT(g5557)
--	I13335 = NOT(g8206)
--	g7770 = NOT(I12475)
--	I14914 = NOT(g9533)
--	g4515 = NOT(I7916)
--	g4204 = NOT(I7429)
--	I15127 = NOT(g9919)
--	I16546 = NOT(g10724)
--	g8561 = NOT(I13776)
--	g2320 = NOT(g18)
--	I10907 = NOT(g6705)
--	g7725 = NOT(I12360)
--	I8842 = NOT(g4556)
--	g7532 = NOT(I11932)
--	I7308 = NOT(g3070)
--	g3874 = NOT(g2920)
--	I8192 = NOT(g3566)
--	I12208 = NOT(g7124)
--	I8298 = NOT(g4437)
--	I8085 = NOT(g3664)
--	I13965 = NOT(g8451)
--	g8004 = NOT(I12838)
--	g6921 = NOT(I11037)
--	g8986 = NOT(I14379)
--	I5494 = NOT(g1690)
--	I13131 = NOT(g7979)
--	I14239 = NOT(g8803)
--	I15956 = NOT(g10402)
--	g2617 = NOT(g1997)
--	g2906 = NOT(I6071)
--	I14567 = NOT(g9027)
--	g2789 = NOT(g2276)
--	g5619 = NOT(g4840)
--	g5167 = NOT(g4682)
--	I15980 = NOT(g10414)
--	
--	g11103 = AND(g2250, g10937)
--	g9900 = AND(g9845, g8327)
--	g11095 = AND(g845, g10950)
--	g3880 = AND(g3186, g2023)
--	g4973 = AND(g1645, g4467)
--	g7389 = AND(g7001, g3880)
--	g7888 = AND(g7465, g7025)
--	g4969 = AND(g1642, g4463)
--	g8224 = AND(g1882, g7887)
--	g2892 = AND(g1980, g1976)
--	g5686 = AND(g158, g5361)
--	g10308 = AND(g10217, g9085)
--	g4123 = AND(g2695, g3037)
--	g8120 = AND(g1909, g7944)
--	g6788 = AND(g287, g5876)
--	g5598 = AND(g778, g4824)
--	g9694 = AND(g278, g9432)
--	g10495 = AND(g10431, g3971)
--	g2945 = AND(g2411, g1684)
--	g11190 = AND(g5623, g11065)
--	g8789 = AND(g8639, g8719)
--	g9852 = AND(g9728, g9563)
--	g5625 = AND(g1053, g4399)
--	g4875 = AND(g995, g3914)
--	g9701 = AND(g1574, g9474)
--	g7138 = AND(g6055, g6707)
--	g10752 = AND(g10692, g3586)
--	g11211 = AND(g11058, g5534)
--	g11024 = AND(g435, g10974)
--	g8547 = AND(g8307, g7693)
--	g10669 = AND(g10577, g9429)
--	g7707 = AND(g691, g7206)
--	g4884 = AND(g3813, g2971)
--	g4839 = AND(g225, g3946)
--	g9870 = AND(g1561, g9816)
--	g6640 = AND(g5281, g5801)
--	g9650 = AND(g2797, g9240)
--	g5687 = AND(g139, g5361)
--	g7957 = AND(g2885, g7527)
--	g3512 = AND(g2050, g2971)
--	g8244 = AND(g7847, g4336)
--	g7449 = AND(g6868, g4355)
--	g4235 = AND(g1011, g3914)
--	g4343 = AND(g345, g3586)
--	g11296 = AND(g5482, g11241)
--	g9594 = AND(g1, g9292)
--	g6829 = AND(g213, g6596)
--	g4334 = AND(g1160, g3703)
--	g9943 = AND(g9923, g9367)
--	g5525 = AND(g1721, g4292)
--	g4548 = AND(g440, g3990)
--	g8876 = AND(g8105, g6764, g8858)
--	g6733 = AND(g5678, g4324)
--	g4804 = AND(g476, g3458)
--	g10705 = AND(g10564, g4840)
--	g9934 = AND(g9913, g9624)
--	g6225 = AND(g566, g5082)
--	g6324 = AND(g1240, g5949)
--	g10686 = AND(g10612, g3863)
--	g6540 = AND(g1223, g6072)
--	g8663 = AND(g8538, g4013)
--	g11581 = AND(g1308, g11539)
--	g6206 = AND(g560, g5068)
--	g4518 = AND(g452, g3975)
--	g3989 = AND(g248, g3164)
--	g7730 = AND(g7260, g2347)
--	g5174 = AND(g1235, g4681)
--	g7504 = AND(g7148, g2847)
--	g7185 = AND(g1887, g6724)
--	g2563 = AND(I5689, I5690)
--	g7881 = AND(g7612, g3810)
--	g11070 = AND(g2008, g10913)
--	g9859 = AND(g9736, g9573)
--	g8877 = AND(g8103, g6764, g8858)
--	g11590 = AND(g2274, g11561)
--	g6199 = AND(g557, g5062)
--	g9266 = AND(g8932, g3398)
--	g5545 = AND(g1730, g4321)
--	g5180 = AND(g4541, g4533)
--	g5591 = AND(g1615, g4514)
--	g8556 = AND(g8412, g8029)
--	g11094 = AND(g374, g10883)
--	g5853 = AND(g5044, g1927)
--	g6245 = AND(g575, g5098)
--	g4360 = AND(g1861, g3748)
--	g8930 = AND(g8100, g6368, g8828)
--	g5507 = AND(g4310, g3528)
--	g11150 = AND(g3087, g10913)
--	g8464 = AND(g8302, g7416)
--	g9692 = AND(g272, g9432)
--	g4996 = AND(g1428, g4682)
--	g7131 = AND(g6044, g6700)
--	g11019 = AND(g421, g10974)
--	g9960 = AND(g9951, g9536)
--	g11196 = AND(g4912, g11068)
--	g11018 = AND(g7286, g10974)
--	g6819 = AND(g243, g6596)
--	g10595 = AND(g10550, g4347)
--	g10494 = AND(g10433, g3945)
--	g10623 = AND(g10544, g4536)
--	g4878 = AND(g1868, g3531)
--	g5204 = AND(g4838, g2126)
--	g8844 = AND(g8609, g8709)
--	g6701 = AND(g6185, g4228)
--	g10782 = AND(g10725, g5146)
--	g5100 = AND(g1791, g4606)
--	g4882 = AND(g1089, g3638)
--	g8731 = AND(g8622, g7918)
--	g6215 = AND(g1504, g5128)
--	g6886 = AND(g1932, g6420)
--	g3586 = AND(g3323, g2191)
--	g8557 = AND(g8415, g8033)
--	g8966 = AND(g8081, g6778, g8849)
--	g8071 = AND(g691, g7826)
--	g11597 = AND(g11576, g5446)
--	g9828 = AND(g9722, g9785)
--	g2918 = AND(g2411, g1672)
--	g9830 = AND(g9725, g9785)
--	g8955 = AND(g8110, g6368, g8828)
--	g9592 = AND(g4, g9292)
--	g5123 = AND(g1618, g4669)
--	g7059 = AND(g6078, g6714)
--	g8254 = AND(g2773, g7909)
--	g7459 = AND(g7148, g2814)
--	g11102 = AND(g861, g10950)
--	g7718 = AND(g709, g7221)
--	g7535 = AND(g7148, g2874)
--	g9703 = AND(g1577, g9474)
--	g5528 = AND(g4322, g3537)
--	g5151 = AND(g4478, g2733)
--	g9932 = AND(g9911, g9624)
--	g5530 = AND(g1636, g4305)
--	g3506 = AND(g986, g2760)
--	g8769 = AND(g8629, g5151)
--	g6887 = AND(g6187, g6566)
--	g6228 = AND(g5605, g713)
--	g6322 = AND(g1275, g5949)
--	g3111 = AND(I6337, I6338)
--	g8967 = AND(g8085, g6778, g8849)
--	g5010 = AND(g1458, g4640)
--	g3275 = AND(g115, g2356)
--	g10809 = AND(g4811, g10754)
--	g2895 = AND(g2411, g1678)
--	g7721 = AND(g736, g7237)
--	g9866 = AND(g1549, g9802)
--	g9716 = AND(g1534, g9490)
--	g10808 = AND(g10744, g3829)
--	g3374 = AND(g1231, g3047)
--	g4492 = AND(g1786, g3685)
--	g8822 = AND(g8614, g8752)
--	g10560 = AND(g10487, g4575)
--	g11456 = AND(g3765, g3517, g11422)
--	g9848 = AND(g9724, g9557)
--	g4714 = AND(g646, g3333)
--	g6550 = AND(g1231, g6089)
--	g5172 = AND(g4555, g4549)
--	g10642 = AND(g10612, g3829)
--	g3284 = AND(g2531, g677)
--	g9699 = AND(g284, g9432)
--	g9855 = AND(g302, g9772)
--	g5618 = AND(g1630, g4551)
--	g6891 = AND(g1950, g6435)
--	g7940 = AND(g7620, g4013)
--	g11085 = AND(g312, g10897)
--	g4736 = AND(g396, g3379)
--	g4968 = AND(g1432, g4682)
--	g8837 = AND(g8646, g8697)
--	g9644 = AND(g1182, g9125)
--	g5804 = AND(g1546, g5261)
--	g8462 = AND(g8300, g7406)
--	I6330 = AND(g2549, g2556, g2562, g2570)
--	g11156 = AND(g333, g10934)
--	g6342 = AND(g293, g5886)
--	g9867 = AND(g1552, g9807)
--	g9717 = AND(g1537, g9490)
--	g4871 = AND(g1864, g3523)
--	g10454 = AND(g10435, g3411)
--	g4722 = AND(g426, g3353)
--	g7741 = AND(g6961, g3880)
--	g4500 = AND(g1357, g3941)
--	g9386 = AND(g1327, g9151)
--	g8842 = AND(g8607, g8707)
--	g9599 = AND(g8, g9292)
--	g9274 = AND(g8974, g5708)
--	g5518 = AND(g4317, g3532)
--	g9614 = AND(g1197, g9111)
--	g4838 = AND(g3275, g4122)
--	g9125 = AND(g8966, g6674)
--	g7217 = AND(g4610, g6432)
--	g11557 = AND(g2707, g11519)
--	g2911 = AND(g2411, g1675)
--	g11210 = AND(g11078, g4515)
--	g7466 = AND(g7148, g2821)
--	g9939 = AND(g9918, g9367)
--	g11279 = AND(g4939, g11200)
--	g10518 = AND(g10513, g10440, I16145)
--	g4477 = AND(g1129, g3878)
--	g8708 = AND(g7605, g8592)
--	g7055 = AND(g5900, g6579)
--	g5264 = AND(g1095, g4763)
--	g6329 = AND(g1265, g5949)
--	g6828 = AND(g1377, g6596)
--	g8176 = AND(g5299, g7853)
--	g6830 = AND(g1380, g6596)
--	g8005 = AND(g7510, g6871)
--	g4099 = AND(g770, g3281)
--	g11601 = AND(g1351, g11574)
--	g11187 = AND(g5597, g11061)
--	g6746 = AND(g6228, g6166)
--	g6221 = AND(g782, g5598)
--	g8765 = AND(g8630, g5151)
--	g9622 = AND(g1200, g9111)
--	g11143 = AND(g10923, g4567)
--	g9904 = AND(g9886, g9676)
--	g8733 = AND(g8625, g7920)
--	g8974 = AND(g8094, g6368, g8858)
--	g6624 = AND(g348, g6171)
--	g11169 = AND(g530, g11112)
--	g8073 = AND(g709, g7826)
--	g9841 = AND(g9706, g9512)
--	g5882 = AND(g5592, g3829)
--	g8796 = AND(g8645, g8725)
--	g11168 = AND(g534, g11112)
--	g4269 = AND(g1015, g3914)
--	g5271 = AND(g727, g4772)
--	g10348 = AND(g10272, g3705)
--	g5611 = AND(g1047, g4382)
--	g8069 = AND(g673, g7826)
--	g9695 = AND(g1567, g9474)
--	g10304 = AND(g10211, g9079)
--	g8469 = AND(g8305, g7422)
--	g4712 = AND(g1071, g3638)
--	g6576 = AND(g5762, g5503)
--	g10622 = AND(g10543, g4525)
--	g11015 = AND(g5217, g10827)
--	g5674 = AND(g148, g5361)
--	g9359 = AND(g1308, g9173)
--	g9223 = AND(g6454, g8960)
--	g11556 = AND(g2701, g11519)
--	g9858 = AND(g1595, g9774)
--	g5541 = AND(g4331, g3582)
--	g4534 = AND(g363, g3586)
--	g6198 = AND(g1499, g5128)
--	g6747 = AND(g2214, g5897)
--	g6699 = AND(g6177, g4221)
--	g6855 = AND(g1964, g6392)
--	g3804 = AND(g3098, g2203)
--	g5680 = AND(g153, g5361)
--	g9642 = AND(g2654, g9240)
--	g5744 = AND(g1528, g5191)
--	g10333 = AND(g10262, g3307)
--	g8399 = AND(g6094, g8229)
--	g9447 = AND(g1762, g9030)
--	g4903 = AND(g1849, g4243)
--	g11178 = AND(g516, g11112)
--	g8510 = AND(g8414, g7972)
--	g8245 = AND(g7850, g4339)
--	g6319 = AND(g1296, g5949)
--	g11186 = AND(g5594, g11059)
--	g3908 = AND(g186, g3164)
--	g2951 = AND(g2411, g1681)
--	g6352 = AND(g278, g5894)
--	g9595 = AND(g901, g9205)
--	g4831 = AND(g810, g4109)
--	g5492 = AND(g1654, g4263)
--	g9272 = AND(g8934, g3424)
--	g10312 = AND(g10220, g9094)
--	g6186 = AND(g546, g5042)
--	g9612 = AND(g2652, g9240)
--	g9417 = AND(g1738, g9052)
--	g9935 = AND(g9914, g9624)
--	g8701 = AND(g7597, g8582)
--	g10745 = AND(g10658, g3586)
--	g11216 = AND(g956, g11162)
--	g9328 = AND(g8971, g5708)
--	g11587 = AND(g1327, g11546)
--	g6821 = AND(g237, g6596)
--	g6325 = AND(g1245, g5949)
--	g4560 = AND(g431, g4002)
--	g7368 = AND(g6980, g3880)
--	g6083 = AND(g552, g5619)
--	g6544 = AND(g1227, g6081)
--	g5476 = AND(g1615, g4237)
--	g7743 = AND(g6967, g3880)
--	g4869 = AND(g1083, g3638)
--	g5722 = AND(g1598, g5144)
--	g6790 = AND(g5813, g4398)
--	g8408 = AND(g704, g8139)
--	g10761 = AND(g10700, g10699)
--	g7734 = AND(g6944, g3880)
--	g8136 = AND(g7926, g7045)
--	g6187 = AND(g5569, g2340)
--	g4752 = AND(g401, g3385)
--	g9902 = AND(g9894, g9392)
--	g8768 = AND(g8623, g5151)
--	g5500 = AND(g1657, g4272)
--	g2496 = AND(g374, g369)
--	g6756 = AND(g3010, g5877)
--	g8972 = AND(g8085, g6764, g8858)
--	g6622 = AND(g336, g6165)
--	g11639 = AND(g11612, g7897)
--	g9366 = AND(g1311, g9173)
--	g11230 = AND(g471, g11062)
--	g10328 = AND(g10252, g3307)
--	g5024 = AND(g1284, g4513)
--	g4364 = AND(g1215, g3756)
--	g9649 = AND(g916, g9205)
--	g5795 = AND(g1543, g5251)
--	g5737 = AND(g1524, g5183)
--	g6841 = AND(g1400, g6596)
--	g4054 = AND(g1753, g2793)
--	g6345 = AND(g5823, g4426)
--	g11391 = AND(g11275, g7912)
--	g9851 = AND(g296, g9770)
--	g6763 = AND(g5802, g4381)
--	g4770 = AND(g416, g3415)
--	I16142 = AND(g10511, g10509, g10507)
--	g9698 = AND(g1571, g9474)
--	g4725 = AND(g1032, g3914)
--	g5477 = AND(g1887, g4241)
--	g9964 = AND(g9954, g9536)
--	g5523 = AND(g1663, g4290)
--	g4553 = AND(g435, g3995)
--	g8550 = AND(g8402, g8011)
--	g8845 = AND(g8611, g8711)
--	g2081 = AND(g932, g928)
--	g6359 = AND(g281, g5898)
--	g11586 = AND(g1324, g11545)
--	g11007 = AND(g5147, g10827)
--	g5104 = AND(g1796, g4608)
--	g5099 = AND(g4821, g3829)
--	g6757 = AND(g2221, g5919)
--	g5499 = AND(g1627, g4270)
--	g4389 = AND(g3529, g3092)
--	g6416 = AND(g3497, g5774)
--	g9720 = AND(g1546, g9490)
--	g4990 = AND(g1444, g4682)
--	g9619 = AND(g2772, g9010)
--	I6630 = AND(g2677, g2683, g2689, g2701)
--	g6047 = AND(g2017, g4977)
--	g9652 = AND(g953, g9223)
--	g10515 = AND(g10505, g10469, I16142)
--	g9843 = AND(g9711, g9519)
--	g5273 = AND(g1074, g4776)
--	g11465 = AND(g11434, g5446)
--	g5044 = AND(g4348, g1918)
--	g11237 = AND(g5472, g11109)
--	g9834 = AND(g9731, g9785)
--	g6654 = AND(g363, g6214)
--	g5444 = AND(g1041, g4880)
--	g3714 = AND(g1690, g2991)
--	g11340 = AND(g11285, g4424)
--	g9598 = AND(g2086, g9274)
--	g8097 = AND(g6200, g7851)
--	g8726 = AND(g8608, g7913)
--	g6880 = AND(g4816, g6562)
--	g4338 = AND(g1157, g3707)
--	g5543 = AND(g4874, g4312)
--	g8960 = AND(g8085, g6368, g8828)
--	g4109 = AND(g806, g3287)
--	g10759 = AND(g10698, g10697)
--	g9938 = AND(g9917, g9367)
--	g10758 = AND(g10652, g4013)
--	g4759 = AND(g406, g3392)
--	g9909 = AND(g9891, g9804)
--	g7127 = AND(g6663, g2241)
--	g11165 = AND(g476, g11112)
--	g6234 = AND(g2244, g5151)
--	g6328 = AND(g1260, g5949)
--	g8401 = AND(g677, g8124)
--	g11006 = AND(g5125, g10827)
--	g4865 = AND(g1080, g3638)
--	g4715 = AND(g1077, g3638)
--	g4604 = AND(g3056, g3753, g2325)
--	g5513 = AND(g1675, g4282)
--	g11222 = AND(g965, g11055)
--	g4498 = AND(g1145, g3940)
--	g6554 = AND(g5075, g6183)
--	g7732 = AND(g6935, g3880)
--	g9586 = AND(g2727, g9173)
--	g5178 = AND(g2047, g4401, g4104)
--	g4584 = AND(g3710, g2322)
--	g7472 = AND(g7148, g2829)
--	g11253 = AND(g981, g11072)
--	g5182 = AND(g1240, g4713)
--	g9860 = AND(g1598, g9775)
--	g8703 = AND(g7601, g8585)
--	g11600 = AND(g1346, g11573)
--	g9710 = AND(g1586, g9474)
--	g9645 = AND(g1203, g9111)
--	g11236 = AND(g5469, g11108)
--	g4162 = AND(g3106, g2971)
--	g6090 = AND(g553, g5627)
--	g9691 = AND(g269, g9432)
--	g11372 = AND(g11316, g4266)
--	g6823 = AND(g1368, g6596)
--	g11175 = AND(g501, g11112)
--	g8068 = AND(g664, g7826)
--	g9607 = AND(g12, g9274)
--	g9962 = AND(g9952, g9536)
--	g6348 = AND(g296, g5891)
--	g9659 = AND(g956, g9223)
--	g9358 = AND(g1318, g9151)
--	g3104 = AND(I6316, I6317)
--	g4486 = AND(g1711, g3910)
--	g9587 = AND(g892, g8995)
--	g5632 = AND(g1636, g4563)
--	g9111 = AND(g8965, g6674)
--	g4881 = AND(g991, g3914)
--	g11209 = AND(g11074, g9448)
--	g8848 = AND(g8715, g8713)
--	g4070 = AND(g3263, g2330)
--	g6463 = AND(g5052, g6210)
--	g8699 = AND(g7595, g8579)
--	I5689 = AND(g1419, g1424, g1428, g1432)
--	g7820 = AND(g1896, g7479)
--	g11021 = AND(g448, g10974)
--	g5917 = AND(g1044, g5320)
--	g6619 = AND(g49, g6156)
--	g6318 = AND(g1300, g5949)
--	g6872 = AND(g1896, g6389)
--	g11320 = AND(g11201, g4379)
--	g10514 = AND(g10489, g4580)
--	g4006 = AND(g201, g3228)
--	g9853 = AND(g299, g9771)
--	g11274 = AND(g4913, g11197)
--	g6193 = AND(g2206, g5151)
--	g8119 = AND(g6239, g7890)
--	g9420 = AND(g1747, g9030)
--	g5233 = AND(g1791, g4492)
--	g7581 = AND(g7092, g5420)
--	g6549 = AND(g5515, g6175)
--	g11464 = AND(g11433, g5446)
--	g4801 = AND(g516, g3439)
--	g6834 = AND(g1365, g6596)
--	g4487 = AND(g1718, g3911)
--	g2939 = AND(g2411, g1687)
--	g7060 = AND(g6739, g5521)
--	g5770 = AND(g4466, g5128)
--	g5725 = AND(g1580, g5166)
--	g11641 = AND(g11615, g7901)
--	g2544 = AND(g1341, g1336)
--	g11292 = AND(g11252, g4250)
--	g5532 = AND(g1681, g4307)
--	g11153 = AND(g3771, g10913)
--	g9905 = AND(g9872, g9680)
--	g7739 = AND(g6957, g3880)
--	g6321 = AND(g1284, g5949)
--	g8386 = AND(g6085, g8219)
--	g8975 = AND(g8089, g6764, g8858)
--	g2306 = AND(g1223, g1218)
--	g6625 = AND(g1218, g6178)
--	g7937 = AND(g7606, g4013)
--	g10788 = AND(g8303, g10754)
--	g10325 = AND(g10248, g3307)
--	g8170 = AND(g5270, g7853)
--	g5706 = AND(g1574, g5121)
--	g2756 = AND(g936, g2081)
--	g8821 = AND(g8643, g8751)
--	g10946 = AND(g5225, g10827)
--	g4169 = AND(g2765, g3066)
--	g5029 = AND(g1077, g4521)
--	g11164 = AND(g4889, g11112)
--	g4007 = AND(g2683, g2276)
--	g4059 = AND(g1756, g2796)
--	g4868 = AND(g1027, g3914)
--	g5675 = AND(g131, g5361)
--	g4718 = AND(g650, g3343)
--	g10682 = AND(g10600, g3863)
--	g6687 = AND(g5486, g5840)
--	g7704 = AND(g682, g7197)
--	g4582 = AND(g525, g4055)
--	g4261 = AND(g1019, g3914)
--	g3422 = AND(g225, g3228)
--	g5745 = AND(g1549, g5192)
--	g8387 = AND(g6086, g8220)
--	g7954 = AND(g2874, g7512)
--	g11283 = AND(g4966, g11205)
--	g8461 = AND(g8298, g7403)
--	g10760 = AND(g10695, g10691)
--	g11492 = AND(g11480, g4807)
--	g7032 = AND(g2965, g6626, g5292)
--	g8756 = AND(g7431, g8674)
--	g9151 = AND(g8967, g6674)
--	g6341 = AND(g272, g5885)
--	g10506 = AND(g10390, g2135)
--	g9648 = AND(g16, g9274)
--	g7453 = AND(g7148, g2809)
--	g6525 = AND(g5995, g3102)
--	g6645 = AND(g67, g6202)
--	g5707 = AND(g1595, g5122)
--	g8046 = AND(g7548, g5128)
--	g11091 = AND(g833, g10950)
--	g11174 = AND(g496, g11112)
--	g9010 = AND(g6454, g8930)
--	g8403 = AND(g6101, g8239)
--	g5201 = AND(g1250, g4721)
--	g8841 = AND(g8605, g8704)
--	g6879 = AND(g1914, g6407)
--	g8763 = AND(g7440, g8680)
--	g4502 = AND(g2031, g3938)
--	g9839 = AND(g9702, g9742)
--	g6358 = AND(g5841, g4441)
--	g5575 = AND(g1618, g4501)
--	g4940 = AND(g3500, g4440)
--	g8107 = AND(g6226, g7882)
--	g10240 = AND(g10150, g9103)
--	g11192 = AND(g5628, g11066)
--	g9618 = AND(g910, g9205)
--	g5539 = AND(g1684, g4314)
--	g8416 = AND(g731, g8151)
--	g9693 = AND(g275, g9432)
--	g11553 = AND(g2683, g11519)
--	g8047 = AND(g7557, g5919)
--	g5268 = AND(g1098, g4769)
--	g9555 = AND(g9107, g3391)
--	g6180 = AND(g2190, g5128)
--	g6832 = AND(g1383, g6596)
--	g10633 = AND(g10600, g3829)
--	g7894 = AND(g7617, g3816)
--	g8654 = AND(g8529, g4013)
--	g9621 = AND(g1179, g9125)
--	g6794 = AND(g5819, g4415)
--	g9313 = AND(g8876, g5708)
--	g4883 = AND(g248, g3946)
--	g3412 = AND(g219, g3228)
--	g7661 = AND(g7127, g2251)
--	g2800 = AND(g2399, g2369, g591)
--	g3389 = AND(g207, g3228)
--	g3706 = AND(g471, g3268)
--	g9908 = AND(g9890, g9782)
--	g3429 = AND(g231, g3228)
--	g6628 = AND(g351, g6182)
--	g5470 = AND(g1044, g4222)
--	g7526 = AND(g7148, g2868)
--	g5897 = AND(g2204, g5354)
--	g5025 = AND(g1482, g4640)
--	g6204 = AND(g3738, g4921)
--	g4048 = AND(g1750, g2790)
--	g8935 = AND(g8106, g6778, g8849)
--	g3281 = AND(g766, g2525)
--	g9593 = AND(g898, g9205)
--	g4827 = AND(g213, g3946)
--	g10701 = AND(g10620, g10619)
--	g10777 = AND(g10733, g3015)
--	g8130 = AND(g1936, g7952)
--	g9965 = AND(g9955, g9536)
--	g3684 = AND(g1710, g3015)
--	g11213 = AND(g947, g11157)
--	g5006 = AND(g1462, g4640)
--	g9933 = AND(g9912, g9624)
--	g8554 = AND(g8407, g8020)
--	g9641 = AND(g913, g9205)
--	g6123 = AND(g5630, g4311)
--	g6323 = AND(g1235, g5949)
--	g10766 = AND(g10646, g4840)
--	g6666 = AND(g5301, g5818)
--	g4994 = AND(g1504, g4640)
--	g5755 = AND(g5103, g5354)
--	g11592 = AND(g3717, g11561)
--	g6351 = AND(g6210, g5052)
--	g6875 = AND(g1905, g6400)
--	g4816 = AND(g4070, g2336)
--	g9658 = AND(g947, g9240)
--	g6530 = AND(g6207, g3829)
--	g8366 = AND(g8199, g7265)
--	g9835 = AND(g9735, g9785)
--	g6655 = AND(g5296, g5812)
--	g5445 = AND(g4631, g3875, g2733)
--	g5173 = AND(g3094, g4676)
--	g7970 = AND(g7384, g7703)
--	g3098 = AND(g2331, g2198)
--	g5491 = AND(g1624, g4262)
--	g9271 = AND(g6681, g8949)
--	g11152 = AND(g369, g10903)
--	g9611 = AND(g2651, g9010)
--	g6410 = AND(g2804, g5759)
--	g10451 = AND(g10444, g3365)
--	g4397 = AND(g3475, g2181)
--	g7224 = AND(g5398, g6441)
--	g5602 = AND(g1624, g4535)
--	g4421 = AND(g4112, g2980)
--	g6884 = AND(g5569, g6564)
--	g6839 = AND(g1397, g6596)
--	g8698 = AND(g7591, g8576)
--	g8964 = AND(g8255, g6368, g8849)
--	g8260 = AND(g2775, g7911)
--	g11413 = AND(g11354, g10679)
--	g4950 = AND(g1415, g4682)
--	g5535 = AND(g4327, g3544)
--	g7277 = AND(g6772, g731)
--	g8463 = AND(g8301, g7410)
--	g3268 = AND(g466, g2511)
--	g10785 = AND(g10728, g5177)
--	g6618 = AND(g658, g6016)
--	g6235 = AND(g569, g5089)
--	g10950 = AND(g10788, g6355)
--	g4723 = AND(g3626, g2779)
--	g8720 = AND(g8601, g7905)
--	g6693 = AND(g5494, g5845)
--	g11020 = AND(g452, g10974)
--	g11583 = AND(g1314, g11541)
--	g8118 = AND(g1900, g7941)
--	g8167 = AND(g5253, g7853)
--	g6334 = AND(g1389, g5904)
--	g7892 = AND(g7616, g3815)
--	g8652 = AND(g8523, g4013)
--	g5721 = AND(g1577, g5143)
--	g10367 = AND(g10362, g3375)
--	g9901 = AND(g9893, g9392)
--	g6792 = AND(g290, g5881)
--	g11282 = AND(g4958, g11203)
--	g7945 = AND(g2847, g7473)
--	g8971 = AND(g8081, g6764, g8858)
--	g11302 = AND(g5508, g11244)
--	g4585 = AND(g521, g4060)
--	g6621 = AND(g52, g6164)
--	g5502 = AND(g1932, g4275)
--	g11105 = AND(g3634, g10937)
--	g7709 = AND(g6856, g4333)
--	g8598 = AND(g8471, g7432)
--	g7140 = AND(g6069, g6711)
--	g9600 = AND(g904, g9205)
--	g9864 = AND(g1604, g9778)
--	g11640 = AND(g11613, g7900)
--	g5188 = AND(g4504, g4496)
--	g7435 = AND(g7260, g6572)
--	g7876 = AND(g7609, g3790)
--	g5030 = AND(g1280, g4523)
--	g4058 = AND(g2707, g2276)
--	g6776 = AND(g5809, g4390)
--	g4890 = AND(g630, g4739)
--	g2525 = AND(g762, g758)
--	g10301 = AND(g8892, g10223)
--	g4505 = AND(g354, g3586)
--	g9623 = AND(g17, g9274)
--	g10739 = AND(g10676, g3368)
--	g11027 = AND(g391, g10974)
--	g10738 = AND(g10692, g4840)
--	g8687 = AND(g8558, g8036)
--	g6360 = AND(g302, g5899)
--	g9871 = AND(g1564, g9668)
--	g5108 = AND(g1801, g4614)
--	g11248 = AND(g976, g11071)
--	g4992 = AND(g1407, g4682)
--	g11552 = AND(g2677, g11519)
--	g9651 = AND(g944, g9240)
--	g11204 = AND(g971, g11083)
--	g7824 = AND(g1932, g7479)
--	g4480 = AND(g1133, g3905)
--	g6179 = AND(g5115, g5354)
--	g8710 = AND(g7607, g8595)
--	g7590 = AND(g7102, g5425)
--	g9384 = AND(g968, g9223)
--	g3407 = AND(g2561, g3012)
--	g9838 = AND(g9700, g9754)
--	g3718 = AND(g192, g3164)
--	g10661 = AND(g10594, g3015)
--	g11380 = AND(g11321, g4285)
--	g8879 = AND(g8110, g6764, g8858)
--	g7930 = AND(g7621, g3110)
--	g8962 = AND(g8089, g6368, g8828)
--	g10715 = AND(g2272, g10630)
--	g8659 = AND(g8535, g4013)
--	g3015 = AND(g2028, g2191)
--	g9643 = AND(g950, g9223)
--	g9205 = AND(g6454, g8957)
--	g5538 = AND(g1669, g4313)
--	g4000 = AND(g1744, g2778)
--	g4126 = AND(g2701, g3040)
--	g4400 = AND(g4088, g3829)
--	g2794 = AND(I5886, I5887)
--	g4760 = AND(g486, g3393)
--	g6238 = AND(g572, g5096)
--	g10784 = AND(g10727, g5169)
--	g8174 = AND(g5284, g7853)
--	g6332 = AND(g1374, g5904)
--	g5067 = AND(g305, g4811)
--	g5418 = AND(g1512, g4344)
--	g10297 = AND(g8892, g10211)
--	g6353 = AND(g299, g5895)
--	g11026 = AND(g386, g10974)
--	g11212 = AND(g944, g11155)
--	g6744 = AND(g4828, g6151)
--	g5493 = AND(g1923, g4265)
--	g10671 = AND(g10578, g9431)
--	g4383 = AND(g2517, g3829)
--	g5256 = AND(g4297, g2779)
--	g4220 = AND(g105, g3539)
--	g8380 = AND(g8252, g4240)
--	g7071 = AND(g5916, g6590)
--	g4779 = AND(g501, g3427)
--	g9613 = AND(g1176, g9125)
--	g7705 = AND(g6853, g4328)
--	g9269 = AND(g8933, g3413)
--	g5181 = AND(g4520, g4510)
--	g4977 = AND(g4567, g4807)
--	g7948 = AND(g2855, g7497)
--	g11149 = AND(g324, g10930)
--	g9862 = AND(g1601, g9777)
--	g11387 = AND(g11284, g3629)
--	g7955 = AND(g2877, g7516)
--	g4161 = AND(g2719, g3060)
--	g11148 = AND(g2321, g10913)
--	g9712 = AND(g1528, g9490)
--	g8931 = AND(g8807, g8164)
--	g11097 = AND(g378, g10884)
--	g5421 = AND(g4631, g2733, g3819)
--	g11104 = AND(g2963, g10937)
--	g5263 = AND(g709, g4761)
--	g6092 = AND(g1059, g5320)
--	g4999 = AND(g1499, g4640)
--	I6338 = AND(g2475, g2456, g2451, g2446)
--	g7409 = AND(g4976, g632, g6858)
--	g4103 = AND(g2683, g2997)
--	I6309 = AND(g2446, g2451, g2456, g2475)
--	g6580 = AND(g1801, g5944)
--	g5631 = AND(g1056, g4416)
--	g9414 = AND(g1730, g9052)
--	g9660 = AND(g1188, g9125)
--	g9946 = AND(g9926, g9392)
--	g5257 = AND(g691, g4755)
--	g4732 = AND(g391, g3372)
--	g3108 = AND(I6330, I6331)
--	g4753 = AND(g481, g3386)
--	g9903 = AND(g9885, g9673)
--	g10625 = AND(g10546, g4552)
--	g5605 = AND(g4828, g704)
--	g6623 = AND(g55, g6170)
--	g11228 = AND(g466, g11060)
--	g11011 = AND(g1968, g10809)
--	g6889 = AND(g1941, g6427)
--	g8040 = AND(g7523, g5128)
--	g7822 = AND(g1914, g7479)
--	g8123 = AND(g1918, g7946)
--	g11582 = AND(g1311, g11540)
--	g4316 = AND(g1965, g3400)
--	g10969 = AND(g3625, g10809)
--	g5041 = AND(g3983, g4401)
--	g9335 = AND(g8975, g5708)
--	g9831 = AND(g9727, g9785)
--	g4565 = AND(g534, g4010)
--	g9422 = AND(g1750, g9030)
--	g8648 = AND(g4588, g8511)
--	g8875 = AND(g8255, g6368, g8858)
--	g5168 = AND(g1512, g4679)
--	g7895 = AND(g7503, g7036)
--	g8655 = AND(g8532, g4013)
--	g3396 = AND(g213, g3228)
--	g4914 = AND(g1062, g4436)
--	g9947 = AND(g9927, g9392)
--	g5772 = AND(g1555, g5214)
--	g6838 = AND(g192, g6596)
--	g5531 = AND(g1666, g4306)
--	g6795 = AND(g5036, g5878)
--	g10503 = AND(g10388, g2135)
--	g8010 = AND(g7738, g7413)
--	g8410 = AND(g713, g8143)
--	g6231 = AND(g818, g5608)
--	g10581 = AND(g10531, g9453)
--	g10450 = AND(g10364, g3359)
--	g2804 = AND(g2132, g1891)
--	g3418 = AND(g2379, g3012)
--	g4820 = AND(g186, g3946)
--	g9653 = AND(g1185, g9125)
--	g6205 = AND(g1515, g5151)
--	g10818 = AND(g10730, g4545)
--	g8172 = AND(g5275, g7853)
--	g10496 = AND(g10429, g3977)
--	g5074 = AND(g1771, g4587)
--	g9869 = AND(g1558, g9814)
--	g9719 = AND(g1543, g9490)
--	g10741 = AND(g10635, g4013)
--	g3381 = AND(g940, g2756)
--	g5863 = AND(g5272, g2173)
--	g8693 = AND(g3738, g8509)
--	g5480 = AND(g4279, g3519)
--	g4581 = AND(g3766, g3254)
--	g3685 = AND(g1781, g2981)
--	g5569 = AND(g4816, g2338)
--	g8555 = AND(g8409, g8025)
--	g3263 = AND(g2503, g2328)
--	g9364 = AND(g965, g9223)
--	g4784 = AND(g506, g3432)
--	g9454 = AND(g8994, g5708)
--	I6331 = AND(g2060, g2070, g2074, g2077)
--	g11299 = AND(g5498, g11243)
--	g6983 = AND(g6592, g3105)
--	g7958 = AND(g736, g7697)
--	g4995 = AND(g1474, g4640)
--	g4079 = AND(g2765, g2276)
--	g2264 = AND(g1771, g1766)
--	g2160 = AND(g745, g746)
--	g3257 = AND(g378, g2496)
--	g3101 = AND(I6309, I6310)
--	g5000 = AND(g1470, g4640)
--	g3301 = AND(g1346, g2544)
--	g5126 = AND(g3076, g4638)
--	I5084 = AND(g1462, g1470, g1474, g1478)
--	g9412 = AND(g1727, g9052)
--	g9389 = AND(g1330, g9151)
--	g2379 = AND(g744, g743)
--	g10706 = AND(g10567, g4840)
--	I16145 = AND(g10366, g10447, g10446)
--	g10597 = AND(g10533, g4359)
--	g8965 = AND(g8110, g6778, g8849)
--	g5608 = AND(g814, g4831)
--	g5220 = AND(g1083, g4729)
--	g10624 = AND(g10545, g4544)
--	g10300 = AND(g8892, g10220)
--	g5023 = AND(g1071, g4511)
--	g4432 = AND(g3723, g1975)
--	g4053 = AND(g2701, g2276)
--	g8050 = AND(g7596, g5919)
--	g5588 = AND(g1639, g4508)
--	g6679 = AND(g4631, g6074, g2733)
--	g9963 = AND(g9953, g9536)
--	g3772 = AND(g2542, g3089)
--	g5051 = AND(g4432, g2834)
--	g6831 = AND(g207, g6596)
--	g2981 = AND(g1776, g2264)
--	g8724 = AND(g8606, g7910)
--	g4157 = AND(g2713, g3055)
--	g9707 = AND(g1583, g9474)
--	g8878 = AND(g8099, g6368, g8858)
--	g2132 = AND(g1872, g1882)
--	g10763 = AND(g10639, g4840)
--	g8289 = AND(g6777, g8109, g6475)
--	g7898 = AND(g7511, g7041)
--	g11271 = AND(g5624, g11191)
--	g11461 = AND(g11429, g5446)
--	g5732 = AND(g1604, g5176)
--	g11145 = AND(g315, g10927)
--	g11031 = AND(g411, g10974)
--	g9865 = AND(g1607, g9780)
--	g5944 = AND(g1796, g5233)
--	g9715 = AND(g1531, g9490)
--	g9604 = AND(g1194, g9111)
--	g8799 = AND(g8647, g8727)
--	g11198 = AND(g4919, g11069)
--	g6873 = AND(g3263, g6557)
--	g6632 = AND(g61, g6190)
--	g6095 = AND(g1062, g5320)
--	g3863 = AND(g3323, g2728)
--	g9833 = AND(g9729, g9785)
--	g6653 = AND(g70, g6213)
--	g6102 = AND(g1038, g5320)
--	g7819 = AND(g1887, g7479)
--	g11393 = AND(g11280, g7916)
--	g2511 = AND(g461, g456)
--	g7088 = AND(g2331, g6737)
--	g9584 = AND(g2726, g9173)
--	g9896 = AND(g9883, g9624)
--	g8209 = AND(g4094, g3792, g7980)
--	g6752 = AND(g6187, g2343)
--	g4778 = AND(g421, g3426)
--	g11161 = AND(g1969, g10937)
--	g9268 = AND(g6681, g8947)
--	g5681 = AND(g135, g5361)
--	g7951 = AND(g2868, g7505)
--	g9419 = AND(g1744, g9030)
--	g10268 = AND(g10183, g3307)
--	g5533 = AND(g1724, g4308)
--	g9052 = AND(g8936, g7192)
--	g6786 = AND(g178, g5919)
--	g10670 = AND(g10571, g9091)
--	g11087 = AND(g829, g10950)
--	g4949 = AND(g3505, g4449)
--	g6364 = AND(g5851, g4454)
--	g7825 = AND(g1941, g7479)
--	g3400 = AND(g115, g3164)
--	g4998 = AND(g1304, g4485)
--	g10667 = AND(g10576, g9427)
--	g7136 = AND(g6050, g6704)
--	g6532 = AND(g339, g6057)
--	g9385 = AND(g1324, g9151)
--	I5690 = AND(g1436, g1440, g1444, g1448)
--	g4484 = AND(g1137, g3909)
--	g9897 = AND(g9884, g9624)
--	g9425 = AND(g1753, g9030)
--	g3383 = AND(g186, g3228)
--	g5601 = AND(g1035, g4375)
--	g7943 = AND(g2840, g7467)
--	g11171 = AND(g481, g11112)
--	g3423 = AND(I6630, I6631)
--	g7230 = AND(g6064, g6444)
--	g4952 = AND(g1648, g4457)
--	g8736 = AND(g7439, g8635)
--	g6787 = AND(g266, g5875)
--	g8968 = AND(g8089, g6778, g8849)
--	g10306 = AND(g10214, g9082)
--	g9331 = AND(g8972, g5708)
--	g11459 = AND(g11427, g5446)
--	g4561 = AND(g538, g4003)
--	g11425 = AND(g11350, g10899)
--	g11458 = AND(g11426, g5446)
--	g5739 = AND(g1607, g5185)
--	g7496 = AND(g7148, g2840)
--	g4986 = AND(g1411, g4682)
--	g11010 = AND(g5187, g10827)
--	g3999 = AND(g1741, g2777)
--	g8175 = AND(g5291, g7853)
--	g8722 = AND(g8604, g7908)
--	g4764 = AND(g411, g3404)
--	g7137 = AND(g5590, g6361)
--	g7891 = AND(g7471, g7028)
--	g8651 = AND(g8520, g4013)
--	g5479 = AND(g1845, g4243)
--	g11599 = AND(g1341, g11572)
--	g6684 = AND(g5314, g5836)
--	g6745 = AND(g5605, g6158)
--	g6639 = AND(g357, g6196)
--	g10937 = AND(g4822, g10822)
--	g3696 = AND(g1713, g3015)
--	g4503 = AND(g654, g3943)
--	g6791 = AND(g269, g5880)
--	g5190 = AND(g1245, g4716)
--	g5390 = AND(g3220, g4819)
--	g8384 = AND(g8180, g3397)
--	g4224 = AND(g1092, g3638)
--	g5501 = AND(g1672, g4273)
--	g9173 = AND(g8968, g6674)
--	g6759 = AND(g148, g5919)
--	g8838 = AND(g8602, g8702)
--	g8024 = AND(g7394, g4337)
--	g10666 = AND(g10575, g9424)
--	g11158 = AND(g309, g10935)
--	g9602 = AND(g2650, g9010)
--	g5704 = AND(g143, g5361)
--	g4617 = AND(g3275, g3879)
--	g11561 = AND(g11518, g3015)
--	g9868 = AND(g1555, g9812)
--	g11295 = AND(g5475, g11239)
--	g11144 = AND(g305, g10926)
--	g9718 = AND(g1540, g9490)
--	g3434 = AND(g237, g3228)
--	g4987 = AND(g1440, g4682)
--	g4771 = AND(g496, g3416)
--	g5250 = AND(g1270, g4748)
--	g6098 = AND(g1065, g5320)
--	g9582 = AND(g2725, g9173)
--	g6833 = AND(g186, g6596)
--	g3533 = AND(g1981, g2892)
--	g4892 = AND(g632, g4739)
--	g8104 = AND(g6218, g7880)
--	g9415 = AND(g1733, g9052)
--	g8499 = AND(g8377, g4737)
--	g9664 = AND(g1191, g9125)
--	g10740 = AND(g10676, g3384)
--	g2534 = AND(g798, g794)
--	g8754 = AND(g7420, g8667)
--	g9721 = AND(g9413, g4785)
--	g6162 = AND(g3584, g5200)
--	g4991 = AND(g1508, g4640)
--	g6362 = AND(g5846, g4450)
--	I6631 = AND(g2707, g2713, g2719, g2765)
--	g10685 = AND(g10608, g3863)
--	g4340 = AND(g1153, g3715)
--	g11023 = AND(g440, g10974)
--	g8044 = AND(g7598, g5919)
--	g11224 = AND(g968, g11056)
--	g11571 = AND(g2018, g11561)
--	g4959 = AND(g1520, g4682)
--	g10334 = AND(g10265, g3307)
--	g5626 = AND(g1633, g4557)
--	g9940 = AND(g9920, g9367)
--	g4876 = AND(g1086, g3638)
--	g6728 = AND(g6250, g4318)
--	g6730 = AND(g1872, g6128)
--	g9689 = AND(g263, g9432)
--	g10762 = AND(g10635, g4840)
--	g6070 = AND(g1050, g5320)
--	g9428 = AND(g1756, g9030)
--	g9030 = AND(g8935, g7192)
--	g9430 = AND(g1759, g9030)
--	g8927 = AND(g7872, g8807)
--	g7068 = AND(g5912, g6586)
--	g8014 = AND(g7740, g7419)
--	g11392 = AND(g11278, g7914)
--	g5782 = AND(g1558, g5223)
--	g9910 = AND(g9892, g9809)
--	g4824 = AND(g774, g4099)
--	g6331 = AND(g201, g5904)
--	g4236 = AND(g1098, g3638)
--	g11559 = AND(g2719, g11519)
--	g9609 = AND(g907, g9205)
--	g11558 = AND(g2713, g11519)
--	g6087 = AND(g1056, g5320)
--	g4877 = AND(g243, g3946)
--	g5526 = AND(g1950, g4294)
--	g10751 = AND(g10646, g4013)
--	g10772 = AND(g10655, g4840)
--	g8135 = AND(g1945, g7956)
--	g11544 = AND(g11515, g10584)
--	g5084 = AND(g1776, g4591)
--	g8382 = AND(g6077, g8213)
--	g10230 = AND(g8892, g10145)
--	g5484 = AND(g1896, g4256)
--	g7241 = AND(g6772, g6172)
--	g3942 = AND(g219, g3164)
--	g10638 = AND(g10608, g3829)
--	g4064 = AND(g1759, g2799)
--	g9365 = AND(g1321, g9151)
--	g9861 = AND(g9738, g9579)
--	g8749 = AND(g7604, g8660)
--	g11255 = AND(g456, g11075)
--	g11189 = AND(g5616, g11064)
--	g10510 = AND(g10393, g2135)
--	g8947 = AND(g8056, g6368, g8828)
--	g2917 = AND(g2424, g1657)
--	g5919 = AND(g5216, g2965)
--	g11188 = AND(g5604, g11063)
--	g9846 = AND(g287, g9764)
--	g7818 = AND(g1878, g7479)
--	g11460 = AND(g11428, g5446)
--	g5276 = AND(g736, g4780)
--	g11030 = AND(g406, g10974)
--	g11093 = AND(g841, g10950)
--	g7893 = AND(g7478, g7031)
--	g8653 = AND(g8526, g4013)
--	g10442 = AND(g10311, g2135)
--	g6535 = AND(g345, g6063)
--	g8102 = AND(g6209, g7878)
--	I5085 = AND(g1490, g1494, g1504, g1508)
--	g5004 = AND(g1296, g4499)
--	g3912 = AND(g207, g3164)
--	g7186 = AND(g2503, g6403)
--	g4489 = AND(g348, g3586)
--	g9662 = AND(g2094, g9292)
--	g9418 = AND(g1741, g9052)
--	g11218 = AND(g959, g11053)
--	g4471 = AND(g1121, g3862)
--	g10746 = AND(g10643, g4013)
--	g7125 = AND(g1212, g6648)
--	g7821 = AND(g1905, g7479)
--	g6246 = AND(g178, g5361)
--	g9256 = AND(g6689, g8963)
--	g8042 = AND(g7533, g5128)
--	g10237 = AND(g10145, g9100)
--	g7939 = AND(g2829, g7460)
--	g8786 = AND(g8638, g8716)
--	g10684 = AND(g10604, g3863)
--	g11455 = AND(g11435, g5446)
--	g8364 = AND(g658, g8235)
--	g2990 = AND(g2061, g2557, g1814)
--	g9847 = AND(g290, g9766)
--	g8054 = AND(g7584, g5919)
--	g5617 = AND(g1050, g4391)
--	g6502 = AND(g5981, g3095)
--	g5789 = AND(g1561, g5232)
--	g4009 = AND(g1747, g2789)
--	g11277 = AND(g4920, g11199)
--	g6940 = AND(g6472, g1945)
--	g7061 = AND(g790, g6760)
--	g11595 = AND(g1336, g11575)
--	g5771 = AND(g1534, g5213)
--	g8553 = AND(g8405, g8015)
--	g4836 = AND(g643, g3520)
--	g5547 = AND(g1733, g4326)
--	g6216 = AND(g2232, g5151)
--	g4967 = AND(g1515, g4682)
--	g6671 = AND(g342, g6227)
--	g7200 = AND(g3098, g6418)
--	g3661 = AND(g382, g3257)
--	g7046 = AND(g5892, g6570)
--	g4229 = AND(g999, g3914)
--	g8389 = AND(g6091, g8225)
--	g6430 = AND(g5044, g5791)
--	g8706 = AND(g7602, g8589)
--	g4993 = AND(g1448, g4682)
--	g6247 = AND(g127, g5361)
--	g9257 = AND(g6689, g8964)
--	g11170 = AND(g525, g11112)
--	g7145 = AND(g6082, g6718)
--	g5738 = AND(g1586, g5184)
--	g6826 = AND(g225, g6596)
--	g7191 = AND(g6343, g4323)
--	g3998 = AND(g2677, g2276)
--	g6741 = AND(g3284, g6141)
--	g5478 = AND(g1905, g4242)
--	g11167 = AND(g538, g11112)
--	g11194 = AND(g5637, g11067)
--	g11589 = AND(g1333, g11548)
--	g6638 = AND(g64, g6195)
--	g4921 = AND(g2779, g4431)
--	g7536 = AND(g7148, g2877)
--	g9585 = AND(g889, g8995)
--	g2957 = AND(g2424, g1663)
--	g11588 = AND(g1330, g11547)
--	g5690 = AND(g1567, g5112)
--	g6883 = AND(g1923, g6413)
--	g4837 = AND(g1068, g3638)
--	g8963 = AND(g8056, g6368, g8849)
--	g8791 = AND(g8641, g8721)
--	g6217 = AND(g563, g5073)
--	I6316 = AND(g2082, g2087, g2381, g2395)
--	g11022 = AND(g444, g10974)
--	g5915 = AND(g4168, g4977)
--	g4788 = AND(g511, g3436)
--	g8759 = AND(g7437, g8677)
--	g5110 = AND(g1806, g4618)
--	g11254 = AND(g986, g11073)
--	g6827 = AND(g219, g6596)
--	g8957 = AND(g8081, g6368, g8828)
--	g6333 = AND(g197, g5904)
--	g8049 = AND(g7567, g5919)
--	g4392 = AND(g3273, g3829)
--	g9856 = AND(g1592, g9773)
--	g9411 = AND(g1724, g9052)
--	g5002 = AND(g1494, g4640)
--	g11101 = AND(g857, g10950)
--	g11177 = AND(g511, g11112)
--	g11560 = AND(g2765, g11519)
--	g8098 = AND(g6201, g7852)
--	g3970 = AND(g225, g3164)
--	g4941 = AND(g1038, g4451)
--	g10453 = AND(g10437, g3395)
--	g5877 = AND(g4921, g639)
--	g6662 = AND(g366, g6220)
--	g7935 = AND(g2821, g7454)
--	g6067 = AND(g1047, g5320)
--	I6317 = AND(g2406, g2420, g2434, g2438)
--	g9863 = AND(g9740, g9576)
--	I5886 = AND(g174, g170, g2249, g2254)
--	g6994 = AND(g6758, g3829)
--	g9713 = AND(g1589, g9474)
--	g4431 = AND(g2268, g3533)
--	g4252 = AND(g1007, g3914)
--	g11166 = AND(g542, g11112)
--	g7130 = AND(g6041, g6697)
--	g11009 = AND(g5179, g10827)
--	g7542 = AND(g7148, g2885)
--	g8019 = AND(g7386, g4332)
--	g11008 = AND(g5171, g10827)
--	g3516 = AND(g1209, g3015)
--	g8052 = AND(g7573, g5128)
--	g3987 = AND(g243, g3164)
--	g4765 = AND(g491, g3405)
--	g11555 = AND(g2695, g11519)
--	g9857 = AND(g9734, g9569)
--	g8728 = AND(g8610, g7915)
--	g8730 = AND(g8613, g7917)
--	g8185 = AND(g664, g7997)
--	g5194 = AND(g1610, g4717)
--	g8385 = AND(g6084, g8218)
--	g4610 = AND(g3804, g2212)
--	g7902 = AND(g7661, g6587)
--	g4073 = AND(g3200, g3222)
--	g8070 = AND(g682, g7826)
--	g5731 = AND(g1583, g5175)
--	g11238 = AND(g5474, g11110)
--	g4473 = AND(g1125, g3874)
--	g8470 = AND(g8308, g7427)
--	g5489 = AND(g4287, g3521)
--	g3991 = AND(g1738, g2774)
--	I5887 = AND(g2078, g2083, g166, g2095)
--	g7823 = AND(g1923, g7479)
--	g4069 = AND(g1762, g2802)
--	g11519 = AND(g1317, g3015, g11492)
--	g11176 = AND(g506, g11112)
--	g11092 = AND(g837, g10950)
--	g11154 = AND(g330, g10932)
--	g9608 = AND(g7, g9292)
--	g11637 = AND(g11626, g5446)
--	g2091 = AND(g976, g971)
--	g8406 = AND(g695, g8131)
--	g5254 = AND(g4335, g4165)
--	g7260 = AND(g6752, g2345)
--	g5150 = AND(g1275, g4678)
--	g8766 = AND(g8612, g5151)
--	g9588 = AND(g3272, g9173)
--	g8801 = AND(g8742, g8729)
--	g7063 = AND(g5903, g6582)
--	g10303 = AND(g10208, g9076)
--	g5009 = AND(g1486, g4640)
--	g9665 = AND(g1314, g9151)
--	g8748 = AND(g7670, g8656)
--	g11215 = AND(g953, g11160)
--	g10750 = AND(g10687, g3586)
--	g5769 = AND(g2112, g4921, g3818)
--	g8755 = AND(g7426, g8671)
--	g6673 = AND(g5305, g5822)
--	g5212 = AND(g1255, g4726)
--	g7720 = AND(g727, g7232)
--	g5918 = AND(g2965, g5292, g4609)
--	g8045 = AND(g7547, g5128)
--	g8173 = AND(g7971, g3112)
--	g11349 = AND(g11288, g7964)
--	g7843 = AND(g7599, g5919)
--	g9696 = AND(g281, g9432)
--	g6772 = AND(g6228, g722)
--	g6058 = AND(g1035, g5320)
--	g6531 = AND(g79, g6056)
--	g6743 = AND(g4106, g6146)
--	g6890 = AND(g6752, g6568)
--	g7549 = AND(g7269, g3829)
--	g8169 = AND(g5265, g7853)
--	g11304 = AND(g5520, g11245)
--	g9944 = AND(g9924, g9392)
--	g9240 = AND(g6454, g8962)
--	g8059 = AND(g7592, g5919)
--	g8718 = AND(g8600, g7903)
--	g8767 = AND(g8616, g5151)
--	g9316 = AND(g8877, g5708)
--	g7625 = AND(g673, g7085)
--	g8793 = AND(g8644, g8723)
--	g2940 = AND(g2424, g1654)
--	g4114 = AND(g1351, g3301)
--	g11636 = AND(g11624, g7936)
--	g10949 = AND(g2947, g10809)
--	g4870 = AND(g237, g3946)
--	g3563 = AND(g3275, g2126)
--	g10948 = AND(g2223, g10809)
--	g8246 = AND(g7846, g7442)
--	g5788 = AND(g1540, g5231)
--	g4008 = AND(g2689, g2276)
--	g9596 = AND(g2649, g9010)
--	g5249 = AND(g1089, g4747)
--	g11585 = AND(g1321, g11543)
--	g3089 = AND(g2054, g2050)
--	g4972 = AND(g1436, g4682)
--	g11554 = AND(g2689, g11519)
--	g7586 = AND(g7096, g5423)
--	g10673 = AND(g10580, g9450)
--	g4806 = AND(g3215, g3992, g2493)
--	g5485 = AND(g1914, g4257)
--	g9936 = AND(g9915, g9624)
--	g2910 = AND(g2424, g1660)
--	g9317 = AND(g6109, g8875)
--	g10933 = AND(g10853, g3982)
--	g8388 = AND(g8177, g7689)
--	g4465 = AND(g1117, g3828)
--	g7141 = AND(g6073, g6716)
--	g10508 = AND(g10391, g2135)
--	g4230 = AND(g1095, g3638)
--	g10634 = AND(g10604, g3829)
--	g9601 = AND(g922, g9192)
--	g6126 = AND(g5639, g4319)
--	g6326 = AND(g1250, g5949)
--	g7710 = AND(g700, g7214)
--	g8028 = AND(g7375, g7436)
--	g6760 = AND(g786, g6221)
--	g5640 = AND(g1059, g4427)
--	g5031 = AND(g1478, g4640)
--	g4550 = AND(g342, g3586)
--	g7879 = AND(g7610, g3798)
--	g7962 = AND(g7730, g6712)
--	g9597 = AND(g1170, g9125)
--	g10452 = AND(g10439, g3388)
--	g4891 = AND(g631, g4739)
--	g5005 = AND(g1490, g4640)
--	g6423 = AND(g4348, g5784)
--	g8108 = AND(g1891, g7938)
--	g4807 = AND(g3015, g1289, g3937)
--	g5911 = AND(g3322, g4977)
--	g9937 = AND(g9916, g9624)
--	g9840 = AND(g9704, g9747)
--	g10780 = AND(g10723, g5124)
--	g8217 = AND(g1872, g7883)
--	g11013 = AND(g5209, g10827)
--	g9390 = AND(g1333, g9151)
--	g11214 = AND(g950, g11159)
--	g6327 = AND(g1255, g5949)
--	g4342 = AND(g1149, g3719)
--	g5796 = AND(g1564, g5252)
--	g5473 = AND(g4268, g3518)
--	g6346 = AND(g5038, g5883)
--	g6633 = AND(g354, g6191)
--	g11005 = AND(g5119, g10827)
--	g8365 = AND(g668, g8240)
--	g8048 = AND(g7558, g5919)
--	g4481 = AND(g1713, g3906)
--	g4097 = AND(g2677, g2989)
--	g8055 = AND(g7588, g5128)
--	g4497 = AND(g351, g3586)
--	g9942 = AND(g9922, g9367)
--	g6696 = AND(g5504, g5850)
--	g10731 = AND(g5118, g1850, g10665)
--	g8827 = AND(g8552, g8696)
--	g5540 = AND(g1727, g4315)
--	g4960 = AND(g1403, g4682)
--	g8846 = AND(g8615, g8712)
--	g6508 = AND(g5983, g3096)
--	g6240 = AND(g182, g5361)
--	g7931 = AND(g2809, g7446)
--	g5287 = AND(g3876, g4782)
--	g6472 = AND(g5853, g1936)
--	g11100 = AND(g853, g10950)
--	g11235 = AND(g5443, g11107)
--	g5199 = AND(g1068, g4719)
--	g6316 = AND(g1270, g5949)
--	g7515 = AND(g7148, g2855)
--	g10583 = AND(g10518, g10515)
--	g5781 = AND(g1537, g5222)
--	g8018 = AND(g7742, g7425)
--	g4401 = AND(g2971, g3772)
--	g8994 = AND(g8110, g6778, g8925)
--	g2950 = AND(g2424, g1666)
--	g5510 = AND(g1630, g4280)
--	g6347 = AND(g275, g5890)
--	g9357 = AND(g962, g9223)
--	g4828 = AND(g4106, g695)
--	g11407 = AND(g11339, g5949)
--	g4727 = AND(g386, g3364)
--	g10357 = AND(g10278, g2462)
--	g10743 = AND(g10639, g4013)
--	g5259 = AND(g627, g4739)
--	g5694 = AND(g162, g5361)
--	g10769 = AND(g10652, g4840)
--	g11584 = AND(g1318, g11542)
--	g4932 = AND(g1065, g4442)
--	g10768 = AND(g10649, g4840)
--	g6820 = AND(g1362, g6596)
--	g4068 = AND(g2719, g2276)
--	g6317 = AND(g1304, g5949)
--	g5215 = AND(g4276, g3400)
--	g4576 = AND(g530, g4049)
--	g4866 = AND(g231, g3946)
--	g6775 = AND(g822, g6231)
--	g3829 = AND(g2028, g2728)
--	g10662 = AND(g8892, g10571)
--	g8101 = AND(g6208, g7877)
--	g5825 = AND(g3204, g5318)
--	I6310 = AND(g2396, g2407, g2421, g2435)
--	g7884 = AND(g7457, g7022)
--	g5008 = AND(g1292, g4507)
--	g3974 = AND(g231, g3164)
--	g9949 = AND(g9929, g9392)
--	g2531 = AND(g658, g668)
--	g9292 = AND(g8878, g5708)
--	g10778 = AND(g1027, g10729)
--	g8041 = AND(g7524, g5128)
--	g6079 = AND(g1053, g5320)
--	g7235 = AND(g6663, g6447)
--	g9603 = AND(g1173, g9125)
--	g6840 = AND(g248, g6596)
--	g9850 = AND(g9726, g9560)
--	g7988 = AND(g1878, g7379)
--	g5228 = AND(g1086, g4734)
--	g7134 = AND(g5587, g6354)
--	g5934 = AND(g5215, g1965)
--	g5230 = AND(g1265, g4735)
--	g8168 = AND(g5262, g7853)
--	g9583 = AND(g886, g8995)
--	g10672 = AND(g10579, g9449)
--	g3287 = AND(g802, g2534)
--	g8772 = AND(g8627, g5151)
--	g4893 = AND(g635, g4739)
--	g10331 = AND(g10256, g3307)
--	g8505 = AND(g8309, g4789)
--	g10449 = AND(g10420, g3345)
--	g11273 = AND(g5638, g11195)
--	g8734 = AND(g8626, g7923)
--	g5913 = AND(g1041, g5320)
--	g10448 = AND(g10421, g3335)
--	g6163 = AND(g4572, g5354)
--	g6363 = AND(g284, g5901)
--	g7202 = AND(g6349, g4329)
--	g11463 = AND(g11432, g5446)
--	g8074 = AND(g718, g7826)
--	g4325 = AND(g1166, g3682)
--	g8474 = AND(g8383, g5285)
--	g11234 = AND(g5424, g11106)
--	g5266 = AND(g718, g4766)
--	g4483 = AND(g336, g3586)
--	g5248 = AND(g673, g4738)
--	g11514 = AND(g11491, g5151)
--	g5255 = AND(g682, g4754)
--	g4106 = AND(g3284, g686)
--	g2760 = AND(g981, g2091)
--	g5097 = AND(g1786, g4603)
--	g5726 = AND(g1601, g5167)
--	g5497 = AND(g4296, g3522)
--	g5354 = AND(g2733, g4460)
--	g7933 = AND(g2814, g7450)
--	g9617 = AND(g9, g9274)
--	g9906 = AND(g9873, g9683)
--	g11012 = AND(g5196, g10827)
--	g7050 = AND(g5896, g6575)
--	g10971 = AND(g10849, g3161)
--	g4904 = AND(g1850, g4243)
--	g10369 = AND(g10361, g3382)
--	g8400 = AND(g6097, g8234)
--	g4345 = AND(g1169, g3730)
--	g2161 = AND(I5084, I5085)
--	g5001 = AND(g1300, g4491)
--	g9945 = AND(g9925, g9392)
--	g7271 = AND(g5028, g6499)
--	g9709 = AND(g1524, g9490)
--	g4223 = AND(g1003, g3914)
--	g10716 = AND(g10497, g10675)
--	g11291 = AND(g11247, g4233)
--	g6661 = AND(g73, g6219)
--	g11173 = AND(g491, g11112)
--	g6075 = AND(g549, g5613)
--	g8023 = AND(g7367, g7430)
--	g9907 = AND(g9888, g9686)
--	g10582 = AND(g10532, g9473)
--	g5746 = AND(g1589, g5193)
--	g5221 = AND(g1260, g4730)
--	g9959 = AND(g9950, g9536)
--	g7674 = AND(g7004, g3880)
--	g9690 = AND(g266, g9432)
--	g6627 = AND(g58, g6181)
--	g5703 = AND(g174, g5361)
--	g4522 = AND(g360, g3586)
--	g4115 = AND(g2689, g3009)
--	g7541 = AND(g7075, g3109)
--	g10627 = AND(g10548, g4564)
--	g4047 = AND(g2695, g2276)
--	g6526 = AND(g76, g6052)
--	g2944 = AND(g2424, g1669)
--	g6646 = AND(g360, g6203)
--	g7132 = AND(g6048, g6702)
--	g11029 = AND(g401, g10974)
--	g8051 = AND(g7572, g5128)
--	g8127 = AND(g1927, g7949)
--	g7209 = AND(g3804, g6425)
--	g11028 = AND(g396, g10974)
--	g6439 = AND(g4479, g5919)
--	g10742 = AND(g10655, g3586)
--	g9110 = AND(g8880, g4790)
--	g10681 = AND(g10567, g3586)
--	g4537 = AND(g444, g3988)
--	g9663 = AND(g959, g9223)
--	g5349 = AND(g2126, g4617)
--	g8732 = AND(g8624, g7919)
--	g3807 = AND(g3003, g3062)
--	g8753 = AND(g7414, g8664)
--	g5848 = AND(g3860, g5519)
--	g8508 = AND(g8411, g7967)
--	g8072 = AND(g700, g7826)
--	g5699 = AND(g1592, g5117)
--	g11240 = AND(g5481, g11111)
--	g5398 = AND(g4610, g2224)
--	g6616 = AND(g6105, g3246)
--	g10690 = AND(g10616, g3863)
--	g8043 = AND(g7582, g5128)
--	g9590 = AND(g895, g8995)
--	g4128 = AND(g1976, g2779)
--	g6404 = AND(g2132, g5748)
--	g6647 = AND(g5288, g5808)
--	g10504 = AND(g10389, g2135)
--	g9657 = AND(g919, g9205)
--	g4542 = AND(g366, g3586)
--	g4330 = AND(g1163, g3693)
--	g3497 = AND(g2804, g1900)
--	g5524 = AND(g1678, g4291)
--	g8147 = AND(g2955, g7961)
--	g4554 = AND(g542, g3996)
--	g9899 = AND(g9889, g9367)
--	g5258 = AND(g700, g4756)
--	g7736 = AND(g6951, g3880)
--	g6224 = AND(g1520, g5151)
--	g10626 = AND(g10547, g4558)
--	g6320 = AND(g1292, g5949)
--	g7623 = AND(g664, g7079)
--	g10299 = AND(g8892, g10217)
--	g7889 = AND(g7615, g3814)
--	g10298 = AND(g8892, g10214)
--	g8413 = AND(g722, g8146)
--	g3979 = AND(g237, g3164)
--	g4902 = AND(g1848, g4243)
--	g5211 = AND(g1080, g4724)
--	g4512 = AND(g357, g3586)
--	g7722 = AND(g7127, g6449)
--	g9844 = AND(g9714, g9522)
--	g4490 = AND(g1141, g3913)
--	g4823 = AND(g207, g3946)
--	g6516 = AND(g5993, g3097)
--	g5026 = AND(g1453, g4640)
--	g8820 = AND(g8705, g5422)
--	g10737 = AND(g10687, g4840)
--	g8936 = AND(g8115, g6778, g8849)
--	g10232 = AND(g8892, g10150)
--	g6771 = AND(g263, g5866)
--	g5170 = AND(g1811, g4680)
--	g8117 = AND(g6236, g7886)
--	g4529 = AND(g448, g3980)
--	g4348 = AND(g3497, g1909)
--	g9966 = AND(g9956, g9536)
--	g5280 = AND(g4593, g3052)
--	g7139 = AND(g6060, g6709)
--	g11099 = AND(g382, g10885)
--	g6892 = AND(g6472, g5805)
--	g9705 = AND(g1580, g9474)
--	g10512 = AND(g10395, g2135)
--	g11098 = AND(g849, g10950)
--	g8775 = AND(g8628, g5151)
--	g5083 = AND(g3709, g4586)
--	g5544 = AND(g1687, g4320)
--	g11272 = AND(g5629, g11193)
--	g5483 = AND(g1621, g4254)
--	g9948 = AND(g9928, g9392)
--	g4063 = AND(g2713, g2276)
--	g11462 = AND(g11431, g5446)
--	g6738 = AND(g2531, g6137)
--	g8060 = AND(g7593, g5919)
--	g6244 = AND(g2255, g5151)
--	g11032 = AND(g416, g10974)
--	g10445 = AND(g10315, g2135)
--	g9150 = AND(g8882, g4805)
--	g10316 = AND(g10223, g9097)
--	g5756 = AND(g1531, g5202)
--	g4720 = AND(g1023, g3914)
--	g9409 = AND(g1721, g9052)
--	g8995 = AND(g6454, g8929)
--	g6876 = AND(g4070, g6560)
--	g4989 = AND(g1424, g4682)
--	g9836 = AND(g9737, g9785)
--	g6656 = AND(g2733, g6061, g4631)
--	g5514 = AND(g1941, g4284)
--	g8390 = AND(g8268, g6465)
--	g5003 = AND(g1466, g4640)
--	g9967 = AND(g9957, g9536)
--	g5145 = AND(g1639, g4673)
--	g4834 = AND(g219, g3946)
--	g4971 = AND(g1419, g4682)
--	g10753 = AND(g10649, g4013)
--	g5695 = AND(g166, g5361)
--	g7613 = AND(g6940, g5984)
--	g10736 = AND(g10658, g4840)
--	g11220 = AND(g962, g11054)
--	g7444 = AND(g7277, g5827)
--	g5536 = AND(g4867, g4298)
--	g6663 = AND(g6064, g2237)
--	g4670 = AND(g192, g3946)
--	g6824 = AND(g1371, g6596)
--	g4253 = AND(g1074, g3638)
--	g8250 = AND(g2771, g7907)
--	g8163 = AND(g7960, g3737)
--	g10764 = AND(g10643, g4840)
--	g5757 = AND(g1552, g5203)
--	g10365 = AND(g10319, g2135)
--	g8032 = AND(g7385, g7438)
--	g11591 = AND(g2988, g11561)
--	g8053 = AND(g7583, g5919)
--	g11147 = AND(g321, g10929)
--	g5522 = AND(g1633, g4289)
--	g5115 = AND(g1394, g4572)
--	g9837 = AND(g9697, g9751)
--	g9620 = AND(g2653, g9240)
--	g11151 = AND(g327, g10931)
--	g11172 = AND(g486, g11112)
--	g7885 = AND(g7614, g3812)
--	g6064 = AND(g5398, g2230)
--	g8929 = AND(g8095, g6368, g8828)
--	g5595 = AND(g1621, g4524)
--	g5537 = AND(g4143, g4299)
--	g9842 = AND(g9708, g9516)
--	g4141 = AND(g2707, g3051)
--	g4341 = AND(g339, g3586)
--	g9192 = AND(g6454, g8955)
--	g7679 = AND(g1950, g6863)
--	g7378 = AND(g6990, g3880)
--	g5612 = AND(g1627, g4543)
--	g3939 = AND(g213, g3164)
--	g7135 = AND(g869, g6355)
--	g10970 = AND(g10852, g3390)
--	g11025 = AND(g426, g10974)
--	g9854 = AND(g9730, g9566)
--	g7182 = AND(g1878, g6720)
--	g9941 = AND(g9921, g9367)
--	g6194 = AND(g554, g5043)
--	g5128 = AND(g4474, g2733)
--	g4962 = AND(g1651, g4461)
--	g4358 = AND(g1209, g3747)
--	g8683 = AND(g4803, g8549)
--	g4506 = AND(g1113, g3944)
--	g6471 = AND(g5224, g6014)
--	g8778 = AND(g8688, g2317)
--	g11281 = AND(g4948, g11202)
--	g8735 = AND(g7600, g8632)
--	g11146 = AND(g318, g10928)
--	g3904 = AND(g2948, g2779)
--	g8075 = AND(g727, g7826)
--	g9829 = AND(g9723, g9785)
--	g8949 = AND(g8255, g6368, g8828)
--	g7632 = AND(g7184, g5574)
--	g11290 = AND(g11246, g4226)
--	g6350 = AND(g5837, g4435)
--	g10599 = AND(g10534, g4365)
--	g5902 = AND(g2555, g4977)
--	I6337 = AND(g201, g2421, g2407, g2396)
--	g2276 = AND(g1765, g1610)
--	g6438 = AND(g5853, g5797)
--	g5512 = AND(g1660, g4281)
--	g5090 = AND(g1781, g4592)
--	g7719 = AND(g718, g7227)
--	g2561 = AND(g742, g741)
--	g3695 = AND(g1712, g3015)
--	g8603 = AND(g3983, g8548)
--	g8039 = AND(g7587, g5128)
--	g9610 = AND(g925, g9192)
--	g3536 = AND(g2390, g3103)
--	g5529 = AND(g4129, g4288)
--	g5148 = AND(g3088, g4671)
--	g9124 = AND(g8881, g4802)
--	g9324 = AND(g8879, g5708)
--	g4559 = AND(g2034, g3829)
--	g10561 = AND(g10549, g4583)
--	g5698 = AND(g1571, g5116)
--	g11226 = AND(g461, g11057)
--	g10295 = AND(g8892, g10208)
--	g5260 = AND(g1092, g4758)
--	g10680 = AND(g10564, g3586)
--	g6822 = AND(g231, g6596)
--	g4905 = AND(g1853, g4243)
--	g11551 = AND(g11538, g4013)
--	g3047 = AND(g1227, g2306)
--	g9849 = AND(g293, g9768)
--	g5279 = AND(g1766, g4783)
--	g8404 = AND(g686, g8129)
--	g5720 = AND(g170, g5361)
--	g5318 = AND(g4401, g1857)
--	g8764 = AND(g7443, g8684)
--	g11376 = AND(g11318, g4277)
--	g11297 = AND(g5490, g11242)
--	g9898 = AND(g9887, g9367)
--	
--	g6895 = OR(g6776, g4875)
--	g7189 = OR(g6632, g6053)
--	g9510 = OR(g9125, g9111)
--	g7297 = OR(g7132, g6323)
--	g9088 = OR(g8927, g8381)
--	g9923 = OR(g9865, g9707)
--	g6485 = OR(g5848, g5067)
--	g8771 = OR(g5483, g8652)
--	g5813 = OR(g5617, g4869)
--	g7963 = OR(g7687, g7182)
--	g10643 = OR(g10624, g7736)
--	g9886 = OR(g9607, g9592, g9759)
--	g9951 = OR(g9902, g9899, g9803)
--	g11625 = OR(g6535, g11597)
--	g8945 = OR(g8801, g8710)
--	g10489 = OR(g4961, g10367)
--	g10559 = OR(g4141, g10512)
--	g10558 = OR(g4126, g10510)
--	g11338 = OR(g11283, g11178)
--	g8435 = OR(g8403, g8075)
--	g10544 = OR(g5511, g10495)
--	g6911 = OR(g6342, g5681)
--	g10865 = OR(g5538, g10752)
--	g3698 = OR(g3121, g2480)
--	g8214 = OR(g7472, g8004)
--	g6124 = OR(g5181, g5188)
--	g6469 = OR(g5698, g4959)
--	g5587 = OR(g4714, g3904)
--	g6177 = OR(g5444, g4712)
--	I14585 = OR(g8995, g9205, g9192)
--	g9891 = OR(g9741, g9760)
--	g9913 = OR(g9849, g9691)
--	I5600 = OR(g496, g491, g486, g481)
--	g11257 = OR(g11234, g11019)
--	g8236 = OR(g7526, g8001)
--	g7385 = OR(g7235, g6746)
--	g6898 = OR(g6790, g4881)
--	g6900 = OR(g6787, g6246)
--	g4264 = OR(g4048, g4053)
--	g9726 = OR(g9411, g9420, g9489)
--	g6088 = OR(g5260, g4522)
--	g6923 = OR(g6353, g5695)
--	g8194 = OR(g5168, g7940)
--	g9676 = OR(g9454, g9292, g9274)
--	g11256 = OR(g11186, g11018)
--	g3860 = OR(g3107, g2167)
--	g11280 = OR(g11254, g11153)
--	g9727 = OR(g9650, g9663, g9362, I14866)
--	g4997 = OR(g4581, g4584)
--	g11624 = OR(g11595, g11571)
--	g11300 = OR(g11213, g11091)
--	g4238 = OR(g3999, g4007)
--	g8814 = OR(g7945, g8728)
--	g10401 = OR(g9317, g10291)
--	g8773 = OR(g5491, g8653)
--	g11231 = OR(g11156, g11013)
--	g10864 = OR(g5532, g10751)
--	g9624 = OR(g9316, g9313)
--	g9953 = OR(g9945, g9939, g9669)
--	g6122 = OR(g5172, g5180)
--	g6465 = OR(g5825, g5041)
--	g6934 = OR(g6363, g5720)
--	g7664 = OR(g6855, g4084)
--	g7246 = OR(g6465, g6003)
--	g7203 = OR(g6640, g6058)
--	g6096 = OR(g5268, g4542)
--	g9747 = OR(g9173, g9509)
--	g11314 = OR(g11224, g11102)
--	g10733 = OR(g5227, g10674)
--	g8921 = OR(g8827, g8748)
--	I15054 = OR(g7853, g9782, g9624, g9785)
--	g11269 = OR(g11196, g11031)
--	g5555 = OR(g4389, g4397)
--	g11268 = OR(g11194, g11030)
--	g10485 = OR(g9317, g10376)
--	g10555 = OR(g4103, g10504)
--	g6481 = OR(g5722, g4972)
--	g10712 = OR(g10662, g9531)
--	g11335 = OR(g11279, g11175)
--	g8249 = OR(g8018, g7710)
--	g7638 = OR(g7265, g6488)
--	g10567 = OR(g10514, g7378)
--	g11487 = OR(g6662, g11464)
--	I15210 = OR(g9839, g9964, g9852, g9882)
--	I5805 = OR(g2102, g2099, g2096, g2088)
--	g8941 = OR(g8796, g8706)
--	g11443 = OR(g7130, g11407)
--	g4231 = OR(g3991, g3998)
--	g11278 = OR(g11253, g11150)
--	I15039 = OR(g7853, g9809, g9624, g9785)
--	g11286 = OR(g10670, g11209)
--	g8431 = OR(g8387, g8071)
--	g7133 = OR(g6616, g3067)
--	g11306 = OR(g11216, g11095)
--	g8252 = OR(g7988, g7679)
--	g8812 = OR(g7939, g8724)
--	g7846 = OR(g7722, g7241)
--	g3875 = OR(g3275, g12)
--	g5996 = OR(g5473, g3908)
--	g6592 = OR(g5100, g5882)
--	g8286 = OR(g8107, g7823)
--	g10501 = OR(g4161, g10445)
--	g10728 = OR(g4973, g10642)
--	g8270 = OR(g7894, g3434)
--	g7290 = OR(g7046, g6316)
--	g6068 = OR(g5220, g4497)
--	g6468 = OR(g5690, g4950)
--	g11217 = OR(g11144, g11005)
--	g11478 = OR(g6532, g11455)
--	g9536 = OR(g9335, g9331, g9328, g9324)
--	g5981 = OR(g5074, g4383)
--	g11486 = OR(g6654, g11463)
--	g8377 = OR(g8185, g7958)
--	g8206 = OR(g7459, g8007)
--	g11580 = OR(g11413, g11544)
--	g8287 = OR(g8117, g7824)
--	g11223 = OR(g11147, g11008)
--	g9522 = OR(g9173, g9125)
--	g8199 = OR(g7902, g7444)
--	g5802 = OR(g5601, g4837)
--	g11321 = OR(g11230, g11105)
--	g6524 = OR(g5746, g4996)
--	g10664 = OR(g10240, g10582)
--	g7257 = OR(g6701, g4725)
--	g7301 = OR(g7140, g6327)
--	g10484 = OR(g9317, g10400)
--	g10554 = OR(g4097, g10503)
--	g8259 = OR(g8028, g7719)
--	g11334 = OR(g11277, g11174)
--	g8819 = OR(g7957, g8734)
--	g8923 = OR(g8846, g8763)
--	g8488 = OR(g3664, g8390)
--	g7441 = OR(g7271, g6789)
--	g6026 = OR(g5507, g3970)
--	g10799 = OR(g6225, g10769)
--	g10798 = OR(g6217, g10768)
--	g10805 = OR(g10759, g10760)
--	g10732 = OR(g4358, g10661)
--	g6061 = OR(g5204, g4)
--	g9512 = OR(g9151, g9125)
--	g10013 = OR(I15214, I15215)
--	g8806 = OR(g7931, g8718)
--	g8943 = OR(g8837, g8749)
--	g11293 = OR(g11211, g10818)
--	g11265 = OR(g11189, g11027)
--	g8887 = OR(g8842, g8755)
--	g5838 = OR(g5612, g4866)
--	g6514 = OR(g5738, g4992)
--	g8322 = OR(g8136, g6891)
--	g8230 = OR(g7515, g7991)
--	g5809 = OR(g5611, g4865)
--	g8433 = OR(g8399, g8073)
--	g11579 = OR(g5123, g11551)
--	g10771 = OR(g5533, g10684)
--	g11615 = OR(g11601, g11592)
--	g9367 = OR(g9335, g9331)
--	g9872 = OR(g9617, g9594, g9750)
--	g6522 = OR(g5744, g4994)
--	g8266 = OR(g7885, g3412)
--	g10414 = OR(g10300, g9534)
--	g11275 = OR(g11248, g11148)
--	g11430 = OR(g11387, g4006)
--	g8248 = OR(g8014, g7707)
--	g9686 = OR(g9454, g9292, g9274)
--	g8815 = OR(g7948, g8730)
--	g7183 = OR(g6623, g6046)
--	g5983 = OR(g5084, g4392)
--	g8154 = OR(g7891, g6879)
--	g6537 = OR(g5781, g5005)
--	g4309 = OR(g4069, g4079)
--	g10725 = OR(g4962, g10634)
--	g6243 = OR(g5537, g4774)
--	I6351 = OR(g2405, g2389, g2380, g2372)
--	g9519 = OR(g9173, g9151, g9125)
--	g9740 = OR(g9418, g9505)
--	g8267 = OR(g7889, g3422)
--	g10744 = OR(g10600, g10668, I16427)
--	g6542 = OR(g5789, g5010)
--	g7303 = OR(g7145, g6329)
--	g10652 = OR(g10627, g7743)
--	g5036 = OR(g4871, g4162)
--	g7240 = OR(g6687, g6095)
--	g8221 = OR(g7496, g7993)
--	g6902 = OR(g6794, g4223)
--	I14776 = OR(g8995, g9205, g9192)
--	g10500 = OR(g4157, g10442)
--	g4052 = OR(g2862, g2515)
--	I14858 = OR(g9585, g9595, g9610, g9602)
--	g6529 = OR(g5757, g5000)
--	g11264 = OR(g11188, g11026)
--	I15209 = OR(g8169, g9905, g9934, g9830)
--	g8241 = OR(g7536, g7989)
--	g10795 = OR(g6199, g10764)
--	g11607 = OR(g11586, g11557)
--	g8644 = OR(g8123, g8464)
--	g4682 = OR(g3563, g3348, g1570)
--	g8818 = OR(g7955, g8733)
--	g2984 = OR(g2528, g2522)
--	g9931 = OR(g8931, g9900)
--	g3414 = OR(g2911, g2917)
--	g9515 = OR(g9173, g9151)
--	g10724 = OR(g10312, g10672)
--	g7294 = OR(g7068, g6320)
--	g5189 = OR(g4345, g3496)
--	g8614 = OR(g8365, g8510)
--	g3513 = OR(g3118, g2180)
--	g6909 = OR(g6346, g5684)
--	I5571 = OR(g396, g391, g386, g426)
--	g4283 = OR(g4059, g4063)
--	g8939 = OR(g8791, g8701)
--	g2514 = OR(I5599, I5600)
--	g11327 = OR(g11297, g11167)
--	g8187 = OR(g7542, g7998)
--	g11606 = OR(g11585, g11556)
--	g11303 = OR(g11214, g11092)
--	g5309 = OR(g3664, g4401)
--	g9528 = OR(g9151, g9125, g9111)
--	g8200 = OR(g7535, g8008)
--	g2522 = OR(g833, g829, I5629)
--	g2315 = OR(g1163, g1166, g1113, I5363)
--	g6506 = OR(g5731, g4989)
--	g10649 = OR(g10626, g7741)
--	g8159 = OR(g7895, g6886)
--	g7626 = OR(g7060, g5267)
--	g10770 = OR(g5525, g10682)
--	g9566 = OR(g9052, g9030)
--	g11483 = OR(g6633, g11460)
--	g8811 = OR(g7935, g8722)
--	g8642 = OR(g5236, g5205, g8465)
--	g6545 = OR(g5795, g5025)
--	g10767 = OR(g5500, g10681)
--	g11326 = OR(g11296, g11166)
--	g10898 = OR(g4220, g10777)
--	g11252 = OR(g11099, g10969)
--	g10719 = OR(g10303, g10666)
--	g4609 = OR(g3400, g119)
--	g6507 = OR(g5732, g4990)
--	g10718 = OR(g6238, g10706)
--	g10521 = OR(I16148, I16149)
--	g7075 = OR(g5104, g6530)
--	g7292 = OR(g7055, g6318)
--	g10861 = OR(g5523, g10745)
--	g8417 = OR(g8246, g7721)
--	g6515 = OR(g5739, g4993)
--	I14855 = OR(g9583, g9593, g9601, g9596)
--	I15205 = OR(g9838, g9963, g9850, g9878)
--	I15051 = OR(g7853, g9673, g9624, g9785)
--	g9724 = OR(g9409, g9419, g9615)
--	g6528 = OR(g5756, g4999)
--	g8823 = OR(g8778, g8693)
--	g7503 = OR(g6887, g6430)
--	g8148 = OR(g7884, g6872)
--	g8649 = OR(g8499, g4519)
--	g3584 = OR(g2863, g2516)
--	g10776 = OR(g5544, g10758)
--	g9680 = OR(g9454, g9292, g9274)
--	g10859 = OR(g5512, g10742)
--	I14866 = OR(g9590, g9609, g9619)
--	g7299 = OR(g7138, g6325)
--	g10858 = OR(g5501, g10741)
--	g8193 = OR(g5145, g7937)
--	g9511 = OR(g9151, g9125, g9111)
--	g7738 = OR(g7200, g6738)
--	g7244 = OR(g6699, g4720)
--	g3425 = OR(g2895, g2910)
--	g7478 = OR(g6884, g6423)
--	g9714 = OR(g9664, g9366, g9654)
--	g10025 = OR(I15224, I15225)
--	g6908 = OR(g6345, g4229)
--	g5028 = OR(g4836, g4128)
--	g8253 = OR(g8023, g7718)
--	g8938 = OR(g8789, g8699)
--	g8813 = OR(g7943, g8726)
--	g9736 = OR(g9430, g9416)
--	g9968 = OR(I15171, I15172)
--	g8552 = OR(g8217, g8388)
--	g5910 = OR(g5023, g4341)
--	g11249 = OR(g6162, g11143)
--	g11482 = OR(g6628, g11459)
--	g9722 = OR(g9612, g9643, g9410, I14855)
--	I15204 = OR(g8168, g9904, g9933, g9829)
--	g7236 = OR(g6684, g6092)
--	I14596 = OR(g8995, g9205, g9192)
--	g8645 = OR(g8127, g8469)
--	g11647 = OR(g6622, g11637)
--	g6777 = OR(g5691, g5052)
--	g9737 = OR(g9657, g9658, g9655)
--	I16149 = OR(g10472, g10470, g10468, g10467)
--	g11233 = OR(g11085, g10946)
--	g8607 = OR(g8406, g8554)
--	I16148 = OR(g10386, g10384, g10476, g10474)
--	g8158 = OR(g7893, g6883)
--	g5846 = OR(g4932, g4236)
--	g5396 = OR(g4481, g3684)
--	g5803 = OR(g5575, g4820)
--	g11331 = OR(g11272, g11171)
--	g7295 = OR(g7071, g6321)
--	g6541 = OR(g5788, g5009)
--	g8615 = OR(g8413, g8557)
--	g9742 = OR(g9173, g9528)
--	g9926 = OR(g9868, g9715)
--	g9754 = OR(g9173, g9511)
--	g8284 = OR(g8102, g7821)
--	g2204 = OR(g1393, g1394)
--	g7471 = OR(g6880, g6416)
--	g7242 = OR(g6693, g6098)
--	g5847 = OR(g5626, g4877)
--	g6901 = OR(g6788, g6247)
--	g8559 = OR(g8380, g4731)
--	g9729 = OR(g9618, g9357, g9656)
--	g10860 = OR(g5513, g10743)
--	g9927 = OR(g9869, g9716)
--	g10497 = OR(g5052, g10396)
--	g9885 = OR(g9739, g9598, g9662, g9746)
--	g2528 = OR(g861, g857, g853, g849)
--	g11229 = OR(g11154, g11012)
--	g8973 = OR(g8821, g8735)
--	g10658 = OR(g10595, g7674)
--	g10339 = OR(g10232, g9556)
--	I5363 = OR(g1149, g1153, g1157, g1160)
--	g11310 = OR(g11220, g11100)
--	g6500 = OR(g5725, g4986)
--	g10855 = OR(g6075, g10736)
--	g9916 = OR(g9855, g9694)
--	g10411 = OR(g10299, g9529)
--	g11603 = OR(g11582, g11553)
--	I5357 = OR(g1265, g1260, g1255, g1250)
--	g9560 = OR(g9052, g9030)
--	g6672 = OR(g5941, g5259)
--	g9873 = OR(g9623, g9599, g9758)
--	g6523 = OR(g5745, g4995)
--	g10707 = OR(g5545, g10686)
--	I5626 = OR(g521, g525, g530, g534)
--	g9579 = OR(g9052, g9030)
--	g7298 = OR(g7136, g6324)
--	g6551 = OR(g5804, g5031)
--	g6099 = OR(g5273, g4550)
--	g8282 = OR(g8101, g7819)
--	g9917 = OR(g9856, g9695)
--	I15057 = OR(g7853, g9680, g9624, g9785)
--	g7219 = OR(g6661, g6076)
--	g10019 = OR(I15219, I15220)
--	g5857 = OR(g5418, g4670)
--	g9725 = OR(g9642, g9659, g9616, I14862)
--	g11298 = OR(g11212, g11087)
--	g10402 = OR(g10295, g9554)
--	g2521 = OR(g538, g542, g476, I5626)
--	I14751 = OR(g8995, g9205, g9192)
--	g10866 = OR(g5539, g10753)
--	g6534 = OR(g5772, g5003)
--	g11232 = OR(g11158, g11015)
--	g9706 = OR(g9644, g9386, g9591)
--	g10001 = OR(I15204, I15205)
--	g8776 = OR(g5510, g8655)
--	g7225 = OR(g6666, g6079)
--	g9888 = OR(g9648, g9608, g9757)
--	g11261 = OR(g11238, g11023)
--	g9956 = OR(g9948, g9942, g9815)
--	g10923 = OR(g10778, g10715)
--	g8264 = OR(g7879, g3389)
--	g6513 = OR(g5737, g4991)
--	I14835 = OR(g9621, g9645, g9588)
--	g8641 = OR(g8120, g8463)
--	g5361 = OR(g4316, g4093, g126)
--	g11316 = OR(g11226, g11103)
--	I16161 = OR(g10479, g10478, g10477, g10475)
--	g6916 = OR(g6348, g5687)
--	g8777 = OR(g5522, g8659)
--	g2353 = OR(g1403, g1407, g1411, g1415)
--	g7510 = OR(g7186, g6730)
--	g9957 = OR(g9949, g9943, g9776)
--	g2744 = OR(I5804, I5805)
--	g7245 = OR(g6696, g6102)
--	g7291 = OR(g7050, g6317)
--	g8611 = OR(g8410, g8556)
--	I15199 = OR(g8167, g9903, g9932, g9828)
--	g10550 = OR(g4942, g10450)
--	g11330 = OR(g11304, g11170)
--	g10721 = OR(g10306, g10669)
--	g8153 = OR(g7888, g6875)
--	g10773 = OR(g5540, g10685)
--	g3688 = OR(g3144, g2454)
--	I15225 = OR(g9842, g9967, g9859, g9881)
--	g6042 = OR(g5535, g3987)
--	g10655 = OR(g10561, g7389)
--	g11259 = OR(g11236, g11021)
--	g11225 = OR(g11149, g11009)
--	g5914 = OR(g5029, g4343)
--	g11258 = OR(g11235, g11020)
--	g6054 = OR(g5199, g4483)
--	g9728 = OR(g9412, g9422, g9426)
--	g9730 = OR(g9414, g9425, g9423)
--	g5820 = OR(g5595, g4834)
--	g8574 = OR(g5679, g7853, g8465)
--	g11602 = OR(g11581, g11552)
--	g10502 = OR(g4169, g10365)
--	g10557 = OR(g4123, g10508)
--	I15171 = OR(g8175, g9909, g9896, g9835)
--	g11337 = OR(g11282, g11177)
--	g7465 = OR(g6876, g6410)
--	g8262 = OR(g7970, g7625)
--	g8889 = OR(g8844, g8756)
--	g7096 = OR(g6544, g5911)
--	g5995 = OR(g5097, g5099)
--	g8285 = OR(g8104, g7822)
--	g10791 = OR(g6186, g10762)
--	g2499 = OR(I5570, I5571)
--	I14607 = OR(g8995, g9205, g9192)
--	g6049 = OR(g5254, g3718)
--	g9920 = OR(g9860, g9701)
--	g10556 = OR(g4115, g10506)
--	g8643 = OR(g8364, g8508)
--	g5810 = OR(g5588, g4823)
--	g11336 = OR(g11281, g11176)
--	g8742 = OR(g8135, g8598)
--	g8926 = OR(g8848, g8764)
--	g7218 = OR(g6655, g6070)
--	I15224 = OR(g8174, g9908, g9937, g9834)
--	g7293 = OR(g7063, g6319)
--	g11288 = OR(g11204, g11070)
--	g10800 = OR(g6245, g10772)
--	g11308 = OR(g11218, g11098)
--	g8269 = OR(g7892, g3429)
--	g10417 = OR(g10301, g9527)
--	g10936 = OR(g5170, g10808)
--	g9388 = OR(g9240, g9223)
--	g6185 = OR(g5470, g4715)
--	g6470 = OR(g5699, g4960)
--	g6897 = OR(g6771, g6240)
--	g8885 = OR(g8841, g8754)
--	g11260 = OR(g11237, g11022)
--	g11488 = OR(g6671, g11465)
--	g6105 = OR(g5279, g4559)
--	g10807 = OR(g10701, g10761)
--	g10639 = OR(g10623, g7734)
--	g4556 = OR(g3536, g2916)
--	g8288 = OR(g8119, g7825)
--	g6755 = OR(g6106, g5479)
--	I14862 = OR(g9587, g9600, g9611)
--	I16160 = OR(g10394, g10392, g10482, g10481)
--	I15042 = OR(g7853, g9686, g9624, g9785)
--	g11610 = OR(g11589, g11560)
--	g9711 = OR(g9660, g9390, g9359, g9589)
--	g6045 = OR(g5541, g3989)
--	g11270 = OR(g11198, g11032)
--	g7258 = OR(g6549, g5913)
--	g6059 = OR(g5211, g4489)
--	g10007 = OR(I15209, I15210)
--	g11267 = OR(g11192, g11029)
--	g11294 = OR(g6576, g11210)
--	g9509 = OR(g9151, g9125, g9111)
--	g7211 = OR(g6647, g6067)
--	g5404 = OR(g4487, g3696)
--	g4089 = OR(g1959, g3318)
--	I15219 = OR(g8172, g9907, g9936, g9833)
--	g11219 = OR(g11145, g11006)
--	g6015 = OR(g5497, g3942)
--	g10720 = OR(g10304, g10667)
--	g8265 = OR(g7881, g3396)
--	g5224 = OR(g4360, g3512)
--	g9700 = OR(g9358, g9667, I14827)
--	g7106 = OR(g6554, g5917)
--	g8770 = OR(g5476, g8651)
--	g11201 = OR(g11152, g11011)
--	g9950 = OR(g9901, g9898, g9779)
--	g9723 = OR(g9620, g9652, g9391, I14858)
--	g2309 = OR(I5357, I5358)
--	g11266 = OR(g11190, g11028)
--	g10727 = OR(g4969, g10638)
--	g10863 = OR(g5531, g10750)
--	g8429 = OR(g8385, g8069)
--	g9751 = OR(g9515, g9510)
--	g8281 = OR(g8097, g7818)
--	g6910 = OR(g6341, g5680)
--	g8639 = OR(g8118, g8462)
--	g9673 = OR(g9454, g9292, g9274)
--	g11285 = OR(g11255, g11161)
--	g11305 = OR(g11215, g11093)
--	I15177 = OR(g9844, g9960, g9863, g9876)
--	g9734 = OR(g9415, g9428, g9421)
--	I14827 = OR(g9603, g9614, g9584)
--	g5824 = OR(g5602, g4839)
--	g8715 = OR(g8416, g8687)
--	g5762 = OR(g5178, g5186)
--	g6538 = OR(g5782, g5006)
--	g5590 = OR(g4718, g4723)
--	g10726 = OR(g10316, g10673)
--	g3120 = OR(I6350, I6351)
--	g9573 = OR(g9052, g9030)
--	g4640 = OR(g3348, g3563, g1527)
--	g6093 = OR(g5264, g4534)
--	g8162 = OR(g7898, g6889)
--	g8268 = OR(g7962, g7613)
--	g9569 = OR(g9052, g9030)
--	g11485 = OR(g6646, g11462)
--	g10797 = OR(g6206, g10766)
--	I14779 = OR(g8995, g9205, g9192)
--	g10408 = OR(g10298, g9553)
--	g10635 = OR(g10622, g7732)
--	g2305 = OR(I5351, I5352)
--	I15176 = OR(g8176, g9910, g9897, g9836)
--	g3435 = OR(g2945, g2950)
--	g9924 = OR(g9866, g9709)
--	g10711 = OR(g5547, g10690)
--	g5814 = OR(g5591, g4827)
--	g5038 = OR(g4878, g4884)
--	I15215 = OR(g9840, g9965, g9854, g9879)
--	g8226 = OR(g7504, g8002)
--	g7367 = OR(g7224, g6744)
--	g7457 = OR(g6873, g6404)
--	g5229 = OR(g4364, g3516)
--	g5993 = OR(g5090, g4400)
--	g8283 = OR(g8098, g7820)
--	g7971 = OR(g5110, g7549)
--	g8602 = OR(g8401, g8550)
--	g8920 = OR(g8845, g8759)
--	g10663 = OR(g10237, g10581)
--	g6074 = OR(g5349, g1)
--	g8261 = OR(g7876, g3383)
--	g10862 = OR(g5524, g10746)
--	g5837 = OR(g5640, g4224)
--	g11333 = OR(g11274, g11173)
--	g6080 = OR(g5249, g4512)
--	g6480 = OR(g5721, g4971)
--	g7740 = OR(g7209, g6741)
--	g10702 = OR(g10562, g3877)
--	g9697 = OR(g9665, g9606, I14822)
--	g8203 = OR(g7453, g7999)
--	g9914 = OR(g9851, g9692)
--	g10564 = OR(g10560, g7368)
--	g11484 = OR(g6639, g11461)
--	g5842 = OR(g5618, g4870)
--	I15200 = OR(g9837, g9962, g9848, g9880)
--	g11609 = OR(g11588, g11559)
--	I14582 = OR(g8995, g9205, g9192)
--	g8940 = OR(g8793, g8703)
--	g11312 = OR(g11222, g11101)
--	g11608 = OR(g11587, g11558)
--	g6000 = OR(g5480, g3912)
--	g8428 = OR(g8382, g8068)
--	g8430 = OR(g8386, g8070)
--	g9922 = OR(g9864, g9705)
--	g8247 = OR(g8010, g7704)
--	g3438 = OR(g2939, g2944)
--	I5576 = OR(g431, g435, g440, g444)
--	g6924 = OR(g6362, g4261)
--	g5405 = OR(g4476, g3440)
--	g8638 = OR(g8108, g8461)
--	g8609 = OR(g8408, g8555)
--	g9995 = OR(I15199, I15200)
--	g8883 = OR(g8838, g8753)
--	I15214 = OR(g8170, g9906, g9935, g9831)
--	g2538 = OR(g1466, g1458, I5649)
--	g11329 = OR(g11302, g11169)
--	g4255 = OR(g4009, g4047)
--	g11328 = OR(g11299, g11168)
--	g9704 = OR(g9385, g9605, I14835)
--	I5352 = OR(g1129, g1125, g1121, g1117)
--	g8774 = OR(g5499, g8654)
--	g9954 = OR(g9946, g9940, g9781)
--	g10405 = OR(g10297, g9530)
--	g9363 = OR(g9205, g9192)
--	g5849 = OR(g4949, g4260)
--	I5599 = OR(g516, g511, g506, g501)
--	g7204 = OR(g6645, g6062)
--	g7300 = OR(g7139, g6326)
--	g4293 = OR(g4064, g4068)
--	g9912 = OR(g9847, g9690)
--	g6533 = OR(g5771, g5002)
--	g8816 = OR(g7951, g8731)
--	g9929 = OR(g9871, g9718)
--	g5819 = OR(g5625, g4876)
--	I14831 = OR(g9613, g9622, g9586)
--	g5852 = OR(g5632, g4883)
--	g8263 = OR(g8032, g7720)
--	g3431 = OR(g2951, g2957)
--	g9683 = OR(g9454, g9292, g9274)
--	g8631 = OR(g8474, g7449)
--	g6922 = OR(g6352, g5694)
--	g8817 = OR(g7954, g8732)
--	g9735 = OR(g9649, g9651, g9384, g9361)
--	g8605 = OR(g8404, g8553)
--	g11263 = OR(g11187, g11025)
--	g6739 = OR(g5769, g5780)
--	g11332 = OR(g11273, g11172)
--	g7143 = OR(g6619, g6039)
--	g6479 = OR(g5707, g4968)
--	I15048 = OR(g7853, g9683, g9624, g9785)
--	g6501 = OR(g5726, g4987)
--	g9702 = OR(g9365, g9647, I14831)
--	g11221 = OR(g11146, g11007)
--	g9952 = OR(g9944, g9938, g9817)
--	g11613 = OR(g11600, g11591)
--	g7621 = OR(g5108, g6994)
--	g3399 = OR(g2918, g2940)
--	g11605 = OR(g11584, g11555)
--	g4274 = OR(g4054, g4058)
--	I14602 = OR(g8995, g9205, g9192)
--	I15033 = OR(g7853, g9804, g9624, g9785)
--	g10717 = OR(g6235, g10705)
--	I5629 = OR(g845, g841, g837)
--	g9925 = OR(g9867, g9712)
--	g3819 = OR(g3275, g9)
--	g6912 = OR(g6350, g4235)
--	g10723 = OR(g4952, g10633)
--	g6929 = OR(g6360, g5704)
--	g10646 = OR(g10625, g7739)
--	g9516 = OR(g9151, g9125)
--	g6626 = OR(g5934, g123)
--	I6350 = OR(g2445, g2437, g2433, g2419)
--	g11325 = OR(g11295, g11165)
--	I5366 = OR(g1280, g1284, g1292, g1296)
--	I5649 = OR(g1499, g1486, g1482)
--	g6894 = OR(g6763, g4868)
--	g9738 = OR(g9417, g9447, g9506)
--	g8383 = OR(g8163, g5051)
--	g8779 = OR(g5530, g8663)
--	g8161 = OR(g8005, g7185)
--	g8451 = OR(g3440, g8366)
--	g9915 = OR(g9853, g9693)
--	g2316 = OR(g1300, g1304, g1270, I5366)
--	g5576 = OR(g4675, g3664)
--	g10857 = OR(g6090, g10738)
--	g10793 = OR(g6194, g10763)
--	g7511 = OR(g6890, g6438)
--	g8944 = OR(g8799, g8708)
--	g10765 = OR(g5492, g10680)
--	g10549 = OR(g4951, g10451)
--	g7092 = OR(g6540, g5902)
--	g11604 = OR(g11583, g11554)
--	g8434 = OR(g8400, g8074)
--	g6546 = OR(g5796, g5026)
--	g3354 = OR(g2920, g2124)
--	g9928 = OR(g9870, g9717)
--	g11262 = OR(g11240, g11024)
--	g9785 = OR(g9010, g8995, g9388, g9363)
--	g5867 = OR(g3440, g4921)
--	g8210 = OR(g7466, g7995)
--	g10533 = OR(g4933, g10449)
--	g9563 = OR(g9052, g9030)
--	g6906 = OR(g6791, g5674)
--	g7375 = OR(g7230, g6745)
--	g7651 = OR(g7135, g4084)
--	I5570 = OR(g416, g411, g406, g401)
--	g9731 = OR(g9641, g9364, g9387)
--	g11247 = OR(g11097, g10949)
--	I15045 = OR(g7853, g9676, g9624, g9785)
--	g10856 = OR(g6083, g10737)
--	g9557 = OR(g9052, g9030)
--	g7184 = OR(g6625, g6047)
--	g11612 = OR(g11599, g11590)
--	g7384 = OR(g7088, g6618)
--	g11324 = OR(g11271, g11164)
--	g8922 = OR(g8822, g8736)
--	I5358 = OR(g1245, g1240, g1235, g1275)
--	g9955 = OR(g9947, g9941, g9808)
--	g2501 = OR(g448, g452, g421, I5576)
--	g7231 = OR(g6673, g6087)
--	g6078 = OR(g4503, g5256)
--	g6478 = OR(g5706, g4967)
--	g6907 = OR(g6792, g5675)
--	g6035 = OR(g5518, g3974)
--	g8937 = OR(g8786, g8698)
--	g7742 = OR(g7217, g6743)
--	g10722 = OR(g10308, g10671)
--	g9918 = OR(g9858, g9698)
--	g5403 = OR(g4486, g3695)
--	g7926 = OR(g7435, g6892)
--	g6915 = OR(g6347, g5686)
--	g5841 = OR(g4914, g4230)
--	I15220 = OR(g9841, g9966, g9857, g9877)
--	g10529 = OR(I16160, I16161)
--	g11246 = OR(g11094, g10948)
--	g6002 = OR(g5489, g3939)
--	g7712 = OR(g7125, g3540)
--	g8810 = OR(g7933, g8720)
--	g9921 = OR(g9862, g9703)
--	g8432 = OR(g8389, g8072)
--	I15172 = OR(g9843, g9959, g9861, g9874)
--	I14822 = OR(g9597, g9604, g9582)
--	g6928 = OR(g6359, g5703)
--	g8157 = OR(g7965, g7623)
--	g6930 = OR(g6364, g4269)
--	g7660 = OR(g7059, g6583)
--	g6899 = OR(g6463, g5471)
--	g9392 = OR(g9328, g9324)
--	g11318 = OR(g11228, g11104)
--	I16427 = OR(g10683, g10608, g10604)
--	g11227 = OR(g11151, g11010)
--	g11058 = OR(g10933, g5280)
--	I5351 = OR(g1145, g1141, g1137, g1133)
--	g9708 = OR(g9653, g9389, g9646)
--	g6071 = OR(g5228, g4505)
--	g9911 = OR(g9846, g9689)
--	g7102 = OR(g6550, g5915)
--	g7302 = OR(g7141, g6328)
--	g6038 = OR(g5528, g3979)
--	g4239 = OR(g4000, g4008)
--	g8646 = OR(g8224, g8547)
--	g9974 = OR(I15176, I15177)
--	g5823 = OR(g5631, g4882)
--	g6918 = OR(g6358, g4252)
--	g7265 = OR(g6756, g6204)
--	I5804 = OR(g2111, g2109, g2106, g2104)
--	g5851 = OR(g4941, g4253)
--	g11481 = OR(g6624, g11458)
--	g10336 = OR(g10230, g9572)
--	g7296 = OR(g7131, g6322)
--	g4300 = OR(g3546, g2391)
--	g8647 = OR(g8130, g8470)
--	
--	g8546 = NAND(g3983, g8390)
--	g2516 = NAND(I5612, I5613)
--	g2987 = NAND(g2481, g883)
--	I5593 = NAND(g1703, I5591)
--	g8970 = NAND(g5548, g8839)
--	I10519 = NAND(g6231, g822)
--	I11279 = NAND(g305, I11278)
--	g7990 = NAND(g7011, g6995, g7562, g7550)
--	I11278 = NAND(g305, g6485)
--	g3978 = NAND(g3207, g1822)
--	I5264 = NAND(g456, I5263)
--	I8640 = NAND(g4278, g516)
--	I6761 = NAND(g2943, I6760)
--	I17400 = NAND(g11418, g11416)
--	I5450 = NAND(g1235, I5449)
--	I16060 = NAND(g10372, I16058)
--	I6746 = NAND(g2938, g1453)
--	I11975 = NAND(g1462, I11973)
--	I12136 = NAND(g7110, g131)
--	I11937 = NAND(g1458, I11935)
--	g2959 = NAND(I6167, I6168)
--	I5878 = NAND(g2120, g2115)
--	g2517 = NAND(I5619, I5620)
--	g5552 = NAND(g4777, g4401)
--	I6468 = NAND(g23, I6467)
--	I8796 = NAND(g4672, I8795)
--	g10392 = NAND(I15891, I15892)
--	I5611 = NAND(g1280, g1284)
--	g8738 = NAND(g8688, g4921)
--	I6716 = NAND(g201, I6714)
--	g2310 = NAND(g591, g605)
--	I7685 = NAND(g3460, I7683)
--	g3056 = NAND(g2374, g599)
--	I12108 = NAND(g135, I12106)
--	g3529 = NAND(g2310, g3062, g2325)
--	I6747 = NAND(g2938, I6746)
--	g2236 = NAND(I5230, I5231)
--	g7584 = NAND(I12075, I12076)
--	I15870 = NAND(g10358, g2713)
--	I16067 = NAND(g2765, I16065)
--	I7562 = NAND(g3533, g654)
--	I13531 = NAND(g8253, I13529)
--	I8797 = NAND(g1145, I8795)
--	I17584 = NAND(g11354, g11515)
--	I11936 = NAND(g7004, I11935)
--	I15257 = NAND(g9984, I15256)
--	g8402 = NAND(I13505, I13506)
--	g8824 = NAND(g8502, g8501, g8739)
--	I6186 = NAND(g2511, g466)
--	g11496 = NAND(I17504, I17505)
--	I16001 = NAND(g2683, I15999)
--	I6125 = NAND(g2215, I6124)
--	I11909 = NAND(g1474, I11907)
--	I12040 = NAND(g1466, I12038)
--	I13909 = NAND(g1432, I13907)
--	g3625 = NAND(I6771, I6772)
--	I11908 = NAND(g6967, I11907)
--	g10470 = NAND(I16008, I16009)
--	I13908 = NAND(g8526, I13907)
--	g3813 = NAND(I7034, I7035)
--	I8650 = NAND(g4824, g778)
--	g6207 = NAND(I9947, I9948)
--	I16066 = NAND(g10428, I16065)
--	g2948 = NAND(I6144, I6145)
--	I11242 = NAND(g6760, I11241)
--	g10467 = NAND(I15993, I15994)
--	I6187 = NAND(g2511, I6186)
--	g6488 = NAND(g6027, g6019)
--	I5500 = NAND(g1255, g1007)
--	I11974 = NAND(g7001, I11973)
--	I12062 = NAND(g1478, I12060)
--	g5300 = NAND(I8771, I8772)
--	I5184 = NAND(g1415, g1515)
--	I13293 = NAND(g1882, g8161)
--	I6200 = NAND(g2525, I6199)
--	I13265 = NAND(g1909, g8154)
--	I5024 = NAND(g995, I5023)
--	I7863 = NAND(g4099, g774)
--	g8705 = NAND(I13991, I13992)
--	g8471 = NAND(I13660, I13661)
--	I15256 = NAND(g9984, g9980)
--	I6145 = NAND(g646, I6143)
--	I13992 = NAND(g8688, I13990)
--	I11510 = NAND(g1806, I11508)
--	g10853 = NAND(g10731, g5034)
--	I5231 = NAND(g148, I5229)
--	I12047 = NAND(g1486, I12045)
--	I10771 = NAND(g1801, I10769)
--	g10477 = NAND(I16045, I16046)
--	g7582 = NAND(I12061, I12062)
--	I5104 = NAND(g431, g435)
--	g8409 = NAND(I13530, I13531)
--	I6447 = NAND(g2264, g1776)
--	I4956 = NAND(g327, I4954)
--	I5613 = NAND(g1284, I5611)
--	I8481 = NAND(g3530, I8479)
--	g5278 = NAND(I8739, I8740)
--	I6880 = NAND(g3301, I6879)
--	I15431 = NAND(g10047, I15430)
--	g5548 = NAND(g1840, g4401)
--	g7671 = NAND(g7011, g6995, g6984, g6974)
--	I12020 = NAND(g7119, I12019)
--	g10665 = NAND(I16331, I16332)
--	I16469 = NAND(g10518, I16467)
--	I5014 = NAND(g1007, I5013)
--	I13523 = NAND(g8249, I13521)
--	I16039 = NAND(g2707, I16037)
--	I16468 = NAND(g10716, I16467)
--	I12046 = NAND(g6951, I12045)
--	g4476 = NAND(g3807, g3071)
--	g10476 = NAND(I16038, I16039)
--	I16038 = NAND(g10427, I16037)
--	I8676 = NAND(g4374, g1027)
--	I12113 = NAND(g7093, g162)
--	I8761 = NAND(g4616, g1129)
--	g3204 = NAND(g2571, g2061)
--	I15993 = NAND(g10422, I15992)
--	I5036 = NAND(g1019, I5034)
--	I14263 = NAND(g8843, g1814)
--	g8298 = NAND(I13249, I13250)
--	I5135 = NAND(g521, g525)
--	g2405 = NAND(I5485, I5486)
--	I7034 = NAND(g3089, I7033)
--	I15443 = NAND(g10122, I15441)
--	I6166 = NAND(g2236, g153)
--	I8624 = NAND(g4267, g511)
--	I16015 = NAND(g10425, g2695)
--	I8677 = NAND(g4374, I8676)
--	I8576 = NAND(g4234, I8575)
--	I14613 = NAND(g9204, I14612)
--	I8716 = NAND(g4601, I8715)
--	g3530 = NAND(I6715, I6716)
--	g8405 = NAND(I13514, I13515)
--	g4104 = NAND(g3215, g3247, g2439, g3200)
--	I12003 = NAND(g7082, I12002)
--	g2177 = NAND(I5127, I5128)
--	g3010 = NAND(g2382, g2399)
--	g5179 = NAND(I8576, I8577)
--	I17395 = NAND(g11414, I17393)
--	g7067 = NAND(I11279, I11280)
--	g7994 = NAND(g7011, g7574, g6984, g7550)
--	I6167 = NAND(g2236, I6166)
--	I5265 = NAND(g461, I5263)
--	I6989 = NAND(g2760, I6988)
--	I13274 = NAND(g8158, I13272)
--	I10507 = NAND(g6221, g786)
--	I13530 = NAND(g704, I13529)
--	I5164 = NAND(g1508, g1499)
--	g9107 = NAND(I14443, I14444)
--	I9559 = NAND(g782, I9557)
--	I8577 = NAND(g496, I8575)
--	g2510 = NAND(I5592, I5593)
--	g8177 = NAND(I13077, I13078)
--	I8717 = NAND(g4052, I8715)
--	I5296 = NAND(g794, I5295)
--	g5209 = NAND(I8625, I8626)
--	g7950 = NAND(g7395, g7390, g7380, g7273)
--	g2088 = NAND(I4911, I4912)
--	I16000 = NAND(g10423, I15999)
--	I5371 = NAND(g971, g976)
--	g2215 = NAND(I5185, I5186)
--	g7101 = NAND(g6617, g2364)
--	I5675 = NAND(g1218, g1223)
--	I8544 = NAND(g4218, I8543)
--	g6577 = NAND(I10520, I10521)
--	I5297 = NAND(g798, I5295)
--	I13537 = NAND(g658, g8157)
--	I13283 = NAND(g1927, g8159)
--	g4749 = NAND(g3710, g2061)
--	I11982 = NAND(g1482, I11980)
--	I8514 = NAND(g4873, I8513)
--	I13091 = NAND(g1840, I13089)
--	g2943 = NAND(I6125, I6126)
--	I15908 = NAND(g10302, I15906)
--	I6879 = NAND(g3301, g1351)
--	I8763 = NAND(g1129, I8761)
--	I5449 = NAND(g1235, g991)
--	g8825 = NAND(g8502, g8738, g8506)
--	I16007 = NAND(g10424, g2689)
--	I5865 = NAND(g2107, g2105)
--	I5604 = NAND(g1149, g1153)
--	g2433 = NAND(I5517, I5518)
--	I6111 = NAND(g1494, I6109)
--	g2096 = NAND(I4929, I4930)
--	I13522 = NAND(g695, I13521)
--	I10770 = NAND(g5944, I10769)
--	g6027 = NAND(g4566, g4921)
--	g7992 = NAND(g7011, g7574, g6984, g6974)
--	I5539 = NAND(g1270, I5538)
--	I17394 = NAND(g11415, I17393)
--	I13553 = NAND(g668, I13552)
--	I8642 = NAND(g516, I8640)
--	g7573 = NAND(I12046, I12047)
--	g11416 = NAND(I17296, I17297)
--	g6003 = NAND(g5552, g5548)
--	g8934 = NAND(I14278, I14279)
--	I15992 = NAND(g10422, g2677)
--	I7683 = NAND(g1023, g3460)
--	I4910 = NAND(g386, g318)
--	g3209 = NAND(g2550, g2061, g2564, g2571)
--	I6794 = NAND(g143, I6792)
--	I10521 = NAND(g822, I10519)
--	I5486 = NAND(g1011, I5484)
--	I15442 = NAND(g10035, I15441)
--	g6858 = NAND(I10931, I10932)
--	I5185 = NAND(g1415, I5184)
--	g5304 = NAND(I8779, I8780)
--	g2354 = NAND(g1515, g1520)
--	I15615 = NAND(g10043, g10153)
--	I17281 = NAND(g11360, g11357)
--	I5470 = NAND(g999, I5468)
--	I11509 = NAND(g6580, I11508)
--	I5025 = NAND(g1275, I5023)
--	I11508 = NAND(g6580, g1806)
--	I15430 = NAND(g10047, g10044)
--	I14612 = NAND(g9204, g611)
--	g4675 = NAND(g4073, g3247)
--	I14272 = NAND(g1822, I14270)
--	g2979 = NAND(I6208, I6209)
--	I17290 = NAND(g11363, I17288)
--	g5269 = NAND(I8716, I8717)
--	g4297 = NAND(I7563, I7564)
--	I12002 = NAND(g7082, g153)
--	I5006 = NAND(g421, I5005)
--	I12128 = NAND(g170, I12126)
--	I5105 = NAND(g431, I5104)
--	I6323 = NAND(g2050, I6322)
--	g7588 = NAND(I12093, I12094)
--	I6666 = NAND(g2776, I6664)
--	g3623 = NAND(I6761, I6762)
--	I5373 = NAND(g976, I5371)
--	I8529 = NAND(g481, I8527)
--	I5283 = NAND(g758, I5282)
--	I7224 = NAND(g2981, I7223)
--	I5007 = NAND(g312, I5005)
--	I5459 = NAND(g1240, g1003)
--	I17297 = NAND(g11369, I17295)
--	g8746 = NAND(g8617, g6517, g6509)
--	I6143 = NAND(g1976, g646)
--	I5015 = NAND(g1011, I5013)
--	g8932 = NAND(I14264, I14265)
--	I16073 = NAND(g845, I16072)
--	I6988 = NAND(g2760, g986)
--	g3205 = NAND(g1814, g2571)
--	I8652 = NAND(g778, I8650)
--	I9558 = NAND(g5598, I9557)
--	I5203 = NAND(g369, I5202)
--	g7533 = NAND(I11936, I11937)
--	g3634 = NAND(I6806, I6807)
--	I6792 = NAND(g2959, g143)
--	g3304 = NAND(I6468, I6469)
--	I12145 = NAND(g158, I12143)
--	g7596 = NAND(I12127, I12128)
--	I13302 = NAND(g8162, I13300)
--	I5502 = NAND(g1007, I5500)
--	I9574 = NAND(g5608, g818)
--	g3273 = NAND(I6448, I6449)
--	I8670 = NAND(g4831, I8669)
--	I7035 = NAND(g1868, I7033)
--	I15453 = NAND(g10051, I15451)
--	I8625 = NAND(g4267, I8624)
--	I7876 = NAND(g4109, I7875)
--	I14203 = NAND(g8825, I14202)
--	I15607 = NAND(g10149, g10144)
--	g2274 = NAND(I5324, I5325)
--	I8740 = NAND(g1121, I8738)
--	I17296 = NAND(g11373, I17295)
--	g10507 = NAND(g10434, g5859)
--	g2325 = NAND(g611, g617)
--	I8606 = NAND(g506, I8604)
--	I12087 = NAND(g1470, I12085)
--	I13249 = NAND(g1891, I13248)
--	I13248 = NAND(g1891, g8148)
--	I13552 = NAND(g668, g8262)
--	g2106 = NAND(I4979, I4980)
--	I12069 = NAND(g139, I12067)
--	g9204 = NAND(g6019, g8942)
--	I12068 = NAND(g7116, I12067)
--	I17503 = NAND(g11475, g7603)
--	I7877 = NAND(g810, I7875)
--	I5165 = NAND(g1508, I5164)
--	g6740 = NAND(g6131, g2550)
--	I6289 = NAND(g981, I6287)
--	I6777 = NAND(g2892, g650)
--	g5171 = NAND(I8562, I8563)
--	I15891 = NAND(g853, I15890)
--	I13090 = NAND(g8006, I13089)
--	g11474 = NAND(I17460, I17461)
--	g7942 = NAND(g7395, g6847, g7380, g7369)
--	I5538 = NAND(g1270, g1023)
--	I7563 = NAND(g3533, I7562)
--	I13513 = NAND(g686, g8248)
--	g2107 = NAND(I4986, I4987)
--	g2223 = NAND(I5203, I5204)
--	I13505 = NAND(g677, I13504)
--	I6209 = NAND(g802, I6207)
--	I12086 = NAND(g6980, I12085)
--	I8545 = NAND(g486, I8543)
--	I8180 = NAND(g1786, I8178)
--	g2115 = NAND(I5014, I5015)
--	I8591 = NAND(g501, I8589)
--	I10931 = NAND(g6395, I10930)
--	I17402 = NAND(g11416, I17400)
--	g8307 = NAND(I13294, I13295)
--	I12144 = NAND(g7089, I12143)
--	I10520 = NAND(g6231, I10519)
--	I5263 = NAND(g456, g461)
--	g8757 = NAND(g8599, g4401)
--	I6714 = NAND(g2961, g201)
--	I14211 = NAND(g599, I14209)
--	I8515 = NAND(g3513, I8513)
--	g2272 = NAND(I5316, I5317)
--	I9946 = NAND(g5233, g1796)
--	I8750 = NAND(g4613, g1125)
--	I5605 = NAND(g1149, I5604)
--	g8880 = NAND(I14203, I14204)
--	I16051 = NAND(g837, g10371)
--	I16072 = NAND(g845, g10373)
--	g10440 = NAND(g10360, g6037)
--	g8612 = NAND(I13858, I13859)
--	I15872 = NAND(g2713, I15870)
--	I8528 = NAND(g4879, I8527)
--	g8629 = NAND(I13901, I13902)
--	g8542 = NAND(g2571, g1828, g1814, g8390)
--	I9947 = NAND(g5233, I9946)
--	I6838 = NAND(g806, I6836)
--	g7583 = NAND(I12068, I12069)
--	g4803 = NAND(g3664, g2356)
--	I17307 = NAND(g11377, I17305)
--	g4538 = NAND(g3475, g2399)
--	I15452 = NAND(g10058, I15451)
--	I13857 = NAND(g8538, g1448)
--	I14202 = NAND(g8825, g591)
--	I13765 = NAND(g731, g8417)
--	g2260 = NAND(I5296, I5297)
--	g7986 = NAND(g7011, g6995, g6984, g7550)
--	g5226 = NAND(I8670, I8671)
--	g8512 = NAND(g3723, g8366)
--	I16046 = NAND(g10370, I16044)
--	I13504 = NAND(g677, g8247)
--	g10447 = NAND(g10363, g5360)
--	g2167 = NAND(I5105, I5106)
--	I8804 = NAND(g4677, I8803)
--	g10472 = NAND(I16016, I16017)
--	I17487 = NAND(g11474, I17485)
--	I4995 = NAND(g416, g309)
--	I12093 = NAND(g6944, I12092)
--	g7987 = NAND(g7011, g6995, g7562, g6974)
--	g5227 = NAND(I8677, I8678)
--	I5126 = NAND(g1386, g1389)
--	g2321 = NAND(I5372, I5373)
--	g7547 = NAND(I11974, I11975)
--	I17306 = NAND(g11381, I17305)
--	g6548 = NAND(g6132, g6124, g6122)
--	I11995 = NAND(g7107, g127)
--	I7225 = NAND(g1781, I7223)
--	I11261 = NAND(g6775, g826)
--	g8843 = NAND(g8542, g8757, g8545)
--	g2938 = NAND(I6110, I6111)
--	I4942 = NAND(g396, I4941)
--	g10394 = NAND(I15899, I15900)
--	g8549 = NAND(g5527, g8390)
--	g3070 = NAND(g2016, g1206)
--	I4954 = NAND(g401, g327)
--	I5023 = NAND(g995, g1275)
--	g10446 = NAND(g10443, g5350)
--	I16081 = NAND(g10374, I16079)
--	I8641 = NAND(g4278, I8640)
--	I6178 = NAND(g197, I6176)
--	I12075 = NAND(g7098, I12074)
--	I5127 = NAND(g1386, I5126)
--	I5451 = NAND(g991, I5449)
--	g4168 = NAND(I7322, I7323)
--	I6288 = NAND(g2091, I6287)
--	I8179 = NAND(g3685, I8178)
--	I4912 = NAND(g318, I4910)
--	I6805 = NAND(g3268, g471)
--	g3766 = NAND(g2439, g3222, g2493)
--	g3087 = NAND(I6288, I6289)
--	I17486 = NAND(g11384, I17485)
--	I4929 = NAND(g391, I4928)
--	I15890 = NAND(g853, g10286)
--	I16331 = NAND(g10616, I16330)
--	I9575 = NAND(g5608, I9574)
--	I13887 = NAND(g8532, I13886)
--	g5308 = NAND(I8787, I8788)
--	I13529 = NAND(g704, g8253)
--	I6208 = NAND(g2534, I6207)
--	g5217 = NAND(I8641, I8642)
--	I5316 = NAND(g1032, I5315)
--	g2111 = NAND(I5006, I5007)
--	g10366 = NAND(g10285, g5392)
--	I5034 = NAND(g1015, g1019)
--	I13869 = NAND(g1403, I13867)
--	I13868 = NAND(g8523, I13867)
--	I15999 = NAND(g10423, g2683)
--	I13259 = NAND(g1900, I13258)
--	g3261 = NAND(g2229, g2222, g2211, g2202)
--	g10481 = NAND(I16073, I16074)
--	g2180 = NAND(I5136, I5137)
--	g4976 = NAND(g2310, g4604, g3807)
--	g8506 = NAND(g3475, g8366)
--	g2380 = NAND(I5460, I5461)
--	I13258 = NAND(g1900, g8153)
--	I5013 = NAND(g1007, g1011)
--	g5196 = NAND(I8605, I8606)
--	I10930 = NAND(g6395, g5555)
--	I6770 = NAND(g3257, g382)
--	g11449 = NAND(I17401, I17402)
--	g11448 = NAND(I17394, I17395)
--	I15717 = NAND(g10231, I15716)
--	I5317 = NAND(g1027, I5315)
--	I14210 = NAND(g8824, I14209)
--	I17569 = NAND(g1610, I17567)
--	I13878 = NAND(g1444, I13876)
--	g8545 = NAND(g3710, g8390)
--	g2515 = NAND(I5605, I5606)
--	I14443 = NAND(g8970, I14442)
--	g7557 = NAND(I11996, I11997)
--	g8180 = NAND(I13090, I13091)
--	I14279 = NAND(g1828, I14277)
--	I17568 = NAND(g11496, I17567)
--	I13886 = NAND(g8532, g1440)
--	I7322 = NAND(g3047, I7321)
--	I6990 = NAND(g986, I6988)
--	I14278 = NAND(g8847, I14277)
--	I7033 = NAND(g3089, g1868)
--	I9006 = NAND(g4492, g1791)
--	g8507 = NAND(g3738, g8366)
--	I5460 = NAND(g1240, I5459)
--	g4588 = NAND(g3440, g2745)
--	I4986 = NAND(g999, I4985)
--	g3247 = NAND(g1828, g2564, g2571)
--	I8651 = NAND(g4824, I8650)
--	I13545 = NAND(g713, I13544)
--	g8628 = NAND(I13894, I13895)
--	I6138 = NAND(g378, I6136)
--	I12074 = NAND(g7098, g174)
--	g8630 = NAND(I13908, I13909)
--	I13078 = NAND(g7963, I13076)
--	I6109 = NAND(g2205, g1494)
--	g8300 = NAND(I13259, I13260)
--	I5501 = NAND(g1255, I5500)
--	I17586 = NAND(g11515, I17584)
--	I12092 = NAND(g6944, g1490)
--	I13901 = NAND(g8520, I13900)
--	I8795 = NAND(g4672, g1145)
--	I6201 = NAND(g766, I6199)
--	I14217 = NAND(g8826, I14216)
--	I9007 = NAND(g4492, I9006)
--	I13561 = NAND(g8263, I13559)
--	I15716 = NAND(g10231, g10229)
--	I6449 = NAND(g1776, I6447)
--	I13295 = NAND(g8161, I13293)
--	I4987 = NAND(g1003, I4985)
--	I6715 = NAND(g2961, I6714)
--	I17493 = NAND(g11475, I17492)
--	I12215 = NAND(g7061, I12214)
--	g2372 = NAND(I5450, I5451)
--	g7062 = NAND(I11262, I11263)
--	g2988 = NAND(I6225, I6226)
--	I13309 = NAND(g617, I13307)
--	g8839 = NAND(g8750, g4401)
--	g2555 = NAND(I5676, I5677)
--	g3662 = NAND(I6826, I6827)
--	I13308 = NAND(g8190, I13307)
--	g2792 = NAND(I5879, I5880)
--	g4117 = NAND(g3041, g3061)
--	I8543 = NAND(g4218, g486)
--	g11549 = NAND(I17585, I17586)
--	I6881 = NAND(g1351, I6879)
--	I12138 = NAND(g131, I12136)
--	I8729 = NAND(g4605, I8728)
--	I14216 = NAND(g8826, g605)
--	g10384 = NAND(I15871, I15872)
--	I13260 = NAND(g8153, I13258)
--	g2776 = NAND(I5866, I5867)
--	I8513 = NAND(g4873, g3513)
--	I13559 = NAND(g722, g8263)
--	I8178 = NAND(g3685, g1786)
--	g3631 = NAND(I6793, I6794)
--	I6487 = NAND(g2306, g1227)
--	I16080 = NAND(g849, I16079)
--	I13893 = NAND(g8529, g1436)
--	I12115 = NAND(g162, I12113)
--	I6748 = NAND(g1453, I6746)
--	I13544 = NAND(g713, g8259)
--	I5484 = NAND(g1250, g1011)
--	I4928 = NAND(g391, g321)
--	I6226 = NAND(g1346, I6224)
--	I8805 = NAND(g1113, I8803)
--	I4930 = NAND(g321, I4928)
--	I15880 = NAND(g2719, I15878)
--	I14265 = NAND(g1814, I14263)
--	I16031 = NAND(g829, I16030)
--	g3585 = NAND(I6747, I6748)
--	g3041 = NAND(g2364, g2399, g2374, g2382)
--	g8933 = NAND(I14271, I14272)
--	I16330 = NAND(g10616, g4997)
--	I13267 = NAND(g8154, I13265)
--	I13294 = NAND(g1882, I13293)
--	g10231 = NAND(I15616, I15617)
--	I14442 = NAND(g8970, g1834)
--	I6793 = NAND(g2959, I6792)
--	I4966 = NAND(g330, I4964)
--	I8752 = NAND(g1125, I8750)
--	I15432 = NAND(g10044, I15430)
--	I12214 = NAND(g7061, g2518)
--	g10511 = NAND(g10438, g6032)
--	g3011 = NAND(g591, g2382)
--	g5103 = NAND(I8480, I8481)
--	I16087 = NAND(g861, I16086)
--	g3734 = NAND(g3039, g599)
--	I6664 = NAND(g2792, g2776)
--	g8882 = NAND(I14217, I14218)
--	I4955 = NAND(g401, I4954)
--	I8786 = NAND(g4639, g1141)
--	g3992 = NAND(g2571, g2550, g2990)
--	g10480 = NAND(I16066, I16067)
--	I11915 = NAND(g6935, I11914)
--	I8770 = NAND(g4619, g1133)
--	I5516 = NAND(g1260, g1019)
--	g8541 = NAND(g4001, g8390)
--	I6188 = NAND(g466, I6186)
--	g5147 = NAND(I8544, I8545)
--	g8744 = NAND(g8617, g6509, g6971)
--	I5892 = NAND(g750, I5891)
--	g8558 = NAND(I13766, I13767)
--	I15258 = NAND(g9980, I15256)
--	I13266 = NAND(g1909, I13265)
--	I8787 = NAND(g4639, I8786)
--	I6826 = NAND(g3281, I6825)
--	I17283 = NAND(g11357, I17281)
--	g5013 = NAND(g4749, g3247, g3205)
--	I17492 = NAND(g11475, g3623)
--	g8511 = NAND(g5277, g8366)
--	I16079 = NAND(g849, g10374)
--	I5035 = NAND(g1015, I5034)
--	I5517 = NAND(g1260, I5516)
--	I7223 = NAND(g2981, g1781)
--	I16086 = NAND(g861, g10375)
--	g5317 = NAND(I8796, I8797)
--	I15879 = NAND(g10359, I15878)
--	I15878 = NAND(g10359, g2719)
--	I12114 = NAND(g7093, I12113)
--	I12107 = NAND(g7113, I12106)
--	g2500 = NAND(g178, g182)
--	I15994 = NAND(g2677, I15992)
--	g7934 = NAND(g7395, g6847, g7279, g7369)
--	g10469 = NAND(g10430, g5999)
--	I14264 = NAND(g8843, I14263)
--	I6448 = NAND(g2264, I6447)
--	I13285 = NAND(g8159, I13283)
--	g10468 = NAND(I16000, I16001)
--	I6827 = NAND(g770, I6825)
--	g8623 = NAND(I13877, I13878)
--	I13900 = NAND(g8520, g1428)
--	g2795 = NAND(I5892, I5893)
--	I8575 = NAND(g4234, g496)
--	I14209 = NAND(g8824, g599)
--	I13560 = NAND(g722, I13559)
--	I8715 = NAND(g4601, g4052)
--	I8604 = NAND(g4259, g506)
--	I16017 = NAND(g2695, I16015)
--	I4941 = NAND(g396, g324)
--	g2205 = NAND(I5165, I5166)
--	g3753 = NAND(g2382, g2364, g2800)
--	I6467 = NAND(g23, g2479)
--	I14614 = NAND(g611, I14612)
--	g2104 = NAND(I4965, I4966)
--	g2099 = NAND(I4942, I4943)
--	I16023 = NAND(g10426, g2701)
--	g10479 = NAND(I16059, I16060)
--	g8737 = NAND(g2317, g4921, g8688)
--	g5942 = NAND(I9575, I9576)
--	g10478 = NAND(I16052, I16053)
--	I12004 = NAND(g153, I12002)
--	I4911 = NAND(g386, I4910)
--	I11914 = NAND(g6935, g1494)
--	g7960 = NAND(g7409, g5573)
--	I5295 = NAND(g794, g798)
--	I12106 = NAND(g7113, g135)
--	I8728 = NAND(g4605, g1117)
--	g3681 = NAND(I6837, I6838)
--	I11907 = NAND(g6967, g1474)
--	I13907 = NAND(g8526, g1432)
--	I8730 = NAND(g1117, I8728)
--	g8551 = NAND(g3967, g8390)
--	I4980 = NAND(g333, I4978)
--	g2961 = NAND(I6177, I6178)
--	g6019 = NAND(g617, g4921)
--	I16016 = NAND(g10425, I16015)
--	I11935 = NAND(g7004, g1458)
--	I8678 = NAND(g1027, I8676)
--	I17051 = NAND(g10923, g11249)
--	g4482 = NAND(I7864, I7865)
--	g7592 = NAND(I12107, I12108)
--	g3460 = NAND(I6665, I6666)
--	g7932 = NAND(g7395, g6847, g7279, g7273)
--	g7624 = NAND(I12215, I12216)
--	g7953 = NAND(g7395, g7390, g7380, g7369)
--	g8414 = NAND(I13553, I13554)
--	I6168 = NAND(g153, I6166)
--	I5229 = NAND(g182, g148)
--	I6772 = NAND(g382, I6770)
--	I16030 = NAND(g829, g10368)
--	I13284 = NAND(g1927, I13283)
--	I16065 = NAND(g10428, g2765)
--	g2947 = NAND(I6137, I6138)
--	I7321 = NAND(g3047, g1231)
--	g2437 = NAND(I5529, I5530)
--	g2102 = NAND(I4955, I4956)
--	I17282 = NAND(g11360, I17281)
--	I5620 = NAND(g1771, I5618)
--	I8664 = NAND(g476, I8662)
--	g7524 = NAND(I11915, I11916)
--	g7717 = NAND(g6863, g3206)
--	I16467 = NAND(g10716, g10518)
--	I4972 = NAND(g991, I4971)
--	I13554 = NAND(g8262, I13552)
--	I16037 = NAND(g10427, g2707)
--	g8302 = NAND(I13273, I13274)
--	I4943 = NAND(g324, I4941)
--	I5485 = NAND(g1250, I5484)
--	g5527 = NAND(g3978, g4749)
--	I10509 = NAND(g786, I10507)
--	g7599 = NAND(I12144, I12145)
--	I10508 = NAND(g6221, I10507)
--	I6126 = NAND(g1419, I6124)
--	I8671 = NAND(g814, I8669)
--	I6760 = NAND(g2943, g1448)
--	g3626 = NAND(I6778, I6779)
--	I11973 = NAND(g7001, g1462)
--	g2389 = NAND(I5469, I5470)
--	I15617 = NAND(g10153, I15615)
--	g5277 = NAND(g3734, g4538)
--	I5005 = NAND(g421, g312)
--	I6779 = NAND(g650, I6777)
--	I6665 = NAND(g2792, I6664)
--	I8589 = NAND(g4251, g501)
--	g8412 = NAND(I13545, I13546)
--	g2963 = NAND(I6187, I6188)
--	I12045 = NAND(g6951, g1486)
--	I16053 = NAND(g10371, I16051)
--	g2109 = NAND(I4996, I4997)
--	g11418 = NAND(I17306, I17307)
--	I13539 = NAND(g8157, I13537)
--	g10475 = NAND(I16031, I16032)
--	I5324 = NAND(g1336, I5323)
--	I13538 = NAND(g658, I13537)
--	I5469 = NAND(g1245, I5468)
--	I5540 = NAND(g1023, I5538)
--	I17505 = NAND(g7603, I17503)
--	I11241 = NAND(g6760, g790)
--	I8803 = NAND(g4677, g1113)
--	I12061 = NAND(g6961, I12060)
--	I8780 = NAND(g1137, I8778)
--	g8745 = NAND(g8617, g6517, g6964)
--	I4979 = NAND(g411, I4978)
--	g8109 = NAND(g5052, g7853)
--	g8309 = NAND(I13308, I13309)
--	g6758 = NAND(I10770, I10771)
--	I16009 = NAND(g2689, I16007)
--	I15616 = NAND(g10043, I15615)
--	I8662 = NAND(g4286, g476)
--	I16008 = NAND(g10424, I16007)
--	I13515 = NAND(g8248, I13513)
--	I13991 = NAND(g622, I13990)
--	g11276 = NAND(I17052, I17053)
--	I15900 = NAND(g10287, I15898)
--	g2419 = NAND(I5501, I5502)
--	I16074 = NAND(g10373, I16072)
--	I10769 = NAND(g5944, g1801)
--	I7323 = NAND(g1231, I7321)
--	g7978 = NAND(g7697, g3038)
--	I7875 = NAND(g4109, g810)
--	I8562 = NAND(g4227, I8561)
--	I15892 = NAND(g10286, I15890)
--	g3771 = NAND(I6989, I6990)
--	I8605 = NAND(g4259, I8604)
--	g10153 = NAND(I15452, I15453)
--	g5295 = NAND(I8762, I8763)
--	I8751 = NAND(g4613, I8750)
--	I15907 = NAND(g6899, I15906)
--	I5136 = NAND(g521, I5135)
--	I11263 = NAND(g826, I11261)
--	I14204 = NAND(g591, I14202)
--	g8881 = NAND(I14210, I14211)
--	g2105 = NAND(I4972, I4973)
--	g5557 = NAND(g4538, g3071, g3011)
--	I5230 = NAND(g182, I5229)
--	I8669 = NAND(g4831, g814)
--	g10474 = NAND(I16024, I16025)
--	I8772 = NAND(g1133, I8770)
--	g2445 = NAND(I5539, I5540)
--	g8006 = NAND(g5552, g7717)
--	I10932 = NAND(g5555, I10930)
--	I17504 = NAND(g11475, I17503)
--	I5137 = NAND(g525, I5135)
--	g8305 = NAND(I13284, I13285)
--	I5891 = NAND(g750, g2057)
--	I13273 = NAND(g1918, I13272)
--	I8480 = NAND(g4455, I8479)
--	g4144 = NAND(g2160, g3044)
--	I15906 = NAND(g6899, g10302)
--	I5342 = NAND(g315, I5341)
--	I13514 = NAND(g686, I13513)
--	g8407 = NAND(I13522, I13523)
--	g4088 = NAND(I7224, I7225)
--	g4488 = NAND(I7876, I7877)
--	g7598 = NAND(I12137, I12138)
--	g3222 = NAND(g2557, g1814, g1834)
--	I16052 = NAND(g837, I16051)
--	I12127 = NAND(g7103, I12126)
--	g10483 = NAND(I16087, I16088)
--	g8415 = NAND(I13560, I13561)
--	g11415 = NAND(I17289, I17290)
--	g6573 = NAND(I10508, I10509)
--	I5676 = NAND(g1218, I5675)
--	I6778 = NAND(g2892, I6777)
--	g9413 = NAND(I14613, I14614)
--	I8779 = NAND(g4630, I8778)
--	I5592 = NAND(g1696, I5591)
--	g8502 = NAND(g2382, g605, g591, g8366)
--	I15609 = NAND(g10144, I15607)
--	I15608 = NAND(g10149, I15607)
--	g3071 = NAND(g605, g2374, g2382)
--	g10509 = NAND(g10436, g6023)
--	I17461 = NAND(g11448, I17459)
--	I13506 = NAND(g8247, I13504)
--	I5468 = NAND(g1245, g999)
--	g5219 = NAND(I8651, I8652)
--	I5677 = NAND(g1223, I5675)
--	g8826 = NAND(g8739, g8737, g8648)
--	I17393 = NAND(g11415, g11414)
--	I5866 = NAND(g2107, I5865)
--	I12126 = NAND(g7103, g170)
--	I4978 = NAND(g411, g333)
--	g7587 = NAND(I12086, I12087)
--	g5286 = NAND(I8751, I8752)
--	g8308 = NAND(I13301, I13302)
--	I7864 = NAND(g4099, I7863)
--	I11981 = NAND(g6957, I11980)
--	I12060 = NAND(g6961, g1478)
--	g5225 = NAND(I8663, I8664)
--	g11538 = NAND(I17568, I17569)
--	I13767 = NAND(g8417, I13765)
--	g10396 = NAND(I15907, I15908)
--	I11262 = NAND(g6775, I11261)
--	I13990 = NAND(g622, g8688)
--	I6224 = NAND(g2544, g1346)
--	I5867 = NAND(g2105, I5865)
--	g2493 = NAND(g1834, g1840)
--	I5893 = NAND(g2057, I5891)
--	g3062 = NAND(g2369, g591, g611)
--	I13521 = NAND(g695, g8249)
--	I5186 = NAND(g1515, I5184)
--	I6771 = NAND(g3257, I6770)
--	I5325 = NAND(g1341, I5323)
--	I17459 = NAND(g11449, g11448)
--	I9557 = NAND(g5598, g782)
--	g11414 = NAND(I17282, I17283)
--	I12067 = NAND(g7116, g139)
--	I12094 = NAND(g1490, I12092)
--	I4964 = NAND(g406, g330)
--	I13272 = NAND(g1918, g8158)
--	I9948 = NAND(g1796, I9946)
--	g10302 = NAND(I15717, I15718)
--	I16332 = NAND(g4997, I16330)
--	I5106 = NAND(g435, I5104)
--	g8847 = NAND(g8760, g8683)
--	g2257 = NAND(I5283, I5284)
--	I12019 = NAND(g7119, g166)
--	I15441 = NAND(g10035, g10122)
--	I11997 = NAND(g127, I11995)
--	I8739 = NAND(g4607, I8738)
--	I5461 = NAND(g1003, I5459)
--	I13766 = NAND(g731, I13765)
--	I8479 = NAND(g4455, g3530)
--	I17295 = NAND(g11373, g11369)
--	I14271 = NAND(g8840, I14270)
--	I4971 = NAND(g991, g995)
--	g8301 = NAND(I13266, I13267)
--	I6110 = NAND(g2205, I6109)
--	g10482 = NAND(I16080, I16081)
--	g10779 = NAND(I16468, I16469)
--	I6762 = NAND(g1448, I6760)
--	I17289 = NAND(g11366, I17288)
--	I5315 = NAND(g1032, g1027)
--	I17288 = NAND(g11366, g11363)
--	I13859 = NAND(g1448, I13857)
--	g7548 = NAND(I11981, I11982)
--	I13858 = NAND(g8538, I13857)
--	I11996 = NAND(g7107, I11995)
--	g8743 = NAND(g8617, g6971, g6964)
--	I5880 = NAND(g2115, I5878)
--	g10513 = NAND(g10441, g5345)
--	g8411 = NAND(I13538, I13539)
--	I8626 = NAND(g511, I8624)
--	g10505 = NAND(g10432, g5938)
--	I5612 = NAND(g1280, I5611)
--	g4821 = NAND(I8179, I8180)
--	I12076 = NAND(g174, I12074)
--	I12085 = NAND(g6980, g1470)
--	g7567 = NAND(I12020, I12021)
--	I5128 = NAND(g1389, I5126)
--	I6489 = NAND(g1227, I6487)
--	g7593 = NAND(I12114, I12115)
--	I8778 = NAND(g4630, g1137)
--	g10149 = NAND(I15442, I15443)
--	I13902 = NAND(g1428, I13900)
--	I13301 = NAND(g1936, I13300)
--	g3215 = NAND(g2564, g1822)
--	g7996 = NAND(g7011, g7574, g7562, g6974)
--	I4985 = NAND(g999, g1003)
--	I14444 = NAND(g1834, I14442)
--	g8000 = NAND(g7011, g7574, g7562, g7550)
--	I5166 = NAND(g1499, I5164)
--	I17460 = NAND(g11449, I17459)
--	g3008 = NAND(g2444, g878)
--	I6836 = NAND(g3287, g806)
--	I5529 = NAND(g1265, I5528)
--	g10229 = NAND(I15608, I15609)
--	I13661 = NAND(g8322, I13659)
--	I13895 = NAND(g1436, I13893)
--	g2303 = NAND(I5342, I5343)
--	I12039 = NAND(g6990, I12038)
--	g5592 = NAND(I9007, I9008)
--	I12038 = NAND(g6990, g1466)
--	g3322 = NAND(I6488, I6489)
--	I8561 = NAND(g4227, g491)
--	I8527 = NAND(g4879, g481)
--	I12143 = NAND(g7089, g158)
--	I5619 = NAND(g1766, I5618)
--	g10386 = NAND(I15879, I15880)
--	I11980 = NAND(g6957, g1482)
--	I6837 = NAND(g3287, I6836)
--	I4973 = NAND(g995, I4971)
--	I13888 = NAND(g1440, I13886)
--	g7558 = NAND(I12003, I12004)
--	I17494 = NAND(g3623, I17492)
--	g11491 = NAND(I17493, I17494)
--	I16045 = NAND(g833, I16044)
--	I7684 = NAND(g1023, I7683)
--	g4130 = NAND(g3044, g2518)
--	I8771 = NAND(g4619, I8770)
--	I13546 = NAND(g8259, I13544)
--	I13089 = NAND(g8006, g1840)
--	g2117 = NAND(I5024, I5025)
--	g5119 = NAND(I8514, I8515)
--	g5319 = NAND(I8804, I8805)
--	I15899 = NAND(g857, I15898)
--	I5606 = NAND(g1153, I5604)
--	I15898 = NAND(g857, g10287)
--	I16032 = NAND(g10368, I16030)
--	I17401 = NAND(g11418, I17400)
--	I13659 = NAND(g1945, g8322)
--	I8738 = NAND(g4607, g1121)
--	I13250 = NAND(g8148, I13248)
--	I15718 = NAND(g10229, I15716)
--	I9008 = NAND(g1791, I9006)
--	I6176 = NAND(g2177, g197)
--	I7865 = NAND(g774, I7863)
--	g5274 = NAND(I8729, I8730)
--	I5341 = NAND(g315, g426)
--	I17305 = NAND(g11381, g11377)
--	I17053 = NAND(g11249, I17051)
--	g5125 = NAND(I8528, I8529)
--	I12216 = NAND(g2518, I12214)
--	I6225 = NAND(g2544, I6224)
--	I5879 = NAND(g2120, I5878)
--	g3221 = NAND(g1834, g2564)
--	I14270 = NAND(g8840, g1822)
--	I6124 = NAND(g2215, g1419)
--	I6324 = NAND(g1864, I6322)
--	I13867 = NAND(g8523, g1403)
--	I13894 = NAND(g8529, I13893)
--	I6469 = NAND(g2479, I6467)
--	I8663 = NAND(g4286, I8662)
--	g7523 = NAND(I11908, I11909)
--	I6177 = NAND(g2177, I6176)
--	g5187 = NAND(I8590, I8591)
--	I6287 = NAND(g2091, g981)
--	I8762 = NAND(g4616, I8761)
--	I15871 = NAND(g10358, I15870)
--	g8840 = NAND(g8542, g8541, g8760)
--	g2250 = NAND(I5264, I5265)
--	I8590 = NAND(g4251, I8589)
--	I6199 = NAND(g2525, g766)
--	I14218 = NAND(g605, I14216)
--	g8190 = NAND(g6027, g7978)
--	I5284 = NAND(g762, I5282)
--	I17485 = NAND(g11384, g11474)
--	I4965 = NAND(g406, I4964)
--	I5591 = NAND(g1696, g1703)
--	g8501 = NAND(g3760, g8366)
--	I15451 = NAND(g10058, g10051)
--	g8942 = NAND(g8823, g4921)
--	I13877 = NAND(g8535, I13876)
--	g7269 = NAND(I11509, I11510)
--	I4996 = NAND(g416, I4995)
--	I6144 = NAND(g1976, I6143)
--	I17567 = NAND(g11496, g1610)
--	g7572 = NAND(I12039, I12040)
--	I6207 = NAND(g2534, g802)
--	I14277 = NAND(g8847, g1828)
--	I16059 = NAND(g841, I16058)
--	I16025 = NAND(g2701, I16023)
--	I8563 = NAND(g491, I8561)
--	g3524 = NAND(g3209, g3221)
--	I16058 = NAND(g841, g10372)
--	I5204 = NAND(g374, I5202)
--	I6488 = NAND(g2306, I6487)
--	g3818 = NAND(g3056, g3071, g2310, g3003)
--	I16044 = NAND(g833, g10370)
--	g3717 = NAND(I6880, I6881)
--	I13077 = NAND(g1872, I13076)
--	g10043 = NAND(I15257, I15258)
--	I11280 = NAND(g6485, I11278)
--	I6825 = NAND(g3281, g770)
--	I4997 = NAND(g309, I4995)
--	I13300 = NAND(g1936, g8162)
--	I5323 = NAND(g1336, g1341)
--	I6136 = NAND(g2496, g378)
--	g5935 = NAND(I9558, I9559)
--	I5528 = NAND(g1265, g1015)
--	I6806 = NAND(g3268, I6805)
--	I5530 = NAND(g1015, I5528)
--	g10886 = NAND(g10807, g10805)
--	g3106 = NAND(I6323, I6324)
--	I13876 = NAND(g8535, g1444)
--	I6322 = NAND(g2050, g1864)
--	g3061 = NAND(g611, g2374)
--	g2439 = NAND(g1814, g1828)
--	g7947 = NAND(g7395, g7390, g7279, g7369)
--	I9576 = NAND(g818, I9574)
--	I13660 = NAND(g1945, I13659)
--	g3200 = NAND(g1822, g2061)
--	g4374 = NAND(I7684, I7685)
--	I11916 = NAND(g1494, I11914)
--	I5372 = NAND(g971, I5371)
--	g3003 = NAND(g599, g2399)
--	g8627 = NAND(I13887, I13888)
--	I5618 = NAND(g1766, g1771)
--	I6137 = NAND(g2496, I6136)
--	I5343 = NAND(g426, I5341)
--	I5282 = NAND(g758, g762)
--	I13307 = NAND(g8190, g617)
--	I13076 = NAND(g1872, g7963)
--	I6807 = NAND(g471, I6805)
--	I11243 = NAND(g790, I11241)
--	I17585 = NAND(g11354, I17584)
--	I12137 = NAND(g7110, I12136)
--	I7564 = NAND(g654, I7562)
--	g2970 = NAND(I6200, I6201)
--	g10144 = NAND(I15431, I15432)
--	I8788 = NAND(g1141, I8786)
--	g7054 = NAND(I11242, I11243)
--	I17052 = NAND(g10923, I17051)
--	g2120 = NAND(I5035, I5036)
--	g8616 = NAND(I13868, I13869)
--	I5202 = NAND(g369, g374)
--	I16088 = NAND(g10375, I16086)
--	I16024 = NAND(g10426, I16023)
--	g11490 = NAND(I17486, I17487)
--	I5518 = NAND(g1019, I5516)
--	g5118 = NAND(g2439, g4806, g4073)
--	I12021 = NAND(g166, I12019)
--	
--	g6392 = NOR(g5859, g5938)
--	g5938 = NOR(g2764, g4988)
--	g2478 = NOR(g1610, g1737)
--	g10374 = NOR(g10347, g3463)
--	g4278 = NOR(g3800, g2593, g2586, g3776)
--	g10424 = NOR(g10292, g4620)
--	g10383 = NOR(g10318, g2998)
--	g3118 = NOR(g2521, g2514)
--	g9815 = NOR(g9392, g9367)
--	g11077 = NOR(g10970, g10971)
--	g9746 = NOR(g9454, g9274, g9292)
--	g3879 = NOR(g3141, g2354, g2353)
--	g10285 = NOR(g10276, g3566)
--	g11480 = NOR(g11456, g4567)
--	g4076 = NOR(g1707, g2864)
--	g10570 = NOR(g10542, g10324)
--	g10239 = NOR(g9317, g10179)
--	g10594 = NOR(g10480, g10521)
--	g9426 = NOR(g9052, g9030)
--	g10382 = NOR(g10314, g2998)
--	g4672 = NOR(g3501, g2669, g2662, g3479)
--	g5360 = NOR(g2071, g4225)
--	g9387 = NOR(g9010, g9240, g9223, I14596)
--	g10438 = NOR(g10356, g3566)
--	g4613 = NOR(g3077, g3491, g2662, g2655)
--	g9391 = NOR(g9010, g9240, g9223, I14602)
--	g4572 = NOR(g3419, g3408, g3628)
--	g9757 = NOR(g9454, g9274, g9292)
--	g9416 = NOR(g9052, g9030)
--	g9874 = NOR(g9519, g9536, g9579, I15033)
--	g9654 = NOR(g9125, g9173)
--	g9880 = NOR(g9751, g9536, g9557, I15051)
--	g4873 = NOR(g3292, g2593, g2586, g3776)
--	g2807 = NOR(g22, g2320)
--	g10441 = NOR(g10351, g3566)
--	g4639 = NOR(g3501, g2669, g2662, g2655)
--	g10435 = NOR(g10332, g3507)
--	g10849 = NOR(g10739, g3903)
--	g9606 = NOR(g9125, g9111, g9173, g9151)
--	g9879 = NOR(g9747, g9536, g9566, I15048)
--	g9506 = NOR(g9052, g9030)
--	g6155 = NOR(g4974, g2864)
--	g6355 = NOR(g6032, g6023)
--	g9615 = NOR(g9052, g9030)
--	g10371 = NOR(g10344, g3463)
--	g9591 = NOR(g9125, g9151)
--	g10359 = NOR(g10227, g4620)
--	g10434 = NOR(g10352, g3566)
--	g10358 = NOR(g10226, g4620)
--	g9750 = NOR(g9454, g9274, g9292)
--	g10291 = NOR(g10247, g3113)
--	g4227 = NOR(g3292, g3793, g2586, g2579)
--	g9655 = NOR(g9010, g9240, g9223, I14776)
--	g9410 = NOR(g9010, g9240, g9223, I14607)
--	g9667 = NOR(g9125, g9111, g9173, g9151)
--	g10563 = NOR(g10539, g10322)
--	g9776 = NOR(g9392, g9367)
--	g10324 = NOR(g9317, g10244)
--	g4455 = NOR(g3543, g3419, g3408)
--	g9878 = NOR(g9754, g9536, g9560, I15045)
--	g10360 = NOR(g10277, g3566)
--	g9882 = NOR(g9742, g9536, g9563, I15057)
--	g10370 = NOR(g10343, g3463)
--	g4605 = NOR(g3077, g2669, g3485, g2655)
--	g10420 = NOR(g10329, g3744)
--	g10562 = NOR(g10483, g10529)
--	g10427 = NOR(g10296, g4620)
--	g5780 = NOR(g2112, g4921)
--	g10385 = NOR(g10321, g2998)
--	g10376 = NOR(g10323, g3113)
--	g10426 = NOR(g10294, g4620)
--	g4601 = NOR(g3077, g2669, g2662, g3479)
--	g5573 = NOR(g4117, g4432)
--	g9808 = NOR(g9392, g9367)
--	g5999 = NOR(g2753, g4953)
--	g9759 = NOR(g9454, g9274, g9292)
--	g6037 = NOR(g3305, g5614)
--	g10287 = NOR(g10275, g3463)
--	g5034 = NOR(g3524, g4593)
--	g9362 = NOR(g9010, g9240, g9223, I14585)
--	g9881 = NOR(g9516, g9536, g9573, I15054)
--	g10443 = NOR(g10353, g3566)
--	g10286 = NOR(g10271, g3463)
--	g4276 = NOR(g4065, g3261, g2500)
--	g4616 = NOR(g3077, g3491, g2662, g3479)
--	g10363 = NOR(g10355, g3566)
--	g2862 = NOR(g2315, g2305)
--	g10373 = NOR(g10346, g3463)
--	g10423 = NOR(g10290, g4620)
--	g9758 = NOR(g9454, g9274, g9292)
--	g9589 = NOR(g9125, g9173, g9151)
--	g9803 = NOR(g9392, g9367)
--	g10430 = NOR(g10349, g3566)
--	g9421 = NOR(g9052, g9030)
--	g10362 = NOR(g10228, g3507)
--	g2791 = NOR(g2187, g750)
--	g9817 = NOR(g9392, g9367)
--	g9605 = NOR(g9125, g9111, g9173, g9151)
--	g10372 = NOR(g10345, g3463)
--	g9669 = NOR(g9392, g9367)
--	g10422 = NOR(g10289, g4620)
--	g10436 = NOR(g10354, g3566)
--	g5556 = NOR(g4787, g2695, g2299, g2031)
--	g4286 = NOR(g3800, g2593, g3784, g2579)
--	g4974 = NOR(g4502, g3714)
--	g9779 = NOR(g9392, g9367)
--	g9423 = NOR(g9052, g9030)
--	g5350 = NOR(g4163, g4872)
--	g9361 = NOR(g9010, g9240, g9223, I14582)
--	g2459 = NOR(g1645, g1642, g1651, g1648)
--	g10381 = NOR(g10310, g2998)
--	g4259 = NOR(g3292, g3793, g3784, g3776)
--	g10522 = NOR(g10486, g10239)
--	g5392 = NOR(g3369, g4258)
--	g4122 = NOR(g3291, g2410, g2538)
--	g6023 = NOR(g2763, g4975)
--	g3462 = NOR(g2187, g2795)
--	g4218 = NOR(g3292, g2593, g3784, g3776)
--	g4267 = NOR(g3800, g2593, g2586, g2579)
--	g4677 = NOR(g3501, g2669, g3485, g2655)
--	g9646 = NOR(g9125, g9151)
--	g2863 = NOR(g2316, g2309)
--	g9616 = NOR(g9010, g9240, g9223, I14751)
--	g6032 = NOR(g3430, g5039)
--	g9647 = NOR(g9125, g9111, g9173, g9151)
--	g5859 = NOR(g3362, g4943)
--	g10433 = NOR(g10330, g3507)
--	g10368 = NOR(g10342, g3463)
--	g4251 = NOR(g3292, g3793, g3784, g2579)
--	g9876 = NOR(g9522, g9536, g9576, I15039)
--	g9656 = NOR(g9010, g9240, g9223, I14779)
--	g8303 = NOR(g8209, g4811)
--	g10429 = NOR(g10326, g3507)
--	g10428 = NOR(g10335, g4620)
--	g4234 = NOR(g3292, g3793, g2586, g3776)
--	g9877 = NOR(g9512, g9536, g9569, I15042)
--	g5186 = NOR(g2047, g4401)
--	g9489 = NOR(g9052, g9030)
--	g4619 = NOR(g3077, g3491, g3485, g2655)
--	g10432 = NOR(g10350, g3566)
--	g5345 = NOR(g2754, g4835)
--	g5763 = NOR(g5350, g5345)
--	g10375 = NOR(g10288, g3463)
--	g4879 = NOR(g3292, g2593, g3784, g2579)
--	g4607 = NOR(g3077, g2669, g3485, g3479)
--	g10425 = NOR(g10293, g4620)
--	g3107 = NOR(g2501, g2499)
--	g10322 = NOR(g9317, g10272)
--	g4630 = NOR(g3077, g3491, g3485, g3479)
--	g10364 = NOR(g10327, g3744)
--	g9781 = NOR(g9392, g9367)
--
-- VHDL Output
-- =============
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.MATH_REAL.ALL;

entity s15850 is
	port (
		CLK: in std_logic;
		G18: in std_logic;
		G23: in std_logic;
		G27: in std_logic;
		G28: in std_logic;
		G29: in std_logic;
		G30: in std_logic;
		G31: in std_logic;
		G41: in std_logic;
		G42: in std_logic;
		G43: in std_logic;
		G44: in std_logic;
		G45: in std_logic;
		G46: in std_logic;
		G47: in std_logic;
		G48: in std_logic;
		G82: in std_logic;
		G83: in std_logic;
		G84: in std_logic;
		G85: in std_logic;
		G86: in std_logic;
		G87: in std_logic;
		G88: in std_logic;
		G89: in std_logic;
		G90: in std_logic;
		G91: in std_logic;
		G92: in std_logic;
		G93: in std_logic;
		G94: in std_logic;
		G95: in std_logic;
		G96: in std_logic;
		G99: in std_logic;
		G100: in std_logic;
		G101: in std_logic;
		G102: in std_logic;
		G103: in std_logic;
		G104: in std_logic;
		G109: in std_logic;
		G741: in std_logic;
		G742: in std_logic;
		G743: in std_logic;
		G744: in std_logic;
		G750: in std_logic;
		G872: in std_logic;
		G873: in std_logic;
		G877: in std_logic;
		G881: in std_logic;
		G886: in std_logic;
		G889: in std_logic;
		G892: in std_logic;
		G895: in std_logic;
		G898: in std_logic;
		G901: in std_logic;
		G904: in std_logic;
		G907: in std_logic;
		G910: in std_logic;
		G913: in std_logic;
		G916: in std_logic;
		G919: in std_logic;
		G922: in std_logic;
		G925: in std_logic;
		G1170: in std_logic;
		G1173: in std_logic;
		G1176: in std_logic;
		G1179: in std_logic;
		G1182: in std_logic;
		G1185: in std_logic;
		G1188: in std_logic;
		G1191: in std_logic;
		G1194: in std_logic;
		G1197: in std_logic;
		G1200: in std_logic;
		G1203: in std_logic;
		G1696: in std_logic;
		G1700: in std_logic;
		G1712: in std_logic;
		G1960: in std_logic;
		G1961: in std_logic;
		G1957: out std_logic;
		G2355: out std_logic;
		G2601: out std_logic;
		G2602: out std_logic;
		G2603: out std_logic;
		G2604: out std_logic;
		G2605: out std_logic;
		G2606: out std_logic;
		G2607: out std_logic;
		G2608: out std_logic;
		G2609: out std_logic;
		G2610: out std_logic;
		G2611: out std_logic;
		G2612: out std_logic;
		G2648: out std_logic;
		G2986: out std_logic;
		G3007: out std_logic;
		G3069: out std_logic;
		G3327: out std_logic;
		G4171: out std_logic;
		G4172: out std_logic;
		G4173: out std_logic;
		G4174: out std_logic;
		G4175: out std_logic;
		G4176: out std_logic;
		G4177: out std_logic;
		G4178: out std_logic;
		G4179: out std_logic;
		G4180: out std_logic;
		G4181: out std_logic;
		G4191: out std_logic;
		G4192: out std_logic;
		G4193: out std_logic;
		G4194: out std_logic;
		G4195: out std_logic;
		G4196: out std_logic;
		G4197: out std_logic;
		G4198: out std_logic;
		G4199: out std_logic;
		G4200: out std_logic;
		G4201: out std_logic;
		G4202: out std_logic;
		G4203: out std_logic;
		G4204: out std_logic;
		G4205: out std_logic;
		G4206: out std_logic;
		G4207: out std_logic;
		G4208: out std_logic;
		G4209: out std_logic;
		G4210: out std_logic;
		G4211: out std_logic;
		G4212: out std_logic;
		G4213: out std_logic;
		G4214: out std_logic;
		G4215: out std_logic;
		G4216: out std_logic;
		G4887: out std_logic;
		G4888: out std_logic;
		G5101: out std_logic;
		G5105: out std_logic;
		G5658: out std_logic;
		G5659: out std_logic;
		G5816: out std_logic;
		G6253: out std_logic;
		G6254: out std_logic;
		G6255: out std_logic;
		G6256: out std_logic;
		G6257: out std_logic;
		G6258: out std_logic;
		G6259: out std_logic;
		G6260: out std_logic;
		G6261: out std_logic;
		G6262: out std_logic;
		G6263: out std_logic;
		G6264: out std_logic;
		G6265: out std_logic;
		G6266: out std_logic;
		G6267: out std_logic;
		G6268: out std_logic;
		G6269: out std_logic;
		G6270: out std_logic;
		G6271: out std_logic;
		G6272: out std_logic;
		G6273: out std_logic;
		G6274: out std_logic;
		G6275: out std_logic;
		G6276: out std_logic;
		G6277: out std_logic;
		G6278: out std_logic;
		G6279: out std_logic;
		G6280: out std_logic;
		G6281: out std_logic;
		G6282: out std_logic;
		G6283: out std_logic;
		G6284: out std_logic;
		G6285: out std_logic;
		G6842: out std_logic;
		G6920: out std_logic;
		G6926: out std_logic;
		G6932: out std_logic;
		G6942: out std_logic;
		G6949: out std_logic;
		G6955: out std_logic;
		G7744: out std_logic;
		G8061: out std_logic;
		G8062: out std_logic;
		G8271: out std_logic;
		G8313: out std_logic;
		G8316: out std_logic;
		G8318: out std_logic;
		G8323: out std_logic;
		G8328: out std_logic;
		G8331: out std_logic;
		G8335: out std_logic;
		G8340: out std_logic;
		G8347: out std_logic;
		G8349: out std_logic;
		G8352: out std_logic;
		G8561: out std_logic;
		G8562: out std_logic;
		G8563: out std_logic;
		G8564: out std_logic;
		G8565: out std_logic;
		G8566: out std_logic;
		G8976: out std_logic;
		G8977: out std_logic;
		G8978: out std_logic;
		G8979: out std_logic;
		G8980: out std_logic;
		G8981: out std_logic;
		G8982: out std_logic;
		G8983: out std_logic;
		G8984: out std_logic;
		G8985: out std_logic;
		G8986: out std_logic;
		G9451: out std_logic;
		G9961: out std_logic;
		G10377: out std_logic;
		G10379: out std_logic;
		G10455: out std_logic;
		G10457: out std_logic;
		G10459: out std_logic;
		G10461: out std_logic;
		G10463: out std_logic;
		G10465: out std_logic;
		G10628: out std_logic;
		G10801: out std_logic;
		G11163: out std_logic;
		G11206: out std_logic;
		G11489: out std_logic
	);
end entity;

architecture RTL of s15850 is
	attribute dont_touch: boolean;

	signal G1: std_logic; attribute dont_touch of G1: signal is true;
	signal G4: std_logic; attribute dont_touch of G4: signal is true;
	signal G7: std_logic; attribute dont_touch of G7: signal is true;
	signal G8: std_logic; attribute dont_touch of G8: signal is true;
	signal G9: std_logic; attribute dont_touch of G9: signal is true;
	signal G12: std_logic; attribute dont_touch of G12: signal is true;
	signal G16: std_logic; attribute dont_touch of G16: signal is true;
	signal G17: std_logic; attribute dont_touch of G17: signal is true;
	signal G22: std_logic; attribute dont_touch of G22: signal is true;
	signal G26: std_logic; attribute dont_touch of G26: signal is true;
	signal G32: std_logic; attribute dont_touch of G32: signal is true;
	signal G33: std_logic; attribute dont_touch of G33: signal is true;
	signal G34: std_logic; attribute dont_touch of G34: signal is true;
	signal G35: std_logic; attribute dont_touch of G35: signal is true;
	signal G36: std_logic; attribute dont_touch of G36: signal is true;
	signal G37: std_logic; attribute dont_touch of G37: signal is true;
	signal G38: std_logic; attribute dont_touch of G38: signal is true;
	signal G39: std_logic; attribute dont_touch of G39: signal is true;
	signal G40: std_logic; attribute dont_touch of G40: signal is true;
	signal G49: std_logic; attribute dont_touch of G49: signal is true;
	signal G52: std_logic; attribute dont_touch of G52: signal is true;
	signal G55: std_logic; attribute dont_touch of G55: signal is true;
	signal G58: std_logic; attribute dont_touch of G58: signal is true;
	signal G61: std_logic; attribute dont_touch of G61: signal is true;
	signal G64: std_logic; attribute dont_touch of G64: signal is true;
	signal G67: std_logic; attribute dont_touch of G67: signal is true;
	signal G70: std_logic; attribute dont_touch of G70: signal is true;
	signal G73: std_logic; attribute dont_touch of G73: signal is true;
	signal G76: std_logic; attribute dont_touch of G76: signal is true;
	signal G79: std_logic; attribute dont_touch of G79: signal is true;
	signal G97: std_logic; attribute dont_touch of G97: signal is true;
	signal G98: std_logic; attribute dont_touch of G98: signal is true;
	signal G105: std_logic; attribute dont_touch of G105: signal is true;
	signal G108: std_logic; attribute dont_touch of G108: signal is true;
	signal G110: std_logic; attribute dont_touch of G110: signal is true;
	signal G113: std_logic; attribute dont_touch of G113: signal is true;
	signal G114: std_logic; attribute dont_touch of G114: signal is true;
	signal G115: std_logic; attribute dont_touch of G115: signal is true;
	signal G119: std_logic; attribute dont_touch of G119: signal is true;
	signal G123: std_logic; attribute dont_touch of G123: signal is true;
	signal G126: std_logic; attribute dont_touch of G126: signal is true;
	signal G127: std_logic; attribute dont_touch of G127: signal is true;
	signal G131: std_logic; attribute dont_touch of G131: signal is true;
	signal G135: std_logic; attribute dont_touch of G135: signal is true;
	signal G139: std_logic; attribute dont_touch of G139: signal is true;
	signal G143: std_logic; attribute dont_touch of G143: signal is true;
	signal G148: std_logic; attribute dont_touch of G148: signal is true;
	signal G153: std_logic; attribute dont_touch of G153: signal is true;
	signal G158: std_logic; attribute dont_touch of G158: signal is true;
	signal G162: std_logic; attribute dont_touch of G162: signal is true;
	signal G166: std_logic; attribute dont_touch of G166: signal is true;
	signal G170: std_logic; attribute dont_touch of G170: signal is true;
	signal G174: std_logic; attribute dont_touch of G174: signal is true;
	signal G178: std_logic; attribute dont_touch of G178: signal is true;
	signal G182: std_logic; attribute dont_touch of G182: signal is true;
	signal G186: std_logic; attribute dont_touch of G186: signal is true;
	signal G192: std_logic; attribute dont_touch of G192: signal is true;
	signal G197: std_logic; attribute dont_touch of G197: signal is true;
	signal G201: std_logic; attribute dont_touch of G201: signal is true;
	signal G207: std_logic; attribute dont_touch of G207: signal is true;
	signal G213: std_logic; attribute dont_touch of G213: signal is true;
	signal G219: std_logic; attribute dont_touch of G219: signal is true;
	signal G225: std_logic; attribute dont_touch of G225: signal is true;
	signal G231: std_logic; attribute dont_touch of G231: signal is true;
	signal G237: std_logic; attribute dont_touch of G237: signal is true;
	signal G243: std_logic; attribute dont_touch of G243: signal is true;
	signal G248: std_logic; attribute dont_touch of G248: signal is true;
	signal G253: std_logic; attribute dont_touch of G253: signal is true;
	signal G254: std_logic; attribute dont_touch of G254: signal is true;
	signal G255: std_logic; attribute dont_touch of G255: signal is true;
	signal G256: std_logic; attribute dont_touch of G256: signal is true;
	signal G257: std_logic; attribute dont_touch of G257: signal is true;
	signal G258: std_logic; attribute dont_touch of G258: signal is true;
	signal G259: std_logic; attribute dont_touch of G259: signal is true;
	signal G260: std_logic; attribute dont_touch of G260: signal is true;
	signal G261: std_logic; attribute dont_touch of G261: signal is true;
	signal G262: std_logic; attribute dont_touch of G262: signal is true;
	signal G263: std_logic; attribute dont_touch of G263: signal is true;
	signal G266: std_logic; attribute dont_touch of G266: signal is true;
	signal G269: std_logic; attribute dont_touch of G269: signal is true;
	signal G272: std_logic; attribute dont_touch of G272: signal is true;
	signal G275: std_logic; attribute dont_touch of G275: signal is true;
	signal G278: std_logic; attribute dont_touch of G278: signal is true;
	signal G281: std_logic; attribute dont_touch of G281: signal is true;
	signal G284: std_logic; attribute dont_touch of G284: signal is true;
	signal G287: std_logic; attribute dont_touch of G287: signal is true;
	signal G290: std_logic; attribute dont_touch of G290: signal is true;
	signal G293: std_logic; attribute dont_touch of G293: signal is true;
	signal G296: std_logic; attribute dont_touch of G296: signal is true;
	signal G299: std_logic; attribute dont_touch of G299: signal is true;
	signal G302: std_logic; attribute dont_touch of G302: signal is true;
	signal G305: std_logic; attribute dont_touch of G305: signal is true;
	signal G309: std_logic; attribute dont_touch of G309: signal is true;
	signal G312: std_logic; attribute dont_touch of G312: signal is true;
	signal G315: std_logic; attribute dont_touch of G315: signal is true;
	signal G318: std_logic; attribute dont_touch of G318: signal is true;
	signal G321: std_logic; attribute dont_touch of G321: signal is true;
	signal G324: std_logic; attribute dont_touch of G324: signal is true;
	signal G327: std_logic; attribute dont_touch of G327: signal is true;
	signal G330: std_logic; attribute dont_touch of G330: signal is true;
	signal G333: std_logic; attribute dont_touch of G333: signal is true;
	signal G336: std_logic; attribute dont_touch of G336: signal is true;
	signal G339: std_logic; attribute dont_touch of G339: signal is true;
	signal G342: std_logic; attribute dont_touch of G342: signal is true;
	signal G345: std_logic; attribute dont_touch of G345: signal is true;
	signal G348: std_logic; attribute dont_touch of G348: signal is true;
	signal G351: std_logic; attribute dont_touch of G351: signal is true;
	signal G354: std_logic; attribute dont_touch of G354: signal is true;
	signal G357: std_logic; attribute dont_touch of G357: signal is true;
	signal G360: std_logic; attribute dont_touch of G360: signal is true;
	signal G363: std_logic; attribute dont_touch of G363: signal is true;
	signal G366: std_logic; attribute dont_touch of G366: signal is true;
	signal G369: std_logic; attribute dont_touch of G369: signal is true;
	signal G374: std_logic; attribute dont_touch of G374: signal is true;
	signal G378: std_logic; attribute dont_touch of G378: signal is true;
	signal G382: std_logic; attribute dont_touch of G382: signal is true;
	signal G386: std_logic; attribute dont_touch of G386: signal is true;
	signal G391: std_logic; attribute dont_touch of G391: signal is true;
	signal G396: std_logic; attribute dont_touch of G396: signal is true;
	signal G401: std_logic; attribute dont_touch of G401: signal is true;
	signal G406: std_logic; attribute dont_touch of G406: signal is true;
	signal G411: std_logic; attribute dont_touch of G411: signal is true;
	signal G416: std_logic; attribute dont_touch of G416: signal is true;
	signal G421: std_logic; attribute dont_touch of G421: signal is true;
	signal G426: std_logic; attribute dont_touch of G426: signal is true;
	signal G431: std_logic; attribute dont_touch of G431: signal is true;
	signal G435: std_logic; attribute dont_touch of G435: signal is true;
	signal G440: std_logic; attribute dont_touch of G440: signal is true;
	signal G444: std_logic; attribute dont_touch of G444: signal is true;
	signal G448: std_logic; attribute dont_touch of G448: signal is true;
	signal G452: std_logic; attribute dont_touch of G452: signal is true;
	signal G456: std_logic; attribute dont_touch of G456: signal is true;
	signal G461: std_logic; attribute dont_touch of G461: signal is true;
	signal G466: std_logic; attribute dont_touch of G466: signal is true;
	signal G471: std_logic; attribute dont_touch of G471: signal is true;
	signal G476: std_logic; attribute dont_touch of G476: signal is true;
	signal G481: std_logic; attribute dont_touch of G481: signal is true;
	signal G486: std_logic; attribute dont_touch of G486: signal is true;
	signal G491: std_logic; attribute dont_touch of G491: signal is true;
	signal G496: std_logic; attribute dont_touch of G496: signal is true;
	signal G501: std_logic; attribute dont_touch of G501: signal is true;
	signal G506: std_logic; attribute dont_touch of G506: signal is true;
	signal G511: std_logic; attribute dont_touch of G511: signal is true;
	signal G516: std_logic; attribute dont_touch of G516: signal is true;
	signal G521: std_logic; attribute dont_touch of G521: signal is true;
	signal G525: std_logic; attribute dont_touch of G525: signal is true;
	signal G530: std_logic; attribute dont_touch of G530: signal is true;
	signal G534: std_logic; attribute dont_touch of G534: signal is true;
	signal G538: std_logic; attribute dont_touch of G538: signal is true;
	signal G542: std_logic; attribute dont_touch of G542: signal is true;
	signal G546: std_logic; attribute dont_touch of G546: signal is true;
	signal G549: std_logic; attribute dont_touch of G549: signal is true;
	signal G552: std_logic; attribute dont_touch of G552: signal is true;
	signal G553: std_logic; attribute dont_touch of G553: signal is true;
	signal G554: std_logic; attribute dont_touch of G554: signal is true;
	signal G557: std_logic; attribute dont_touch of G557: signal is true;
	signal G560: std_logic; attribute dont_touch of G560: signal is true;
	signal G563: std_logic; attribute dont_touch of G563: signal is true;
	signal G566: std_logic; attribute dont_touch of G566: signal is true;
	signal G569: std_logic; attribute dont_touch of G569: signal is true;
	signal G572: std_logic; attribute dont_touch of G572: signal is true;
	signal G575: std_logic; attribute dont_touch of G575: signal is true;
	signal G578: std_logic; attribute dont_touch of G578: signal is true;
	signal G579: std_logic; attribute dont_touch of G579: signal is true;
	signal G580: std_logic; attribute dont_touch of G580: signal is true;
	signal G581: std_logic; attribute dont_touch of G581: signal is true;
	signal G582: std_logic; attribute dont_touch of G582: signal is true;
	signal G583: std_logic; attribute dont_touch of G583: signal is true;
	signal G584: std_logic; attribute dont_touch of G584: signal is true;
	signal G585: std_logic; attribute dont_touch of G585: signal is true;
	signal G586: std_logic; attribute dont_touch of G586: signal is true;
	signal G587: std_logic; attribute dont_touch of G587: signal is true;
	signal G588: std_logic; attribute dont_touch of G588: signal is true;
	signal G589: std_logic; attribute dont_touch of G589: signal is true;
	signal G590: std_logic; attribute dont_touch of G590: signal is true;
	signal G591: std_logic; attribute dont_touch of G591: signal is true;
	signal G599: std_logic; attribute dont_touch of G599: signal is true;
	signal G605: std_logic; attribute dont_touch of G605: signal is true;
	signal G611: std_logic; attribute dont_touch of G611: signal is true;
	signal G617: std_logic; attribute dont_touch of G617: signal is true;
	signal G622: std_logic; attribute dont_touch of G622: signal is true;
	signal G627: std_logic; attribute dont_touch of G627: signal is true;
	signal G630: std_logic; attribute dont_touch of G630: signal is true;
	signal G631: std_logic; attribute dont_touch of G631: signal is true;
	signal G632: std_logic; attribute dont_touch of G632: signal is true;
	signal G635: std_logic; attribute dont_touch of G635: signal is true;
	signal G636: std_logic; attribute dont_touch of G636: signal is true;
	signal G639: std_logic; attribute dont_touch of G639: signal is true;
	signal G643: std_logic; attribute dont_touch of G643: signal is true;
	signal G646: std_logic; attribute dont_touch of G646: signal is true;
	signal G650: std_logic; attribute dont_touch of G650: signal is true;
	signal G654: std_logic; attribute dont_touch of G654: signal is true;
	signal G658: std_logic; attribute dont_touch of G658: signal is true;
	signal G664: std_logic; attribute dont_touch of G664: signal is true;
	signal G668: std_logic; attribute dont_touch of G668: signal is true;
	signal G673: std_logic; attribute dont_touch of G673: signal is true;
	signal G677: std_logic; attribute dont_touch of G677: signal is true;
	signal G682: std_logic; attribute dont_touch of G682: signal is true;
	signal G686: std_logic; attribute dont_touch of G686: signal is true;
	signal G691: std_logic; attribute dont_touch of G691: signal is true;
	signal G695: std_logic; attribute dont_touch of G695: signal is true;
	signal G700: std_logic; attribute dont_touch of G700: signal is true;
	signal G704: std_logic; attribute dont_touch of G704: signal is true;
	signal G709: std_logic; attribute dont_touch of G709: signal is true;
	signal G713: std_logic; attribute dont_touch of G713: signal is true;
	signal G718: std_logic; attribute dont_touch of G718: signal is true;
	signal G722: std_logic; attribute dont_touch of G722: signal is true;
	signal G727: std_logic; attribute dont_touch of G727: signal is true;
	signal G731: std_logic; attribute dont_touch of G731: signal is true;
	signal G736: std_logic; attribute dont_touch of G736: signal is true;
	signal G745: std_logic; attribute dont_touch of G745: signal is true;
	signal G746: std_logic; attribute dont_touch of G746: signal is true;
	signal G754: std_logic; attribute dont_touch of G754: signal is true;
	signal G755: std_logic; attribute dont_touch of G755: signal is true;
	signal G756: std_logic; attribute dont_touch of G756: signal is true;
	signal G757: std_logic; attribute dont_touch of G757: signal is true;
	signal G758: std_logic; attribute dont_touch of G758: signal is true;
	signal G762: std_logic; attribute dont_touch of G762: signal is true;
	signal G766: std_logic; attribute dont_touch of G766: signal is true;
	signal G770: std_logic; attribute dont_touch of G770: signal is true;
	signal G774: std_logic; attribute dont_touch of G774: signal is true;
	signal G778: std_logic; attribute dont_touch of G778: signal is true;
	signal G782: std_logic; attribute dont_touch of G782: signal is true;
	signal G786: std_logic; attribute dont_touch of G786: signal is true;
	signal G790: std_logic; attribute dont_touch of G790: signal is true;
	signal G794: std_logic; attribute dont_touch of G794: signal is true;
	signal G798: std_logic; attribute dont_touch of G798: signal is true;
	signal G802: std_logic; attribute dont_touch of G802: signal is true;
	signal G806: std_logic; attribute dont_touch of G806: signal is true;
	signal G810: std_logic; attribute dont_touch of G810: signal is true;
	signal G814: std_logic; attribute dont_touch of G814: signal is true;
	signal G818: std_logic; attribute dont_touch of G818: signal is true;
	signal G822: std_logic; attribute dont_touch of G822: signal is true;
	signal G826: std_logic; attribute dont_touch of G826: signal is true;
	signal G829: std_logic; attribute dont_touch of G829: signal is true;
	signal G833: std_logic; attribute dont_touch of G833: signal is true;
	signal G837: std_logic; attribute dont_touch of G837: signal is true;
	signal G841: std_logic; attribute dont_touch of G841: signal is true;
	signal G845: std_logic; attribute dont_touch of G845: signal is true;
	signal G849: std_logic; attribute dont_touch of G849: signal is true;
	signal G853: std_logic; attribute dont_touch of G853: signal is true;
	signal G857: std_logic; attribute dont_touch of G857: signal is true;
	signal G861: std_logic; attribute dont_touch of G861: signal is true;
	signal G865: std_logic; attribute dont_touch of G865: signal is true;
	signal G868: std_logic; attribute dont_touch of G868: signal is true;
	signal G869: std_logic; attribute dont_touch of G869: signal is true;
	signal G874: std_logic; attribute dont_touch of G874: signal is true;
	signal G875: std_logic; attribute dont_touch of G875: signal is true;
	signal G876: std_logic; attribute dont_touch of G876: signal is true;
	signal G878: std_logic; attribute dont_touch of G878: signal is true;
	signal G882: std_logic; attribute dont_touch of G882: signal is true;
	signal G883: std_logic; attribute dont_touch of G883: signal is true;
	signal G928: std_logic; attribute dont_touch of G928: signal is true;
	signal G932: std_logic; attribute dont_touch of G932: signal is true;
	signal G936: std_logic; attribute dont_touch of G936: signal is true;
	signal G940: std_logic; attribute dont_touch of G940: signal is true;
	signal G944: std_logic; attribute dont_touch of G944: signal is true;
	signal G947: std_logic; attribute dont_touch of G947: signal is true;
	signal G950: std_logic; attribute dont_touch of G950: signal is true;
	signal G953: std_logic; attribute dont_touch of G953: signal is true;
	signal G956: std_logic; attribute dont_touch of G956: signal is true;
	signal G959: std_logic; attribute dont_touch of G959: signal is true;
	signal G962: std_logic; attribute dont_touch of G962: signal is true;
	signal G965: std_logic; attribute dont_touch of G965: signal is true;
	signal G968: std_logic; attribute dont_touch of G968: signal is true;
	signal G971: std_logic; attribute dont_touch of G971: signal is true;
	signal G976: std_logic; attribute dont_touch of G976: signal is true;
	signal G981: std_logic; attribute dont_touch of G981: signal is true;
	signal G986: std_logic; attribute dont_touch of G986: signal is true;
	signal G991: std_logic; attribute dont_touch of G991: signal is true;
	signal G995: std_logic; attribute dont_touch of G995: signal is true;
	signal G999: std_logic; attribute dont_touch of G999: signal is true;
	signal G1003: std_logic; attribute dont_touch of G1003: signal is true;
	signal G1007: std_logic; attribute dont_touch of G1007: signal is true;
	signal G1011: std_logic; attribute dont_touch of G1011: signal is true;
	signal G1015: std_logic; attribute dont_touch of G1015: signal is true;
	signal G1019: std_logic; attribute dont_touch of G1019: signal is true;
	signal G1023: std_logic; attribute dont_touch of G1023: signal is true;
	signal G1027: std_logic; attribute dont_touch of G1027: signal is true;
	signal G1032: std_logic; attribute dont_touch of G1032: signal is true;
	signal G1035: std_logic; attribute dont_touch of G1035: signal is true;
	signal G1038: std_logic; attribute dont_touch of G1038: signal is true;
	signal G1041: std_logic; attribute dont_touch of G1041: signal is true;
	signal G1044: std_logic; attribute dont_touch of G1044: signal is true;
	signal G1047: std_logic; attribute dont_touch of G1047: signal is true;
	signal G1050: std_logic; attribute dont_touch of G1050: signal is true;
	signal G1053: std_logic; attribute dont_touch of G1053: signal is true;
	signal G1056: std_logic; attribute dont_touch of G1056: signal is true;
	signal G1059: std_logic; attribute dont_touch of G1059: signal is true;
	signal G1062: std_logic; attribute dont_touch of G1062: signal is true;
	signal G1065: std_logic; attribute dont_touch of G1065: signal is true;
	signal G1068: std_logic; attribute dont_touch of G1068: signal is true;
	signal G1071: std_logic; attribute dont_touch of G1071: signal is true;
	signal G1074: std_logic; attribute dont_touch of G1074: signal is true;
	signal G1077: std_logic; attribute dont_touch of G1077: signal is true;
	signal G1080: std_logic; attribute dont_touch of G1080: signal is true;
	signal G1083: std_logic; attribute dont_touch of G1083: signal is true;
	signal G1086: std_logic; attribute dont_touch of G1086: signal is true;
	signal G1089: std_logic; attribute dont_touch of G1089: signal is true;
	signal G1092: std_logic; attribute dont_touch of G1092: signal is true;
	signal G1095: std_logic; attribute dont_touch of G1095: signal is true;
	signal G1098: std_logic; attribute dont_touch of G1098: signal is true;
	signal G1101: std_logic; attribute dont_touch of G1101: signal is true;
	signal G1104: std_logic; attribute dont_touch of G1104: signal is true;
	signal G1107: std_logic; attribute dont_touch of G1107: signal is true;
	signal G1110: std_logic; attribute dont_touch of G1110: signal is true;
	signal G1113: std_logic; attribute dont_touch of G1113: signal is true;
	signal G1117: std_logic; attribute dont_touch of G1117: signal is true;
	signal G1121: std_logic; attribute dont_touch of G1121: signal is true;
	signal G1125: std_logic; attribute dont_touch of G1125: signal is true;
	signal G1129: std_logic; attribute dont_touch of G1129: signal is true;
	signal G1133: std_logic; attribute dont_touch of G1133: signal is true;
	signal G1137: std_logic; attribute dont_touch of G1137: signal is true;
	signal G1141: std_logic; attribute dont_touch of G1141: signal is true;
	signal G1145: std_logic; attribute dont_touch of G1145: signal is true;
	signal G1149: std_logic; attribute dont_touch of G1149: signal is true;
	signal G1153: std_logic; attribute dont_touch of G1153: signal is true;
	signal G1157: std_logic; attribute dont_touch of G1157: signal is true;
	signal G1160: std_logic; attribute dont_touch of G1160: signal is true;
	signal G1163: std_logic; attribute dont_touch of G1163: signal is true;
	signal G1166: std_logic; attribute dont_touch of G1166: signal is true;
	signal G1169: std_logic; attribute dont_touch of G1169: signal is true;
	signal G1206: std_logic; attribute dont_touch of G1206: signal is true;
	signal G1209: std_logic; attribute dont_touch of G1209: signal is true;
	signal G1212: std_logic; attribute dont_touch of G1212: signal is true;
	signal G1215: std_logic; attribute dont_touch of G1215: signal is true;
	signal G1216: std_logic; attribute dont_touch of G1216: signal is true;
	signal G1217: std_logic; attribute dont_touch of G1217: signal is true;
	signal G1218: std_logic; attribute dont_touch of G1218: signal is true;
	signal G1223: std_logic; attribute dont_touch of G1223: signal is true;
	signal G1227: std_logic; attribute dont_touch of G1227: signal is true;
	signal G1231: std_logic; attribute dont_touch of G1231: signal is true;
	signal G1235: std_logic; attribute dont_touch of G1235: signal is true;
	signal G1240: std_logic; attribute dont_touch of G1240: signal is true;
	signal G1245: std_logic; attribute dont_touch of G1245: signal is true;
	signal G1250: std_logic; attribute dont_touch of G1250: signal is true;
	signal G1255: std_logic; attribute dont_touch of G1255: signal is true;
	signal G1260: std_logic; attribute dont_touch of G1260: signal is true;
	signal G1265: std_logic; attribute dont_touch of G1265: signal is true;
	signal G1270: std_logic; attribute dont_touch of G1270: signal is true;
	signal G1275: std_logic; attribute dont_touch of G1275: signal is true;
	signal G1280: std_logic; attribute dont_touch of G1280: signal is true;
	signal G1284: std_logic; attribute dont_touch of G1284: signal is true;
	signal G1289: std_logic; attribute dont_touch of G1289: signal is true;
	signal G1292: std_logic; attribute dont_touch of G1292: signal is true;
	signal G1296: std_logic; attribute dont_touch of G1296: signal is true;
	signal G1300: std_logic; attribute dont_touch of G1300: signal is true;
	signal G1304: std_logic; attribute dont_touch of G1304: signal is true;
	signal G1308: std_logic; attribute dont_touch of G1308: signal is true;
	signal G1311: std_logic; attribute dont_touch of G1311: signal is true;
	signal G1314: std_logic; attribute dont_touch of G1314: signal is true;
	signal G1317: std_logic; attribute dont_touch of G1317: signal is true;
	signal G1318: std_logic; attribute dont_touch of G1318: signal is true;
	signal G1321: std_logic; attribute dont_touch of G1321: signal is true;
	signal G1324: std_logic; attribute dont_touch of G1324: signal is true;
	signal G1327: std_logic; attribute dont_touch of G1327: signal is true;
	signal G1330: std_logic; attribute dont_touch of G1330: signal is true;
	signal G1333: std_logic; attribute dont_touch of G1333: signal is true;
	signal G1336: std_logic; attribute dont_touch of G1336: signal is true;
	signal G1341: std_logic; attribute dont_touch of G1341: signal is true;
	signal G1346: std_logic; attribute dont_touch of G1346: signal is true;
	signal G1351: std_logic; attribute dont_touch of G1351: signal is true;
	signal G1356: std_logic; attribute dont_touch of G1356: signal is true;
	signal G1357: std_logic; attribute dont_touch of G1357: signal is true;
	signal G1360: std_logic; attribute dont_touch of G1360: signal is true;
	signal G1361: std_logic; attribute dont_touch of G1361: signal is true;
	signal G1362: std_logic; attribute dont_touch of G1362: signal is true;
	signal G1365: std_logic; attribute dont_touch of G1365: signal is true;
	signal G1368: std_logic; attribute dont_touch of G1368: signal is true;
	signal G1371: std_logic; attribute dont_touch of G1371: signal is true;
	signal G1374: std_logic; attribute dont_touch of G1374: signal is true;
	signal G1377: std_logic; attribute dont_touch of G1377: signal is true;
	signal G1380: std_logic; attribute dont_touch of G1380: signal is true;
	signal G1383: std_logic; attribute dont_touch of G1383: signal is true;
	signal G1386: std_logic; attribute dont_touch of G1386: signal is true;
	signal G1389: std_logic; attribute dont_touch of G1389: signal is true;
	signal G1393: std_logic; attribute dont_touch of G1393: signal is true;
	signal G1394: std_logic; attribute dont_touch of G1394: signal is true;
	signal G1397: std_logic; attribute dont_touch of G1397: signal is true;
	signal G1400: std_logic; attribute dont_touch of G1400: signal is true;
	signal G1403: std_logic; attribute dont_touch of G1403: signal is true;
	signal G1407: std_logic; attribute dont_touch of G1407: signal is true;
	signal G1411: std_logic; attribute dont_touch of G1411: signal is true;
	signal G1415: std_logic; attribute dont_touch of G1415: signal is true;
	signal G1419: std_logic; attribute dont_touch of G1419: signal is true;
	signal G1424: std_logic; attribute dont_touch of G1424: signal is true;
	signal G1428: std_logic; attribute dont_touch of G1428: signal is true;
	signal G1432: std_logic; attribute dont_touch of G1432: signal is true;
	signal G1436: std_logic; attribute dont_touch of G1436: signal is true;
	signal G1440: std_logic; attribute dont_touch of G1440: signal is true;
	signal G1444: std_logic; attribute dont_touch of G1444: signal is true;
	signal G1448: std_logic; attribute dont_touch of G1448: signal is true;
	signal G1453: std_logic; attribute dont_touch of G1453: signal is true;
	signal G1458: std_logic; attribute dont_touch of G1458: signal is true;
	signal G1462: std_logic; attribute dont_touch of G1462: signal is true;
	signal G1466: std_logic; attribute dont_touch of G1466: signal is true;
	signal G1470: std_logic; attribute dont_touch of G1470: signal is true;
	signal G1474: std_logic; attribute dont_touch of G1474: signal is true;
	signal G1478: std_logic; attribute dont_touch of G1478: signal is true;
	signal G1482: std_logic; attribute dont_touch of G1482: signal is true;
	signal G1486: std_logic; attribute dont_touch of G1486: signal is true;
	signal G1490: std_logic; attribute dont_touch of G1490: signal is true;
	signal G1494: std_logic; attribute dont_touch of G1494: signal is true;
	signal G1499: std_logic; attribute dont_touch of G1499: signal is true;
	signal G1504: std_logic; attribute dont_touch of G1504: signal is true;
	signal G1508: std_logic; attribute dont_touch of G1508: signal is true;
	signal G1512: std_logic; attribute dont_touch of G1512: signal is true;
	signal G1515: std_logic; attribute dont_touch of G1515: signal is true;
	signal G1520: std_logic; attribute dont_touch of G1520: signal is true;
	signal G1524: std_logic; attribute dont_touch of G1524: signal is true;
	signal G1527: std_logic; attribute dont_touch of G1527: signal is true;
	signal G1528: std_logic; attribute dont_touch of G1528: signal is true;
	signal G1531: std_logic; attribute dont_touch of G1531: signal is true;
	signal G1534: std_logic; attribute dont_touch of G1534: signal is true;
	signal G1537: std_logic; attribute dont_touch of G1537: signal is true;
	signal G1540: std_logic; attribute dont_touch of G1540: signal is true;
	signal G1543: std_logic; attribute dont_touch of G1543: signal is true;
	signal G1546: std_logic; attribute dont_touch of G1546: signal is true;
	signal G1549: std_logic; attribute dont_touch of G1549: signal is true;
	signal G1552: std_logic; attribute dont_touch of G1552: signal is true;
	signal G1555: std_logic; attribute dont_touch of G1555: signal is true;
	signal G1558: std_logic; attribute dont_touch of G1558: signal is true;
	signal G1561: std_logic; attribute dont_touch of G1561: signal is true;
	signal G1564: std_logic; attribute dont_touch of G1564: signal is true;
	signal G1567: std_logic; attribute dont_touch of G1567: signal is true;
	signal G1570: std_logic; attribute dont_touch of G1570: signal is true;
	signal G1571: std_logic; attribute dont_touch of G1571: signal is true;
	signal G1574: std_logic; attribute dont_touch of G1574: signal is true;
	signal G1577: std_logic; attribute dont_touch of G1577: signal is true;
	signal G1580: std_logic; attribute dont_touch of G1580: signal is true;
	signal G1583: std_logic; attribute dont_touch of G1583: signal is true;
	signal G1586: std_logic; attribute dont_touch of G1586: signal is true;
	signal G1589: std_logic; attribute dont_touch of G1589: signal is true;
	signal G1592: std_logic; attribute dont_touch of G1592: signal is true;
	signal G1595: std_logic; attribute dont_touch of G1595: signal is true;
	signal G1598: std_logic; attribute dont_touch of G1598: signal is true;
	signal G1601: std_logic; attribute dont_touch of G1601: signal is true;
	signal G1604: std_logic; attribute dont_touch of G1604: signal is true;
	signal G1607: std_logic; attribute dont_touch of G1607: signal is true;
	signal G1610: std_logic; attribute dont_touch of G1610: signal is true;
	signal G1615: std_logic; attribute dont_touch of G1615: signal is true;
	signal G1618: std_logic; attribute dont_touch of G1618: signal is true;
	signal G1621: std_logic; attribute dont_touch of G1621: signal is true;
	signal G1624: std_logic; attribute dont_touch of G1624: signal is true;
	signal G1627: std_logic; attribute dont_touch of G1627: signal is true;
	signal G1630: std_logic; attribute dont_touch of G1630: signal is true;
	signal G1633: std_logic; attribute dont_touch of G1633: signal is true;
	signal G1636: std_logic; attribute dont_touch of G1636: signal is true;
	signal G1639: std_logic; attribute dont_touch of G1639: signal is true;
	signal G1642: std_logic; attribute dont_touch of G1642: signal is true;
	signal G1645: std_logic; attribute dont_touch of G1645: signal is true;
	signal G1648: std_logic; attribute dont_touch of G1648: signal is true;
	signal G1651: std_logic; attribute dont_touch of G1651: signal is true;
	signal G1654: std_logic; attribute dont_touch of G1654: signal is true;
	signal G1657: std_logic; attribute dont_touch of G1657: signal is true;
	signal G1660: std_logic; attribute dont_touch of G1660: signal is true;
	signal G1663: std_logic; attribute dont_touch of G1663: signal is true;
	signal G1666: std_logic; attribute dont_touch of G1666: signal is true;
	signal G1669: std_logic; attribute dont_touch of G1669: signal is true;
	signal G1672: std_logic; attribute dont_touch of G1672: signal is true;
	signal G1675: std_logic; attribute dont_touch of G1675: signal is true;
	signal G1678: std_logic; attribute dont_touch of G1678: signal is true;
	signal G1681: std_logic; attribute dont_touch of G1681: signal is true;
	signal G1684: std_logic; attribute dont_touch of G1684: signal is true;
	signal G1687: std_logic; attribute dont_touch of G1687: signal is true;
	signal G1690: std_logic; attribute dont_touch of G1690: signal is true;
	signal G1703: std_logic; attribute dont_touch of G1703: signal is true;
	signal G1707: std_logic; attribute dont_touch of G1707: signal is true;
	signal G1710: std_logic; attribute dont_touch of G1710: signal is true;
	signal G1711: std_logic; attribute dont_touch of G1711: signal is true;
	signal G1713: std_logic; attribute dont_touch of G1713: signal is true;
	signal G1718: std_logic; attribute dont_touch of G1718: signal is true;
	signal G1721: std_logic; attribute dont_touch of G1721: signal is true;
	signal G1724: std_logic; attribute dont_touch of G1724: signal is true;
	signal G1727: std_logic; attribute dont_touch of G1727: signal is true;
	signal G1730: std_logic; attribute dont_touch of G1730: signal is true;
	signal G1733: std_logic; attribute dont_touch of G1733: signal is true;
	signal G1736: std_logic; attribute dont_touch of G1736: signal is true;
	signal G1737: std_logic; attribute dont_touch of G1737: signal is true;
	signal G1738: std_logic; attribute dont_touch of G1738: signal is true;
	signal G1741: std_logic; attribute dont_touch of G1741: signal is true;
	signal G1744: std_logic; attribute dont_touch of G1744: signal is true;
	signal G1747: std_logic; attribute dont_touch of G1747: signal is true;
	signal G1750: std_logic; attribute dont_touch of G1750: signal is true;
	signal G1753: std_logic; attribute dont_touch of G1753: signal is true;
	signal G1756: std_logic; attribute dont_touch of G1756: signal is true;
	signal G1759: std_logic; attribute dont_touch of G1759: signal is true;
	signal G1762: std_logic; attribute dont_touch of G1762: signal is true;
	signal G1765: std_logic; attribute dont_touch of G1765: signal is true;
	signal G1766: std_logic; attribute dont_touch of G1766: signal is true;
	signal G1771: std_logic; attribute dont_touch of G1771: signal is true;
	signal G1776: std_logic; attribute dont_touch of G1776: signal is true;
	signal G1781: std_logic; attribute dont_touch of G1781: signal is true;
	signal G1786: std_logic; attribute dont_touch of G1786: signal is true;
	signal G1791: std_logic; attribute dont_touch of G1791: signal is true;
	signal G1796: std_logic; attribute dont_touch of G1796: signal is true;
	signal G1801: std_logic; attribute dont_touch of G1801: signal is true;
	signal G1806: std_logic; attribute dont_touch of G1806: signal is true;
	signal G1810: std_logic; attribute dont_touch of G1810: signal is true;
	signal G1811: std_logic; attribute dont_touch of G1811: signal is true;
	signal G1814: std_logic; attribute dont_touch of G1814: signal is true;
	signal G1822: std_logic; attribute dont_touch of G1822: signal is true;
	signal G1828: std_logic; attribute dont_touch of G1828: signal is true;
	signal G1834: std_logic; attribute dont_touch of G1834: signal is true;
	signal G1840: std_logic; attribute dont_touch of G1840: signal is true;
	signal G1845: std_logic; attribute dont_touch of G1845: signal is true;
	signal G1848: std_logic; attribute dont_touch of G1848: signal is true;
	signal G1849: std_logic; attribute dont_touch of G1849: signal is true;
	signal G1850: std_logic; attribute dont_touch of G1850: signal is true;
	signal G1853: std_logic; attribute dont_touch of G1853: signal is true;
	signal G1854: std_logic; attribute dont_touch of G1854: signal is true;
	signal G1857: std_logic; attribute dont_touch of G1857: signal is true;
	signal G1861: std_logic; attribute dont_touch of G1861: signal is true;
	signal G1864: std_logic; attribute dont_touch of G1864: signal is true;
	signal G1868: std_logic; attribute dont_touch of G1868: signal is true;
	signal G1872: std_logic; attribute dont_touch of G1872: signal is true;
	signal G1878: std_logic; attribute dont_touch of G1878: signal is true;
	signal G1882: std_logic; attribute dont_touch of G1882: signal is true;
	signal G1887: std_logic; attribute dont_touch of G1887: signal is true;
	signal G1891: std_logic; attribute dont_touch of G1891: signal is true;
	signal G1896: std_logic; attribute dont_touch of G1896: signal is true;
	signal G1900: std_logic; attribute dont_touch of G1900: signal is true;
	signal G1905: std_logic; attribute dont_touch of G1905: signal is true;
	signal G1909: std_logic; attribute dont_touch of G1909: signal is true;
	signal G1914: std_logic; attribute dont_touch of G1914: signal is true;
	signal G1918: std_logic; attribute dont_touch of G1918: signal is true;
	signal G1923: std_logic; attribute dont_touch of G1923: signal is true;
	signal G1927: std_logic; attribute dont_touch of G1927: signal is true;
	signal G1932: std_logic; attribute dont_touch of G1932: signal is true;
	signal G1936: std_logic; attribute dont_touch of G1936: signal is true;
	signal G1941: std_logic; attribute dont_touch of G1941: signal is true;
	signal G1945: std_logic; attribute dont_touch of G1945: signal is true;
	signal G1950: std_logic; attribute dont_touch of G1950: signal is true;
	signal G1955: std_logic; attribute dont_touch of G1955: signal is true;
	signal G1956: std_logic; attribute dont_touch of G1956: signal is true;
	signal G1958: std_logic; attribute dont_touch of G1958: signal is true;
	signal G1959: std_logic; attribute dont_touch of G1959: signal is true;
	signal G1962: std_logic; attribute dont_touch of G1962: signal is true;
	signal G1963: std_logic; attribute dont_touch of G1963: signal is true;
	signal G1964: std_logic; attribute dont_touch of G1964: signal is true;
	signal G1965: std_logic; attribute dont_touch of G1965: signal is true;
	signal G1968: std_logic; attribute dont_touch of G1968: signal is true;
	signal G1969: std_logic; attribute dont_touch of G1969: signal is true;
	signal G1972: std_logic; attribute dont_touch of G1972: signal is true;
	signal G1973: std_logic; attribute dont_touch of G1973: signal is true;
	signal G1974: std_logic; attribute dont_touch of G1974: signal is true;
	signal G1975: std_logic; attribute dont_touch of G1975: signal is true;
	signal G1976: std_logic; attribute dont_touch of G1976: signal is true;
	signal G1980: std_logic; attribute dont_touch of G1980: signal is true;
	signal G1981: std_logic; attribute dont_touch of G1981: signal is true;
	signal G1982: std_logic; attribute dont_touch of G1982: signal is true;
	signal G1983: std_logic; attribute dont_touch of G1983: signal is true;
	signal G1984: std_logic; attribute dont_touch of G1984: signal is true;
	signal G1987: std_logic; attribute dont_touch of G1987: signal is true;
	signal G1988: std_logic; attribute dont_touch of G1988: signal is true;
	signal G1989: std_logic; attribute dont_touch of G1989: signal is true;
	signal G1990: std_logic; attribute dont_touch of G1990: signal is true;
	signal G1991: std_logic; attribute dont_touch of G1991: signal is true;
	signal G1992: std_logic; attribute dont_touch of G1992: signal is true;
	signal G1993: std_logic; attribute dont_touch of G1993: signal is true;
	signal G1994: std_logic; attribute dont_touch of G1994: signal is true;
	signal G1997: std_logic; attribute dont_touch of G1997: signal is true;
	signal G1998: std_logic; attribute dont_touch of G1998: signal is true;
	signal G1999: std_logic; attribute dont_touch of G1999: signal is true;
	signal G2000: std_logic; attribute dont_touch of G2000: signal is true;
	signal G2001: std_logic; attribute dont_touch of G2001: signal is true;
	signal G2002: std_logic; attribute dont_touch of G2002: signal is true;
	signal G2003: std_logic; attribute dont_touch of G2003: signal is true;
	signal G2004: std_logic; attribute dont_touch of G2004: signal is true;
	signal G2005: std_logic; attribute dont_touch of G2005: signal is true;
	signal G2006: std_logic; attribute dont_touch of G2006: signal is true;
	signal G2007: std_logic; attribute dont_touch of G2007: signal is true;
	signal G2008: std_logic; attribute dont_touch of G2008: signal is true;
	signal G2011: std_logic; attribute dont_touch of G2011: signal is true;
	signal G2012: std_logic; attribute dont_touch of G2012: signal is true;
	signal G2013: std_logic; attribute dont_touch of G2013: signal is true;
	signal G2014: std_logic; attribute dont_touch of G2014: signal is true;
	signal G2015: std_logic; attribute dont_touch of G2015: signal is true;
	signal G2016: std_logic; attribute dont_touch of G2016: signal is true;
	signal G2017: std_logic; attribute dont_touch of G2017: signal is true;
	signal G2018: std_logic; attribute dont_touch of G2018: signal is true;
	signal G2021: std_logic; attribute dont_touch of G2021: signal is true;
	signal G2022: std_logic; attribute dont_touch of G2022: signal is true;
	signal G2023: std_logic; attribute dont_touch of G2023: signal is true;
	signal G2024: std_logic; attribute dont_touch of G2024: signal is true;
	signal G2025: std_logic; attribute dont_touch of G2025: signal is true;
	signal G2028: std_logic; attribute dont_touch of G2028: signal is true;
	signal G2031: std_logic; attribute dont_touch of G2031: signal is true;
	signal G2034: std_logic; attribute dont_touch of G2034: signal is true;
	signal G2037: std_logic; attribute dont_touch of G2037: signal is true;
	signal G2038: std_logic; attribute dont_touch of G2038: signal is true;
	signal G2039: std_logic; attribute dont_touch of G2039: signal is true;
	signal G2040: std_logic; attribute dont_touch of G2040: signal is true;
	signal G2041: std_logic; attribute dont_touch of G2041: signal is true;
	signal G2042: std_logic; attribute dont_touch of G2042: signal is true;
	signal G2043: std_logic; attribute dont_touch of G2043: signal is true;
	signal G2044: std_logic; attribute dont_touch of G2044: signal is true;
	signal G2045: std_logic; attribute dont_touch of G2045: signal is true;
	signal G2046: std_logic; attribute dont_touch of G2046: signal is true;
	signal G2047: std_logic; attribute dont_touch of G2047: signal is true;
	signal G2050: std_logic; attribute dont_touch of G2050: signal is true;
	signal G2054: std_logic; attribute dont_touch of G2054: signal is true;
	signal G2055: std_logic; attribute dont_touch of G2055: signal is true;
	signal G2056: std_logic; attribute dont_touch of G2056: signal is true;
	signal G2057: std_logic; attribute dont_touch of G2057: signal is true;
	signal G2060: std_logic; attribute dont_touch of G2060: signal is true;
	signal G2061: std_logic; attribute dont_touch of G2061: signal is true;
	signal G2067: std_logic; attribute dont_touch of G2067: signal is true;
	signal G2068: std_logic; attribute dont_touch of G2068: signal is true;
	signal G2069: std_logic; attribute dont_touch of G2069: signal is true;
	signal G2070: std_logic; attribute dont_touch of G2070: signal is true;
	signal G2071: std_logic; attribute dont_touch of G2071: signal is true;
	signal G2072: std_logic; attribute dont_touch of G2072: signal is true;
	signal G2073: std_logic; attribute dont_touch of G2073: signal is true;
	signal G2074: std_logic; attribute dont_touch of G2074: signal is true;
	signal G2075: std_logic; attribute dont_touch of G2075: signal is true;
	signal G2076: std_logic; attribute dont_touch of G2076: signal is true;
	signal G2077: std_logic; attribute dont_touch of G2077: signal is true;
	signal G2078: std_logic; attribute dont_touch of G2078: signal is true;
	signal G2079: std_logic; attribute dont_touch of G2079: signal is true;
	signal G2080: std_logic; attribute dont_touch of G2080: signal is true;
	signal G2081: std_logic; attribute dont_touch of G2081: signal is true;
	signal G2082: std_logic; attribute dont_touch of G2082: signal is true;
	signal G2083: std_logic; attribute dont_touch of G2083: signal is true;
	signal G2084: std_logic; attribute dont_touch of G2084: signal is true;
	signal G2085: std_logic; attribute dont_touch of G2085: signal is true;
	signal G2086: std_logic; attribute dont_touch of G2086: signal is true;
	signal G2087: std_logic; attribute dont_touch of G2087: signal is true;
	signal G2088: std_logic; attribute dont_touch of G2088: signal is true;
	signal G2089: std_logic; attribute dont_touch of G2089: signal is true;
	signal G2090: std_logic; attribute dont_touch of G2090: signal is true;
	signal G2091: std_logic; attribute dont_touch of G2091: signal is true;
	signal G2094: std_logic; attribute dont_touch of G2094: signal is true;
	signal G2095: std_logic; attribute dont_touch of G2095: signal is true;
	signal G2096: std_logic; attribute dont_touch of G2096: signal is true;
	signal G2097: std_logic; attribute dont_touch of G2097: signal is true;
	signal G2098: std_logic; attribute dont_touch of G2098: signal is true;
	signal G2099: std_logic; attribute dont_touch of G2099: signal is true;
	signal G2100: std_logic; attribute dont_touch of G2100: signal is true;
	signal G2101: std_logic; attribute dont_touch of G2101: signal is true;
	signal G2102: std_logic; attribute dont_touch of G2102: signal is true;
	signal G2103: std_logic; attribute dont_touch of G2103: signal is true;
	signal G2104: std_logic; attribute dont_touch of G2104: signal is true;
	signal G2105: std_logic; attribute dont_touch of G2105: signal is true;
	signal G2106: std_logic; attribute dont_touch of G2106: signal is true;
	signal G2107: std_logic; attribute dont_touch of G2107: signal is true;
	signal G2108: std_logic; attribute dont_touch of G2108: signal is true;
	signal G2109: std_logic; attribute dont_touch of G2109: signal is true;
	signal G2110: std_logic; attribute dont_touch of G2110: signal is true;
	signal G2111: std_logic; attribute dont_touch of G2111: signal is true;
	signal G2112: std_logic; attribute dont_touch of G2112: signal is true;
	signal G2115: std_logic; attribute dont_touch of G2115: signal is true;
	signal G2116: std_logic; attribute dont_touch of G2116: signal is true;
	signal G2117: std_logic; attribute dont_touch of G2117: signal is true;
	signal G2118: std_logic; attribute dont_touch of G2118: signal is true;
	signal G2119: std_logic; attribute dont_touch of G2119: signal is true;
	signal G2120: std_logic; attribute dont_touch of G2120: signal is true;
	signal G2121: std_logic; attribute dont_touch of G2121: signal is true;
	signal G2122: std_logic; attribute dont_touch of G2122: signal is true;
	signal G2123: std_logic; attribute dont_touch of G2123: signal is true;
	signal G2124: std_logic; attribute dont_touch of G2124: signal is true;
	signal G2125: std_logic; attribute dont_touch of G2125: signal is true;
	signal G2126: std_logic; attribute dont_touch of G2126: signal is true;
	signal G2130: std_logic; attribute dont_touch of G2130: signal is true;
	signal G2131: std_logic; attribute dont_touch of G2131: signal is true;
	signal G2132: std_logic; attribute dont_touch of G2132: signal is true;
	signal G2135: std_logic; attribute dont_touch of G2135: signal is true;
	signal G2154: std_logic; attribute dont_touch of G2154: signal is true;
	signal G2155: std_logic; attribute dont_touch of G2155: signal is true;
	signal G2156: std_logic; attribute dont_touch of G2156: signal is true;
	signal G2157: std_logic; attribute dont_touch of G2157: signal is true;
	signal G2158: std_logic; attribute dont_touch of G2158: signal is true;
	signal G2159: std_logic; attribute dont_touch of G2159: signal is true;
	signal G2160: std_logic; attribute dont_touch of G2160: signal is true;
	signal G2161: std_logic; attribute dont_touch of G2161: signal is true;
	signal G2162: std_logic; attribute dont_touch of G2162: signal is true;
	signal G2163: std_logic; attribute dont_touch of G2163: signal is true;
	signal G2164: std_logic; attribute dont_touch of G2164: signal is true;
	signal G2165: std_logic; attribute dont_touch of G2165: signal is true;
	signal G2166: std_logic; attribute dont_touch of G2166: signal is true;
	signal G2167: std_logic; attribute dont_touch of G2167: signal is true;
	signal G2168: std_logic; attribute dont_touch of G2168: signal is true;
	signal G2169: std_logic; attribute dont_touch of G2169: signal is true;
	signal G2170: std_logic; attribute dont_touch of G2170: signal is true;
	signal G2171: std_logic; attribute dont_touch of G2171: signal is true;
	signal G2172: std_logic; attribute dont_touch of G2172: signal is true;
	signal G2173: std_logic; attribute dont_touch of G2173: signal is true;
	signal G2174: std_logic; attribute dont_touch of G2174: signal is true;
	signal G2175: std_logic; attribute dont_touch of G2175: signal is true;
	signal G2176: std_logic; attribute dont_touch of G2176: signal is true;
	signal G2177: std_logic; attribute dont_touch of G2177: signal is true;
	signal G2178: std_logic; attribute dont_touch of G2178: signal is true;
	signal G2179: std_logic; attribute dont_touch of G2179: signal is true;
	signal G2180: std_logic; attribute dont_touch of G2180: signal is true;
	signal G2181: std_logic; attribute dont_touch of G2181: signal is true;
	signal G2184: std_logic; attribute dont_touch of G2184: signal is true;
	signal G2185: std_logic; attribute dont_touch of G2185: signal is true;
	signal G2186: std_logic; attribute dont_touch of G2186: signal is true;
	signal G2187: std_logic; attribute dont_touch of G2187: signal is true;
	signal G2190: std_logic; attribute dont_touch of G2190: signal is true;
	signal G2191: std_logic; attribute dont_touch of G2191: signal is true;
	signal G2194: std_logic; attribute dont_touch of G2194: signal is true;
	signal G2195: std_logic; attribute dont_touch of G2195: signal is true;
	signal G2196: std_logic; attribute dont_touch of G2196: signal is true;
	signal G2197: std_logic; attribute dont_touch of G2197: signal is true;
	signal G2198: std_logic; attribute dont_touch of G2198: signal is true;
	signal G2199: std_logic; attribute dont_touch of G2199: signal is true;
	signal G2200: std_logic; attribute dont_touch of G2200: signal is true;
	signal G2201: std_logic; attribute dont_touch of G2201: signal is true;
	signal G2202: std_logic; attribute dont_touch of G2202: signal is true;
	signal G2203: std_logic; attribute dont_touch of G2203: signal is true;
	signal G2204: std_logic; attribute dont_touch of G2204: signal is true;
	signal G2205: std_logic; attribute dont_touch of G2205: signal is true;
	signal G2206: std_logic; attribute dont_touch of G2206: signal is true;
	signal G2207: std_logic; attribute dont_touch of G2207: signal is true;
	signal G2208: std_logic; attribute dont_touch of G2208: signal is true;
	signal G2209: std_logic; attribute dont_touch of G2209: signal is true;
	signal G2210: std_logic; attribute dont_touch of G2210: signal is true;
	signal G2211: std_logic; attribute dont_touch of G2211: signal is true;
	signal G2212: std_logic; attribute dont_touch of G2212: signal is true;
	signal G2213: std_logic; attribute dont_touch of G2213: signal is true;
	signal G2214: std_logic; attribute dont_touch of G2214: signal is true;
	signal G2215: std_logic; attribute dont_touch of G2215: signal is true;
	signal G2216: std_logic; attribute dont_touch of G2216: signal is true;
	signal G2217: std_logic; attribute dont_touch of G2217: signal is true;
	signal G2218: std_logic; attribute dont_touch of G2218: signal is true;
	signal G2219: std_logic; attribute dont_touch of G2219: signal is true;
	signal G2220: std_logic; attribute dont_touch of G2220: signal is true;
	signal G2221: std_logic; attribute dont_touch of G2221: signal is true;
	signal G2222: std_logic; attribute dont_touch of G2222: signal is true;
	signal G2223: std_logic; attribute dont_touch of G2223: signal is true;
	signal G2224: std_logic; attribute dont_touch of G2224: signal is true;
	signal G2225: std_logic; attribute dont_touch of G2225: signal is true;
	signal G2226: std_logic; attribute dont_touch of G2226: signal is true;
	signal G2227: std_logic; attribute dont_touch of G2227: signal is true;
	signal G2228: std_logic; attribute dont_touch of G2228: signal is true;
	signal G2229: std_logic; attribute dont_touch of G2229: signal is true;
	signal G2230: std_logic; attribute dont_touch of G2230: signal is true;
	signal G2231: std_logic; attribute dont_touch of G2231: signal is true;
	signal G2232: std_logic; attribute dont_touch of G2232: signal is true;
	signal G2233: std_logic; attribute dont_touch of G2233: signal is true;
	signal G2234: std_logic; attribute dont_touch of G2234: signal is true;
	signal G2235: std_logic; attribute dont_touch of G2235: signal is true;
	signal G2236: std_logic; attribute dont_touch of G2236: signal is true;
	signal G2237: std_logic; attribute dont_touch of G2237: signal is true;
	signal G2238: std_logic; attribute dont_touch of G2238: signal is true;
	signal G2239: std_logic; attribute dont_touch of G2239: signal is true;
	signal G2240: std_logic; attribute dont_touch of G2240: signal is true;
	signal G2241: std_logic; attribute dont_touch of G2241: signal is true;
	signal G2242: std_logic; attribute dont_touch of G2242: signal is true;
	signal G2243: std_logic; attribute dont_touch of G2243: signal is true;
	signal G2244: std_logic; attribute dont_touch of G2244: signal is true;
	signal G2245: std_logic; attribute dont_touch of G2245: signal is true;
	signal G2246: std_logic; attribute dont_touch of G2246: signal is true;
	signal G2247: std_logic; attribute dont_touch of G2247: signal is true;
	signal G2248: std_logic; attribute dont_touch of G2248: signal is true;
	signal G2249: std_logic; attribute dont_touch of G2249: signal is true;
	signal G2250: std_logic; attribute dont_touch of G2250: signal is true;
	signal G2251: std_logic; attribute dont_touch of G2251: signal is true;
	signal G2252: std_logic; attribute dont_touch of G2252: signal is true;
	signal G2253: std_logic; attribute dont_touch of G2253: signal is true;
	signal G2254: std_logic; attribute dont_touch of G2254: signal is true;
	signal G2255: std_logic; attribute dont_touch of G2255: signal is true;
	signal G2256: std_logic; attribute dont_touch of G2256: signal is true;
	signal G2257: std_logic; attribute dont_touch of G2257: signal is true;
	signal G2258: std_logic; attribute dont_touch of G2258: signal is true;
	signal G2259: std_logic; attribute dont_touch of G2259: signal is true;
	signal G2260: std_logic; attribute dont_touch of G2260: signal is true;
	signal G2261: std_logic; attribute dont_touch of G2261: signal is true;
	signal G2264: std_logic; attribute dont_touch of G2264: signal is true;
	signal G2267: std_logic; attribute dont_touch of G2267: signal is true;
	signal G2268: std_logic; attribute dont_touch of G2268: signal is true;
	signal G2269: std_logic; attribute dont_touch of G2269: signal is true;
	signal G2270: std_logic; attribute dont_touch of G2270: signal is true;
	signal G2271: std_logic; attribute dont_touch of G2271: signal is true;
	signal G2272: std_logic; attribute dont_touch of G2272: signal is true;
	signal G2273: std_logic; attribute dont_touch of G2273: signal is true;
	signal G2274: std_logic; attribute dont_touch of G2274: signal is true;
	signal G2275: std_logic; attribute dont_touch of G2275: signal is true;
	signal G2276: std_logic; attribute dont_touch of G2276: signal is true;
	signal G2296: std_logic; attribute dont_touch of G2296: signal is true;
	signal G2297: std_logic; attribute dont_touch of G2297: signal is true;
	signal G2298: std_logic; attribute dont_touch of G2298: signal is true;
	signal G2299: std_logic; attribute dont_touch of G2299: signal is true;
	signal G2302: std_logic; attribute dont_touch of G2302: signal is true;
	signal G2303: std_logic; attribute dont_touch of G2303: signal is true;
	signal G2304: std_logic; attribute dont_touch of G2304: signal is true;
	signal G2305: std_logic; attribute dont_touch of G2305: signal is true;
	signal G2306: std_logic; attribute dont_touch of G2306: signal is true;
	signal G2309: std_logic; attribute dont_touch of G2309: signal is true;
	signal G2310: std_logic; attribute dont_touch of G2310: signal is true;
	signal G2315: std_logic; attribute dont_touch of G2315: signal is true;
	signal G2316: std_logic; attribute dont_touch of G2316: signal is true;
	signal G2317: std_logic; attribute dont_touch of G2317: signal is true;
	signal G2320: std_logic; attribute dont_touch of G2320: signal is true;
	signal G2321: std_logic; attribute dont_touch of G2321: signal is true;
	signal G2322: std_logic; attribute dont_touch of G2322: signal is true;
	signal G2325: std_logic; attribute dont_touch of G2325: signal is true;
	signal G2328: std_logic; attribute dont_touch of G2328: signal is true;
	signal G2329: std_logic; attribute dont_touch of G2329: signal is true;
	signal G2330: std_logic; attribute dont_touch of G2330: signal is true;
	signal G2331: std_logic; attribute dont_touch of G2331: signal is true;
	signal G2334: std_logic; attribute dont_touch of G2334: signal is true;
	signal G2335: std_logic; attribute dont_touch of G2335: signal is true;
	signal G2336: std_logic; attribute dont_touch of G2336: signal is true;
	signal G2337: std_logic; attribute dont_touch of G2337: signal is true;
	signal G2338: std_logic; attribute dont_touch of G2338: signal is true;
	signal G2339: std_logic; attribute dont_touch of G2339: signal is true;
	signal G2340: std_logic; attribute dont_touch of G2340: signal is true;
	signal G2341: std_logic; attribute dont_touch of G2341: signal is true;
	signal G2342: std_logic; attribute dont_touch of G2342: signal is true;
	signal G2343: std_logic; attribute dont_touch of G2343: signal is true;
	signal G2344: std_logic; attribute dont_touch of G2344: signal is true;
	signal G2345: std_logic; attribute dont_touch of G2345: signal is true;
	signal G2346: std_logic; attribute dont_touch of G2346: signal is true;
	signal G2347: std_logic; attribute dont_touch of G2347: signal is true;
	signal G2348: std_logic; attribute dont_touch of G2348: signal is true;
	signal G2349: std_logic; attribute dont_touch of G2349: signal is true;
	signal G2350: std_logic; attribute dont_touch of G2350: signal is true;
	signal G2351: std_logic; attribute dont_touch of G2351: signal is true;
	signal G2352: std_logic; attribute dont_touch of G2352: signal is true;
	signal G2353: std_logic; attribute dont_touch of G2353: signal is true;
	signal G2354: std_logic; attribute dont_touch of G2354: signal is true;
	signal G2356: std_logic; attribute dont_touch of G2356: signal is true;
	signal G2363: std_logic; attribute dont_touch of G2363: signal is true;
	signal G2364: std_logic; attribute dont_touch of G2364: signal is true;
	signal G2368: std_logic; attribute dont_touch of G2368: signal is true;
	signal G2369: std_logic; attribute dont_touch of G2369: signal is true;
	signal G2372: std_logic; attribute dont_touch of G2372: signal is true;
	signal G2373: std_logic; attribute dont_touch of G2373: signal is true;
	signal G2374: std_logic; attribute dont_touch of G2374: signal is true;
	signal G2379: std_logic; attribute dont_touch of G2379: signal is true;
	signal G2380: std_logic; attribute dont_touch of G2380: signal is true;
	signal G2381: std_logic; attribute dont_touch of G2381: signal is true;
	signal G2382: std_logic; attribute dont_touch of G2382: signal is true;
	signal G2389: std_logic; attribute dont_touch of G2389: signal is true;
	signal G2390: std_logic; attribute dont_touch of G2390: signal is true;
	signal G2391: std_logic; attribute dont_touch of G2391: signal is true;
	signal G2395: std_logic; attribute dont_touch of G2395: signal is true;
	signal G2396: std_logic; attribute dont_touch of G2396: signal is true;
	signal G2399: std_logic; attribute dont_touch of G2399: signal is true;
	signal G2405: std_logic; attribute dont_touch of G2405: signal is true;
	signal G2406: std_logic; attribute dont_touch of G2406: signal is true;
	signal G2407: std_logic; attribute dont_touch of G2407: signal is true;
	signal G2410: std_logic; attribute dont_touch of G2410: signal is true;
	signal G2411: std_logic; attribute dont_touch of G2411: signal is true;
	signal G2418: std_logic; attribute dont_touch of G2418: signal is true;
	signal G2419: std_logic; attribute dont_touch of G2419: signal is true;
	signal G2420: std_logic; attribute dont_touch of G2420: signal is true;
	signal G2421: std_logic; attribute dont_touch of G2421: signal is true;
	signal G2424: std_logic; attribute dont_touch of G2424: signal is true;
	signal G2431: std_logic; attribute dont_touch of G2431: signal is true;
	signal G2432: std_logic; attribute dont_touch of G2432: signal is true;
	signal G2433: std_logic; attribute dont_touch of G2433: signal is true;
	signal G2434: std_logic; attribute dont_touch of G2434: signal is true;
	signal G2435: std_logic; attribute dont_touch of G2435: signal is true;
	signal G2436: std_logic; attribute dont_touch of G2436: signal is true;
	signal G2437: std_logic; attribute dont_touch of G2437: signal is true;
	signal G2438: std_logic; attribute dont_touch of G2438: signal is true;
	signal G2439: std_logic; attribute dont_touch of G2439: signal is true;
	signal G2444: std_logic; attribute dont_touch of G2444: signal is true;
	signal G2445: std_logic; attribute dont_touch of G2445: signal is true;
	signal G2446: std_logic; attribute dont_touch of G2446: signal is true;
	signal G2449: std_logic; attribute dont_touch of G2449: signal is true;
	signal G2450: std_logic; attribute dont_touch of G2450: signal is true;
	signal G2451: std_logic; attribute dont_touch of G2451: signal is true;
	signal G2454: std_logic; attribute dont_touch of G2454: signal is true;
	signal G2455: std_logic; attribute dont_touch of G2455: signal is true;
	signal G2456: std_logic; attribute dont_touch of G2456: signal is true;
	signal G2459: std_logic; attribute dont_touch of G2459: signal is true;
	signal G2462: std_logic; attribute dont_touch of G2462: signal is true;
	signal G2475: std_logic; attribute dont_touch of G2475: signal is true;
	signal G2478: std_logic; attribute dont_touch of G2478: signal is true;
	signal G2479: std_logic; attribute dont_touch of G2479: signal is true;
	signal G2480: std_logic; attribute dont_touch of G2480: signal is true;
	signal G2481: std_logic; attribute dont_touch of G2481: signal is true;
	signal G2482: std_logic; attribute dont_touch of G2482: signal is true;
	signal G2493: std_logic; attribute dont_touch of G2493: signal is true;
	signal G2496: std_logic; attribute dont_touch of G2496: signal is true;
	signal G2499: std_logic; attribute dont_touch of G2499: signal is true;
	signal G2500: std_logic; attribute dont_touch of G2500: signal is true;
	signal G2501: std_logic; attribute dont_touch of G2501: signal is true;
	signal G2502: std_logic; attribute dont_touch of G2502: signal is true;
	signal G2503: std_logic; attribute dont_touch of G2503: signal is true;
	signal G2506: std_logic; attribute dont_touch of G2506: signal is true;
	signal G2507: std_logic; attribute dont_touch of G2507: signal is true;
	signal G2508: std_logic; attribute dont_touch of G2508: signal is true;
	signal G2509: std_logic; attribute dont_touch of G2509: signal is true;
	signal G2510: std_logic; attribute dont_touch of G2510: signal is true;
	signal G2511: std_logic; attribute dont_touch of G2511: signal is true;
	signal G2514: std_logic; attribute dont_touch of G2514: signal is true;
	signal G2515: std_logic; attribute dont_touch of G2515: signal is true;
	signal G2516: std_logic; attribute dont_touch of G2516: signal is true;
	signal G2517: std_logic; attribute dont_touch of G2517: signal is true;
	signal G2518: std_logic; attribute dont_touch of G2518: signal is true;
	signal G2521: std_logic; attribute dont_touch of G2521: signal is true;
	signal G2522: std_logic; attribute dont_touch of G2522: signal is true;
	signal G2523: std_logic; attribute dont_touch of G2523: signal is true;
	signal G2524: std_logic; attribute dont_touch of G2524: signal is true;
	signal G2525: std_logic; attribute dont_touch of G2525: signal is true;
	signal G2528: std_logic; attribute dont_touch of G2528: signal is true;
	signal G2529: std_logic; attribute dont_touch of G2529: signal is true;
	signal G2530: std_logic; attribute dont_touch of G2530: signal is true;
	signal G2531: std_logic; attribute dont_touch of G2531: signal is true;
	signal G2534: std_logic; attribute dont_touch of G2534: signal is true;
	signal G2537: std_logic; attribute dont_touch of G2537: signal is true;
	signal G2538: std_logic; attribute dont_touch of G2538: signal is true;
	signal G2539: std_logic; attribute dont_touch of G2539: signal is true;
	signal G2540: std_logic; attribute dont_touch of G2540: signal is true;
	signal G2541: std_logic; attribute dont_touch of G2541: signal is true;
	signal G2542: std_logic; attribute dont_touch of G2542: signal is true;
	signal G2543: std_logic; attribute dont_touch of G2543: signal is true;
	signal G2544: std_logic; attribute dont_touch of G2544: signal is true;
	signal G2547: std_logic; attribute dont_touch of G2547: signal is true;
	signal G2548: std_logic; attribute dont_touch of G2548: signal is true;
	signal G2549: std_logic; attribute dont_touch of G2549: signal is true;
	signal G2550: std_logic; attribute dont_touch of G2550: signal is true;
	signal G2554: std_logic; attribute dont_touch of G2554: signal is true;
	signal G2555: std_logic; attribute dont_touch of G2555: signal is true;
	signal G2556: std_logic; attribute dont_touch of G2556: signal is true;
	signal G2557: std_logic; attribute dont_touch of G2557: signal is true;
	signal G2560: std_logic; attribute dont_touch of G2560: signal is true;
	signal G2561: std_logic; attribute dont_touch of G2561: signal is true;
	signal G2562: std_logic; attribute dont_touch of G2562: signal is true;
	signal G2563: std_logic; attribute dont_touch of G2563: signal is true;
	signal G2564: std_logic; attribute dont_touch of G2564: signal is true;
	signal G2569: std_logic; attribute dont_touch of G2569: signal is true;
	signal G2570: std_logic; attribute dont_touch of G2570: signal is true;
	signal G2571: std_logic; attribute dont_touch of G2571: signal is true;
	signal G2578: std_logic; attribute dont_touch of G2578: signal is true;
	signal G2579: std_logic; attribute dont_touch of G2579: signal is true;
	signal G2586: std_logic; attribute dont_touch of G2586: signal is true;
	signal G2593: std_logic; attribute dont_touch of G2593: signal is true;
	signal G2613: std_logic; attribute dont_touch of G2613: signal is true;
	signal G2614: std_logic; attribute dont_touch of G2614: signal is true;
	signal G2617: std_logic; attribute dont_touch of G2617: signal is true;
	signal G2620: std_logic; attribute dont_touch of G2620: signal is true;
	signal G2623: std_logic; attribute dont_touch of G2623: signal is true;
	signal G2626: std_logic; attribute dont_touch of G2626: signal is true;
	signal G2629: std_logic; attribute dont_touch of G2629: signal is true;
	signal G2632: std_logic; attribute dont_touch of G2632: signal is true;
	signal G2635: std_logic; attribute dont_touch of G2635: signal is true;
	signal G2638: std_logic; attribute dont_touch of G2638: signal is true;
	signal G2639: std_logic; attribute dont_touch of G2639: signal is true;
	signal G2640: std_logic; attribute dont_touch of G2640: signal is true;
	signal G2641: std_logic; attribute dont_touch of G2641: signal is true;
	signal G2642: std_logic; attribute dont_touch of G2642: signal is true;
	signal G2643: std_logic; attribute dont_touch of G2643: signal is true;
	signal G2644: std_logic; attribute dont_touch of G2644: signal is true;
	signal G2645: std_logic; attribute dont_touch of G2645: signal is true;
	signal G2646: std_logic; attribute dont_touch of G2646: signal is true;
	signal G2647: std_logic; attribute dont_touch of G2647: signal is true;
	signal G2649: std_logic; attribute dont_touch of G2649: signal is true;
	signal G2650: std_logic; attribute dont_touch of G2650: signal is true;
	signal G2651: std_logic; attribute dont_touch of G2651: signal is true;
	signal G2652: std_logic; attribute dont_touch of G2652: signal is true;
	signal G2653: std_logic; attribute dont_touch of G2653: signal is true;
	signal G2654: std_logic; attribute dont_touch of G2654: signal is true;
	signal G2655: std_logic; attribute dont_touch of G2655: signal is true;
	signal G2662: std_logic; attribute dont_touch of G2662: signal is true;
	signal G2669: std_logic; attribute dont_touch of G2669: signal is true;
	signal G2677: std_logic; attribute dont_touch of G2677: signal is true;
	signal G2683: std_logic; attribute dont_touch of G2683: signal is true;
	signal G2689: std_logic; attribute dont_touch of G2689: signal is true;
	signal G2695: std_logic; attribute dont_touch of G2695: signal is true;
	signal G2701: std_logic; attribute dont_touch of G2701: signal is true;
	signal G2707: std_logic; attribute dont_touch of G2707: signal is true;
	signal G2713: std_logic; attribute dont_touch of G2713: signal is true;
	signal G2719: std_logic; attribute dont_touch of G2719: signal is true;
	signal G2725: std_logic; attribute dont_touch of G2725: signal is true;
	signal G2726: std_logic; attribute dont_touch of G2726: signal is true;
	signal G2727: std_logic; attribute dont_touch of G2727: signal is true;
	signal G2728: std_logic; attribute dont_touch of G2728: signal is true;
	signal G2731: std_logic; attribute dont_touch of G2731: signal is true;
	signal G2732: std_logic; attribute dont_touch of G2732: signal is true;
	signal G2733: std_logic; attribute dont_touch of G2733: signal is true;
	signal G2742: std_logic; attribute dont_touch of G2742: signal is true;
	signal G2743: std_logic; attribute dont_touch of G2743: signal is true;
	signal G2744: std_logic; attribute dont_touch of G2744: signal is true;
	signal G2745: std_logic; attribute dont_touch of G2745: signal is true;
	signal G2748: std_logic; attribute dont_touch of G2748: signal is true;
	signal G2749: std_logic; attribute dont_touch of G2749: signal is true;
	signal G2750: std_logic; attribute dont_touch of G2750: signal is true;
	signal G2751: std_logic; attribute dont_touch of G2751: signal is true;
	signal G2752: std_logic; attribute dont_touch of G2752: signal is true;
	signal G2753: std_logic; attribute dont_touch of G2753: signal is true;
	signal G2754: std_logic; attribute dont_touch of G2754: signal is true;
	signal G2755: std_logic; attribute dont_touch of G2755: signal is true;
	signal G2756: std_logic; attribute dont_touch of G2756: signal is true;
	signal G2757: std_logic; attribute dont_touch of G2757: signal is true;
	signal G2758: std_logic; attribute dont_touch of G2758: signal is true;
	signal G2759: std_logic; attribute dont_touch of G2759: signal is true;
	signal G2760: std_logic; attribute dont_touch of G2760: signal is true;
	signal G2763: std_logic; attribute dont_touch of G2763: signal is true;
	signal G2764: std_logic; attribute dont_touch of G2764: signal is true;
	signal G2765: std_logic; attribute dont_touch of G2765: signal is true;
	signal G2771: std_logic; attribute dont_touch of G2771: signal is true;
	signal G2772: std_logic; attribute dont_touch of G2772: signal is true;
	signal G2773: std_logic; attribute dont_touch of G2773: signal is true;
	signal G2774: std_logic; attribute dont_touch of G2774: signal is true;
	signal G2775: std_logic; attribute dont_touch of G2775: signal is true;
	signal G2776: std_logic; attribute dont_touch of G2776: signal is true;
	signal G2777: std_logic; attribute dont_touch of G2777: signal is true;
	signal G2778: std_logic; attribute dont_touch of G2778: signal is true;
	signal G2779: std_logic; attribute dont_touch of G2779: signal is true;
	signal G2789: std_logic; attribute dont_touch of G2789: signal is true;
	signal G2790: std_logic; attribute dont_touch of G2790: signal is true;
	signal G2791: std_logic; attribute dont_touch of G2791: signal is true;
	signal G2792: std_logic; attribute dont_touch of G2792: signal is true;
	signal G2793: std_logic; attribute dont_touch of G2793: signal is true;
	signal G2794: std_logic; attribute dont_touch of G2794: signal is true;
	signal G2795: std_logic; attribute dont_touch of G2795: signal is true;
	signal G2796: std_logic; attribute dont_touch of G2796: signal is true;
	signal G2797: std_logic; attribute dont_touch of G2797: signal is true;
	signal G2798: std_logic; attribute dont_touch of G2798: signal is true;
	signal G2799: std_logic; attribute dont_touch of G2799: signal is true;
	signal G2800: std_logic; attribute dont_touch of G2800: signal is true;
	signal G2801: std_logic; attribute dont_touch of G2801: signal is true;
	signal G2802: std_logic; attribute dont_touch of G2802: signal is true;
	signal G2803: std_logic; attribute dont_touch of G2803: signal is true;
	signal G2804: std_logic; attribute dont_touch of G2804: signal is true;
	signal G2807: std_logic; attribute dont_touch of G2807: signal is true;
	signal G2808: std_logic; attribute dont_touch of G2808: signal is true;
	signal G2809: std_logic; attribute dont_touch of G2809: signal is true;
	signal G2812: std_logic; attribute dont_touch of G2812: signal is true;
	signal G2813: std_logic; attribute dont_touch of G2813: signal is true;
	signal G2814: std_logic; attribute dont_touch of G2814: signal is true;
	signal G2817: std_logic; attribute dont_touch of G2817: signal is true;
	signal G2818: std_logic; attribute dont_touch of G2818: signal is true;
	signal G2819: std_logic; attribute dont_touch of G2819: signal is true;
	signal G2820: std_logic; attribute dont_touch of G2820: signal is true;
	signal G2821: std_logic; attribute dont_touch of G2821: signal is true;
	signal G2824: std_logic; attribute dont_touch of G2824: signal is true;
	signal G2825: std_logic; attribute dont_touch of G2825: signal is true;
	signal G2826: std_logic; attribute dont_touch of G2826: signal is true;
	signal G2827: std_logic; attribute dont_touch of G2827: signal is true;
	signal G2828: std_logic; attribute dont_touch of G2828: signal is true;
	signal G2829: std_logic; attribute dont_touch of G2829: signal is true;
	signal G2832: std_logic; attribute dont_touch of G2832: signal is true;
	signal G2833: std_logic; attribute dont_touch of G2833: signal is true;
	signal G2834: std_logic; attribute dont_touch of G2834: signal is true;
	signal G2837: std_logic; attribute dont_touch of G2837: signal is true;
	signal G2838: std_logic; attribute dont_touch of G2838: signal is true;
	signal G2839: std_logic; attribute dont_touch of G2839: signal is true;
	signal G2840: std_logic; attribute dont_touch of G2840: signal is true;
	signal G2843: std_logic; attribute dont_touch of G2843: signal is true;
	signal G2844: std_logic; attribute dont_touch of G2844: signal is true;
	signal G2845: std_logic; attribute dont_touch of G2845: signal is true;
	signal G2846: std_logic; attribute dont_touch of G2846: signal is true;
	signal G2847: std_logic; attribute dont_touch of G2847: signal is true;
	signal G2850: std_logic; attribute dont_touch of G2850: signal is true;
	signal G2851: std_logic; attribute dont_touch of G2851: signal is true;
	signal G2852: std_logic; attribute dont_touch of G2852: signal is true;
	signal G2853: std_logic; attribute dont_touch of G2853: signal is true;
	signal G2854: std_logic; attribute dont_touch of G2854: signal is true;
	signal G2855: std_logic; attribute dont_touch of G2855: signal is true;
	signal G2858: std_logic; attribute dont_touch of G2858: signal is true;
	signal G2859: std_logic; attribute dont_touch of G2859: signal is true;
	signal G2860: std_logic; attribute dont_touch of G2860: signal is true;
	signal G2861: std_logic; attribute dont_touch of G2861: signal is true;
	signal G2862: std_logic; attribute dont_touch of G2862: signal is true;
	signal G2863: std_logic; attribute dont_touch of G2863: signal is true;
	signal G2864: std_logic; attribute dont_touch of G2864: signal is true;
	signal G2867: std_logic; attribute dont_touch of G2867: signal is true;
	signal G2868: std_logic; attribute dont_touch of G2868: signal is true;
	signal G2871: std_logic; attribute dont_touch of G2871: signal is true;
	signal G2872: std_logic; attribute dont_touch of G2872: signal is true;
	signal G2873: std_logic; attribute dont_touch of G2873: signal is true;
	signal G2874: std_logic; attribute dont_touch of G2874: signal is true;
	signal G2877: std_logic; attribute dont_touch of G2877: signal is true;
	signal G2880: std_logic; attribute dont_touch of G2880: signal is true;
	signal G2881: std_logic; attribute dont_touch of G2881: signal is true;
	signal G2882: std_logic; attribute dont_touch of G2882: signal is true;
	signal G2883: std_logic; attribute dont_touch of G2883: signal is true;
	signal G2884: std_logic; attribute dont_touch of G2884: signal is true;
	signal G2885: std_logic; attribute dont_touch of G2885: signal is true;
	signal G2888: std_logic; attribute dont_touch of G2888: signal is true;
	signal G2889: std_logic; attribute dont_touch of G2889: signal is true;
	signal G2890: std_logic; attribute dont_touch of G2890: signal is true;
	signal G2891: std_logic; attribute dont_touch of G2891: signal is true;
	signal G2892: std_logic; attribute dont_touch of G2892: signal is true;
	signal G2895: std_logic; attribute dont_touch of G2895: signal is true;
	signal G2896: std_logic; attribute dont_touch of G2896: signal is true;
	signal G2902: std_logic; attribute dont_touch of G2902: signal is true;
	signal G2903: std_logic; attribute dont_touch of G2903: signal is true;
	signal G2904: std_logic; attribute dont_touch of G2904: signal is true;
	signal G2905: std_logic; attribute dont_touch of G2905: signal is true;
	signal G2906: std_logic; attribute dont_touch of G2906: signal is true;
	signal G2907: std_logic; attribute dont_touch of G2907: signal is true;
	signal G2908: std_logic; attribute dont_touch of G2908: signal is true;
	signal G2909: std_logic; attribute dont_touch of G2909: signal is true;
	signal G2910: std_logic; attribute dont_touch of G2910: signal is true;
	signal G2911: std_logic; attribute dont_touch of G2911: signal is true;
	signal G2912: std_logic; attribute dont_touch of G2912: signal is true;
	signal G2913: std_logic; attribute dont_touch of G2913: signal is true;
	signal G2914: std_logic; attribute dont_touch of G2914: signal is true;
	signal G2915: std_logic; attribute dont_touch of G2915: signal is true;
	signal G2916: std_logic; attribute dont_touch of G2916: signal is true;
	signal G2917: std_logic; attribute dont_touch of G2917: signal is true;
	signal G2918: std_logic; attribute dont_touch of G2918: signal is true;
	signal G2919: std_logic; attribute dont_touch of G2919: signal is true;
	signal G2920: std_logic; attribute dont_touch of G2920: signal is true;
	signal G2937: std_logic; attribute dont_touch of G2937: signal is true;
	signal G2938: std_logic; attribute dont_touch of G2938: signal is true;
	signal G2939: std_logic; attribute dont_touch of G2939: signal is true;
	signal G2940: std_logic; attribute dont_touch of G2940: signal is true;
	signal G2941: std_logic; attribute dont_touch of G2941: signal is true;
	signal G2942: std_logic; attribute dont_touch of G2942: signal is true;
	signal G2943: std_logic; attribute dont_touch of G2943: signal is true;
	signal G2944: std_logic; attribute dont_touch of G2944: signal is true;
	signal G2945: std_logic; attribute dont_touch of G2945: signal is true;
	signal G2946: std_logic; attribute dont_touch of G2946: signal is true;
	signal G2947: std_logic; attribute dont_touch of G2947: signal is true;
	signal G2948: std_logic; attribute dont_touch of G2948: signal is true;
	signal G2949: std_logic; attribute dont_touch of G2949: signal is true;
	signal G2950: std_logic; attribute dont_touch of G2950: signal is true;
	signal G2951: std_logic; attribute dont_touch of G2951: signal is true;
	signal G2952: std_logic; attribute dont_touch of G2952: signal is true;
	signal G2955: std_logic; attribute dont_touch of G2955: signal is true;
	signal G2956: std_logic; attribute dont_touch of G2956: signal is true;
	signal G2957: std_logic; attribute dont_touch of G2957: signal is true;
	signal G2958: std_logic; attribute dont_touch of G2958: signal is true;
	signal G2959: std_logic; attribute dont_touch of G2959: signal is true;
	signal G2960: std_logic; attribute dont_touch of G2960: signal is true;
	signal G2961: std_logic; attribute dont_touch of G2961: signal is true;
	signal G2962: std_logic; attribute dont_touch of G2962: signal is true;
	signal G2963: std_logic; attribute dont_touch of G2963: signal is true;
	signal G2964: std_logic; attribute dont_touch of G2964: signal is true;
	signal G2965: std_logic; attribute dont_touch of G2965: signal is true;
	signal G2970: std_logic; attribute dont_touch of G2970: signal is true;
	signal G2971: std_logic; attribute dont_touch of G2971: signal is true;
	signal G2979: std_logic; attribute dont_touch of G2979: signal is true;
	signal G2980: std_logic; attribute dont_touch of G2980: signal is true;
	signal G2981: std_logic; attribute dont_touch of G2981: signal is true;
	signal G2984: std_logic; attribute dont_touch of G2984: signal is true;
	signal G2985: std_logic; attribute dont_touch of G2985: signal is true;
	signal G2987: std_logic; attribute dont_touch of G2987: signal is true;
	signal G2988: std_logic; attribute dont_touch of G2988: signal is true;
	signal G2989: std_logic; attribute dont_touch of G2989: signal is true;
	signal G2990: std_logic; attribute dont_touch of G2990: signal is true;
	signal G2991: std_logic; attribute dont_touch of G2991: signal is true;
	signal G2994: std_logic; attribute dont_touch of G2994: signal is true;
	signal G2997: std_logic; attribute dont_touch of G2997: signal is true;
	signal G2998: std_logic; attribute dont_touch of G2998: signal is true;
	signal G3003: std_logic; attribute dont_touch of G3003: signal is true;
	signal G3008: std_logic; attribute dont_touch of G3008: signal is true;
	signal G3009: std_logic; attribute dont_touch of G3009: signal is true;
	signal G3010: std_logic; attribute dont_touch of G3010: signal is true;
	signal G3011: std_logic; attribute dont_touch of G3011: signal is true;
	signal G3012: std_logic; attribute dont_touch of G3012: signal is true;
	signal G3015: std_logic; attribute dont_touch of G3015: signal is true;
	signal G3037: std_logic; attribute dont_touch of G3037: signal is true;
	signal G3038: std_logic; attribute dont_touch of G3038: signal is true;
	signal G3039: std_logic; attribute dont_touch of G3039: signal is true;
	signal G3040: std_logic; attribute dont_touch of G3040: signal is true;
	signal G3041: std_logic; attribute dont_touch of G3041: signal is true;
	signal G3044: std_logic; attribute dont_touch of G3044: signal is true;
	signal G3047: std_logic; attribute dont_touch of G3047: signal is true;
	signal G3050: std_logic; attribute dont_touch of G3050: signal is true;
	signal G3051: std_logic; attribute dont_touch of G3051: signal is true;
	signal G3052: std_logic; attribute dont_touch of G3052: signal is true;
	signal G3055: std_logic; attribute dont_touch of G3055: signal is true;
	signal G3056: std_logic; attribute dont_touch of G3056: signal is true;
	signal G3060: std_logic; attribute dont_touch of G3060: signal is true;
	signal G3061: std_logic; attribute dont_touch of G3061: signal is true;
	signal G3062: std_logic; attribute dont_touch of G3062: signal is true;
	signal G3066: std_logic; attribute dont_touch of G3066: signal is true;
	signal G3067: std_logic; attribute dont_touch of G3067: signal is true;
	signal G3068: std_logic; attribute dont_touch of G3068: signal is true;
	signal G3070: std_logic; attribute dont_touch of G3070: signal is true;
	signal G3071: std_logic; attribute dont_touch of G3071: signal is true;
	signal G3076: std_logic; attribute dont_touch of G3076: signal is true;
	signal G3077: std_logic; attribute dont_touch of G3077: signal is true;
	signal G3086: std_logic; attribute dont_touch of G3086: signal is true;
	signal G3087: std_logic; attribute dont_touch of G3087: signal is true;
	signal G3088: std_logic; attribute dont_touch of G3088: signal is true;
	signal G3089: std_logic; attribute dont_touch of G3089: signal is true;
	signal G3092: std_logic; attribute dont_touch of G3092: signal is true;
	signal G3093: std_logic; attribute dont_touch of G3093: signal is true;
	signal G3094: std_logic; attribute dont_touch of G3094: signal is true;
	signal G3095: std_logic; attribute dont_touch of G3095: signal is true;
	signal G3096: std_logic; attribute dont_touch of G3096: signal is true;
	signal G3097: std_logic; attribute dont_touch of G3097: signal is true;
	signal G3098: std_logic; attribute dont_touch of G3098: signal is true;
	signal G3101: std_logic; attribute dont_touch of G3101: signal is true;
	signal G3102: std_logic; attribute dont_touch of G3102: signal is true;
	signal G3103: std_logic; attribute dont_touch of G3103: signal is true;
	signal G3104: std_logic; attribute dont_touch of G3104: signal is true;
	signal G3105: std_logic; attribute dont_touch of G3105: signal is true;
	signal G3106: std_logic; attribute dont_touch of G3106: signal is true;
	signal G3107: std_logic; attribute dont_touch of G3107: signal is true;
	signal G3108: std_logic; attribute dont_touch of G3108: signal is true;
	signal G3109: std_logic; attribute dont_touch of G3109: signal is true;
	signal G3110: std_logic; attribute dont_touch of G3110: signal is true;
	signal G3111: std_logic; attribute dont_touch of G3111: signal is true;
	signal G3112: std_logic; attribute dont_touch of G3112: signal is true;
	signal G3113: std_logic; attribute dont_touch of G3113: signal is true;
	signal G3118: std_logic; attribute dont_touch of G3118: signal is true;
	signal G3119: std_logic; attribute dont_touch of G3119: signal is true;
	signal G3120: std_logic; attribute dont_touch of G3120: signal is true;
	signal G3121: std_logic; attribute dont_touch of G3121: signal is true;
	signal G3138: std_logic; attribute dont_touch of G3138: signal is true;
	signal G3141: std_logic; attribute dont_touch of G3141: signal is true;
	signal G3142: std_logic; attribute dont_touch of G3142: signal is true;
	signal G3143: std_logic; attribute dont_touch of G3143: signal is true;
	signal G3144: std_logic; attribute dont_touch of G3144: signal is true;
	signal G3161: std_logic; attribute dont_touch of G3161: signal is true;
	signal G3164: std_logic; attribute dont_touch of G3164: signal is true;
	signal G3186: std_logic; attribute dont_touch of G3186: signal is true;
	signal G3200: std_logic; attribute dont_touch of G3200: signal is true;
	signal G3204: std_logic; attribute dont_touch of G3204: signal is true;
	signal G3205: std_logic; attribute dont_touch of G3205: signal is true;
	signal G3206: std_logic; attribute dont_touch of G3206: signal is true;
	signal G3207: std_logic; attribute dont_touch of G3207: signal is true;
	signal G3208: std_logic; attribute dont_touch of G3208: signal is true;
	signal G3209: std_logic; attribute dont_touch of G3209: signal is true;
	signal G3212: std_logic; attribute dont_touch of G3212: signal is true;
	signal G3213: std_logic; attribute dont_touch of G3213: signal is true;
	signal G3214: std_logic; attribute dont_touch of G3214: signal is true;
	signal G3215: std_logic; attribute dont_touch of G3215: signal is true;
	signal G3219: std_logic; attribute dont_touch of G3219: signal is true;
	signal G3220: std_logic; attribute dont_touch of G3220: signal is true;
	signal G3221: std_logic; attribute dont_touch of G3221: signal is true;
	signal G3222: std_logic; attribute dont_touch of G3222: signal is true;
	signal G3226: std_logic; attribute dont_touch of G3226: signal is true;
	signal G3227: std_logic; attribute dont_touch of G3227: signal is true;
	signal G3228: std_logic; attribute dont_touch of G3228: signal is true;
	signal G3246: std_logic; attribute dont_touch of G3246: signal is true;
	signal G3247: std_logic; attribute dont_touch of G3247: signal is true;
	signal G3252: std_logic; attribute dont_touch of G3252: signal is true;
	signal G3253: std_logic; attribute dont_touch of G3253: signal is true;
	signal G3254: std_logic; attribute dont_touch of G3254: signal is true;
	signal G3255: std_logic; attribute dont_touch of G3255: signal is true;
	signal G3256: std_logic; attribute dont_touch of G3256: signal is true;
	signal G3257: std_logic; attribute dont_touch of G3257: signal is true;
	signal G3260: std_logic; attribute dont_touch of G3260: signal is true;
	signal G3261: std_logic; attribute dont_touch of G3261: signal is true;
	signal G3262: std_logic; attribute dont_touch of G3262: signal is true;
	signal G3263: std_logic; attribute dont_touch of G3263: signal is true;
	signal G3266: std_logic; attribute dont_touch of G3266: signal is true;
	signal G3267: std_logic; attribute dont_touch of G3267: signal is true;
	signal G3268: std_logic; attribute dont_touch of G3268: signal is true;
	signal G3271: std_logic; attribute dont_touch of G3271: signal is true;
	signal G3272: std_logic; attribute dont_touch of G3272: signal is true;
	signal G3273: std_logic; attribute dont_touch of G3273: signal is true;
	signal G3274: std_logic; attribute dont_touch of G3274: signal is true;
	signal G3275: std_logic; attribute dont_touch of G3275: signal is true;
	signal G3281: std_logic; attribute dont_touch of G3281: signal is true;
	signal G3284: std_logic; attribute dont_touch of G3284: signal is true;
	signal G3287: std_logic; attribute dont_touch of G3287: signal is true;
	signal G3290: std_logic; attribute dont_touch of G3290: signal is true;
	signal G3291: std_logic; attribute dont_touch of G3291: signal is true;
	signal G3292: std_logic; attribute dont_touch of G3292: signal is true;
	signal G3301: std_logic; attribute dont_touch of G3301: signal is true;
	signal G3304: std_logic; attribute dont_touch of G3304: signal is true;
	signal G3305: std_logic; attribute dont_touch of G3305: signal is true;
	signal G3306: std_logic; attribute dont_touch of G3306: signal is true;
	signal G3307: std_logic; attribute dont_touch of G3307: signal is true;
	signal G3318: std_logic; attribute dont_touch of G3318: signal is true;
	signal G3321: std_logic; attribute dont_touch of G3321: signal is true;
	signal G3322: std_logic; attribute dont_touch of G3322: signal is true;
	signal G3323: std_logic; attribute dont_touch of G3323: signal is true;
	signal G3326: std_logic; attribute dont_touch of G3326: signal is true;
	signal G3328: std_logic; attribute dont_touch of G3328: signal is true;
	signal G3329: std_logic; attribute dont_touch of G3329: signal is true;
	signal G3330: std_logic; attribute dont_touch of G3330: signal is true;
	signal G3331: std_logic; attribute dont_touch of G3331: signal is true;
	signal G3332: std_logic; attribute dont_touch of G3332: signal is true;
	signal G3333: std_logic; attribute dont_touch of G3333: signal is true;
	signal G3334: std_logic; attribute dont_touch of G3334: signal is true;
	signal G3335: std_logic; attribute dont_touch of G3335: signal is true;
	signal G3336: std_logic; attribute dont_touch of G3336: signal is true;
	signal G3337: std_logic; attribute dont_touch of G3337: signal is true;
	signal G3343: std_logic; attribute dont_touch of G3343: signal is true;
	signal G3344: std_logic; attribute dont_touch of G3344: signal is true;
	signal G3345: std_logic; attribute dont_touch of G3345: signal is true;
	signal G3348: std_logic; attribute dont_touch of G3348: signal is true;
	signal G3351: std_logic; attribute dont_touch of G3351: signal is true;
	signal G3352: std_logic; attribute dont_touch of G3352: signal is true;
	signal G3353: std_logic; attribute dont_touch of G3353: signal is true;
	signal G3354: std_logic; attribute dont_touch of G3354: signal is true;
	signal G3359: std_logic; attribute dont_touch of G3359: signal is true;
	signal G3362: std_logic; attribute dont_touch of G3362: signal is true;
	signal G3363: std_logic; attribute dont_touch of G3363: signal is true;
	signal G3364: std_logic; attribute dont_touch of G3364: signal is true;
	signal G3365: std_logic; attribute dont_touch of G3365: signal is true;
	signal G3368: std_logic; attribute dont_touch of G3368: signal is true;
	signal G3369: std_logic; attribute dont_touch of G3369: signal is true;
	signal G3370: std_logic; attribute dont_touch of G3370: signal is true;
	signal G3371: std_logic; attribute dont_touch of G3371: signal is true;
	signal G3372: std_logic; attribute dont_touch of G3372: signal is true;
	signal G3373: std_logic; attribute dont_touch of G3373: signal is true;
	signal G3374: std_logic; attribute dont_touch of G3374: signal is true;
	signal G3375: std_logic; attribute dont_touch of G3375: signal is true;
	signal G3378: std_logic; attribute dont_touch of G3378: signal is true;
	signal G3379: std_logic; attribute dont_touch of G3379: signal is true;
	signal G3380: std_logic; attribute dont_touch of G3380: signal is true;
	signal G3381: std_logic; attribute dont_touch of G3381: signal is true;
	signal G3382: std_logic; attribute dont_touch of G3382: signal is true;
	signal G3383: std_logic; attribute dont_touch of G3383: signal is true;
	signal G3384: std_logic; attribute dont_touch of G3384: signal is true;
	signal G3385: std_logic; attribute dont_touch of G3385: signal is true;
	signal G3386: std_logic; attribute dont_touch of G3386: signal is true;
	signal G3387: std_logic; attribute dont_touch of G3387: signal is true;
	signal G3388: std_logic; attribute dont_touch of G3388: signal is true;
	signal G3389: std_logic; attribute dont_touch of G3389: signal is true;
	signal G3390: std_logic; attribute dont_touch of G3390: signal is true;
	signal G3391: std_logic; attribute dont_touch of G3391: signal is true;
	signal G3392: std_logic; attribute dont_touch of G3392: signal is true;
	signal G3393: std_logic; attribute dont_touch of G3393: signal is true;
	signal G3394: std_logic; attribute dont_touch of G3394: signal is true;
	signal G3395: std_logic; attribute dont_touch of G3395: signal is true;
	signal G3396: std_logic; attribute dont_touch of G3396: signal is true;
	signal G3397: std_logic; attribute dont_touch of G3397: signal is true;
	signal G3398: std_logic; attribute dont_touch of G3398: signal is true;
	signal G3399: std_logic; attribute dont_touch of G3399: signal is true;
	signal G3400: std_logic; attribute dont_touch of G3400: signal is true;
	signal G3404: std_logic; attribute dont_touch of G3404: signal is true;
	signal G3405: std_logic; attribute dont_touch of G3405: signal is true;
	signal G3406: std_logic; attribute dont_touch of G3406: signal is true;
	signal G3407: std_logic; attribute dont_touch of G3407: signal is true;
	signal G3408: std_logic; attribute dont_touch of G3408: signal is true;
	signal G3411: std_logic; attribute dont_touch of G3411: signal is true;
	signal G3412: std_logic; attribute dont_touch of G3412: signal is true;
	signal G3413: std_logic; attribute dont_touch of G3413: signal is true;
	signal G3414: std_logic; attribute dont_touch of G3414: signal is true;
	signal G3415: std_logic; attribute dont_touch of G3415: signal is true;
	signal G3416: std_logic; attribute dont_touch of G3416: signal is true;
	signal G3417: std_logic; attribute dont_touch of G3417: signal is true;
	signal G3418: std_logic; attribute dont_touch of G3418: signal is true;
	signal G3419: std_logic; attribute dont_touch of G3419: signal is true;
	signal G3422: std_logic; attribute dont_touch of G3422: signal is true;
	signal G3423: std_logic; attribute dont_touch of G3423: signal is true;
	signal G3424: std_logic; attribute dont_touch of G3424: signal is true;
	signal G3425: std_logic; attribute dont_touch of G3425: signal is true;
	signal G3426: std_logic; attribute dont_touch of G3426: signal is true;
	signal G3427: std_logic; attribute dont_touch of G3427: signal is true;
	signal G3428: std_logic; attribute dont_touch of G3428: signal is true;
	signal G3429: std_logic; attribute dont_touch of G3429: signal is true;
	signal G3430: std_logic; attribute dont_touch of G3430: signal is true;
	signal G3431: std_logic; attribute dont_touch of G3431: signal is true;
	signal G3432: std_logic; attribute dont_touch of G3432: signal is true;
	signal G3433: std_logic; attribute dont_touch of G3433: signal is true;
	signal G3434: std_logic; attribute dont_touch of G3434: signal is true;
	signal G3435: std_logic; attribute dont_touch of G3435: signal is true;
	signal G3436: std_logic; attribute dont_touch of G3436: signal is true;
	signal G3437: std_logic; attribute dont_touch of G3437: signal is true;
	signal G3438: std_logic; attribute dont_touch of G3438: signal is true;
	signal G3439: std_logic; attribute dont_touch of G3439: signal is true;
	signal G3440: std_logic; attribute dont_touch of G3440: signal is true;
	signal G3458: std_logic; attribute dont_touch of G3458: signal is true;
	signal G3459: std_logic; attribute dont_touch of G3459: signal is true;
	signal G3460: std_logic; attribute dont_touch of G3460: signal is true;
	signal G3461: std_logic; attribute dont_touch of G3461: signal is true;
	signal G3462: std_logic; attribute dont_touch of G3462: signal is true;
	signal G3463: std_logic; attribute dont_touch of G3463: signal is true;
	signal G3473: std_logic; attribute dont_touch of G3473: signal is true;
	signal G3474: std_logic; attribute dont_touch of G3474: signal is true;
	signal G3475: std_logic; attribute dont_touch of G3475: signal is true;
	signal G3479: std_logic; attribute dont_touch of G3479: signal is true;
	signal G3485: std_logic; attribute dont_touch of G3485: signal is true;
	signal G3491: std_logic; attribute dont_touch of G3491: signal is true;
	signal G3496: std_logic; attribute dont_touch of G3496: signal is true;
	signal G3497: std_logic; attribute dont_touch of G3497: signal is true;
	signal G3500: std_logic; attribute dont_touch of G3500: signal is true;
	signal G3501: std_logic; attribute dont_touch of G3501: signal is true;
	signal G3505: std_logic; attribute dont_touch of G3505: signal is true;
	signal G3506: std_logic; attribute dont_touch of G3506: signal is true;
	signal G3507: std_logic; attribute dont_touch of G3507: signal is true;
	signal G3512: std_logic; attribute dont_touch of G3512: signal is true;
	signal G3513: std_logic; attribute dont_touch of G3513: signal is true;
	signal G3516: std_logic; attribute dont_touch of G3516: signal is true;
	signal G3517: std_logic; attribute dont_touch of G3517: signal is true;
	signal G3518: std_logic; attribute dont_touch of G3518: signal is true;
	signal G3519: std_logic; attribute dont_touch of G3519: signal is true;
	signal G3520: std_logic; attribute dont_touch of G3520: signal is true;
	signal G3521: std_logic; attribute dont_touch of G3521: signal is true;
	signal G3522: std_logic; attribute dont_touch of G3522: signal is true;
	signal G3523: std_logic; attribute dont_touch of G3523: signal is true;
	signal G3524: std_logic; attribute dont_touch of G3524: signal is true;
	signal G3528: std_logic; attribute dont_touch of G3528: signal is true;
	signal G3529: std_logic; attribute dont_touch of G3529: signal is true;
	signal G3530: std_logic; attribute dont_touch of G3530: signal is true;
	signal G3531: std_logic; attribute dont_touch of G3531: signal is true;
	signal G3532: std_logic; attribute dont_touch of G3532: signal is true;
	signal G3533: std_logic; attribute dont_touch of G3533: signal is true;
	signal G3536: std_logic; attribute dont_touch of G3536: signal is true;
	signal G3537: std_logic; attribute dont_touch of G3537: signal is true;
	signal G3538: std_logic; attribute dont_touch of G3538: signal is true;
	signal G3539: std_logic; attribute dont_touch of G3539: signal is true;
	signal G3540: std_logic; attribute dont_touch of G3540: signal is true;
	signal G3543: std_logic; attribute dont_touch of G3543: signal is true;
	signal G3544: std_logic; attribute dont_touch of G3544: signal is true;
	signal G3545: std_logic; attribute dont_touch of G3545: signal is true;
	signal G3546: std_logic; attribute dont_touch of G3546: signal is true;
	signal G3563: std_logic; attribute dont_touch of G3563: signal is true;
	signal G3566: std_logic; attribute dont_touch of G3566: signal is true;
	signal G3582: std_logic; attribute dont_touch of G3582: signal is true;
	signal G3583: std_logic; attribute dont_touch of G3583: signal is true;
	signal G3584: std_logic; attribute dont_touch of G3584: signal is true;
	signal G3585: std_logic; attribute dont_touch of G3585: signal is true;
	signal G3586: std_logic; attribute dont_touch of G3586: signal is true;
	signal G3621: std_logic; attribute dont_touch of G3621: signal is true;
	signal G3622: std_logic; attribute dont_touch of G3622: signal is true;
	signal G3623: std_logic; attribute dont_touch of G3623: signal is true;
	signal G3624: std_logic; attribute dont_touch of G3624: signal is true;
	signal G3625: std_logic; attribute dont_touch of G3625: signal is true;
	signal G3626: std_logic; attribute dont_touch of G3626: signal is true;
	signal G3627: std_logic; attribute dont_touch of G3627: signal is true;
	signal G3628: std_logic; attribute dont_touch of G3628: signal is true;
	signal G3629: std_logic; attribute dont_touch of G3629: signal is true;
	signal G3630: std_logic; attribute dont_touch of G3630: signal is true;
	signal G3631: std_logic; attribute dont_touch of G3631: signal is true;
	signal G3632: std_logic; attribute dont_touch of G3632: signal is true;
	signal G3633: std_logic; attribute dont_touch of G3633: signal is true;
	signal G3634: std_logic; attribute dont_touch of G3634: signal is true;
	signal G3635: std_logic; attribute dont_touch of G3635: signal is true;
	signal G3636: std_logic; attribute dont_touch of G3636: signal is true;
	signal G3637: std_logic; attribute dont_touch of G3637: signal is true;
	signal G3638: std_logic; attribute dont_touch of G3638: signal is true;
	signal G3661: std_logic; attribute dont_touch of G3661: signal is true;
	signal G3662: std_logic; attribute dont_touch of G3662: signal is true;
	signal G3663: std_logic; attribute dont_touch of G3663: signal is true;
	signal G3664: std_logic; attribute dont_touch of G3664: signal is true;
	signal G3681: std_logic; attribute dont_touch of G3681: signal is true;
	signal G3682: std_logic; attribute dont_touch of G3682: signal is true;
	signal G3683: std_logic; attribute dont_touch of G3683: signal is true;
	signal G3684: std_logic; attribute dont_touch of G3684: signal is true;
	signal G3685: std_logic; attribute dont_touch of G3685: signal is true;
	signal G3688: std_logic; attribute dont_touch of G3688: signal is true;
	signal G3693: std_logic; attribute dont_touch of G3693: signal is true;
	signal G3694: std_logic; attribute dont_touch of G3694: signal is true;
	signal G3695: std_logic; attribute dont_touch of G3695: signal is true;
	signal G3696: std_logic; attribute dont_touch of G3696: signal is true;
	signal G3697: std_logic; attribute dont_touch of G3697: signal is true;
	signal G3698: std_logic; attribute dont_touch of G3698: signal is true;
	signal G3703: std_logic; attribute dont_touch of G3703: signal is true;
	signal G3704: std_logic; attribute dont_touch of G3704: signal is true;
	signal G3705: std_logic; attribute dont_touch of G3705: signal is true;
	signal G3706: std_logic; attribute dont_touch of G3706: signal is true;
	signal G3707: std_logic; attribute dont_touch of G3707: signal is true;
	signal G3708: std_logic; attribute dont_touch of G3708: signal is true;
	signal G3709: std_logic; attribute dont_touch of G3709: signal is true;
	signal G3710: std_logic; attribute dont_touch of G3710: signal is true;
	signal G3714: std_logic; attribute dont_touch of G3714: signal is true;
	signal G3715: std_logic; attribute dont_touch of G3715: signal is true;
	signal G3716: std_logic; attribute dont_touch of G3716: signal is true;
	signal G3717: std_logic; attribute dont_touch of G3717: signal is true;
	signal G3718: std_logic; attribute dont_touch of G3718: signal is true;
	signal G3719: std_logic; attribute dont_touch of G3719: signal is true;
	signal G3720: std_logic; attribute dont_touch of G3720: signal is true;
	signal G3721: std_logic; attribute dont_touch of G3721: signal is true;
	signal G3722: std_logic; attribute dont_touch of G3722: signal is true;
	signal G3723: std_logic; attribute dont_touch of G3723: signal is true;
	signal G3726: std_logic; attribute dont_touch of G3726: signal is true;
	signal G3727: std_logic; attribute dont_touch of G3727: signal is true;
	signal G3728: std_logic; attribute dont_touch of G3728: signal is true;
	signal G3729: std_logic; attribute dont_touch of G3729: signal is true;
	signal G3730: std_logic; attribute dont_touch of G3730: signal is true;
	signal G3731: std_logic; attribute dont_touch of G3731: signal is true;
	signal G3732: std_logic; attribute dont_touch of G3732: signal is true;
	signal G3733: std_logic; attribute dont_touch of G3733: signal is true;
	signal G3734: std_logic; attribute dont_touch of G3734: signal is true;
	signal G3735: std_logic; attribute dont_touch of G3735: signal is true;
	signal G3736: std_logic; attribute dont_touch of G3736: signal is true;
	signal G3737: std_logic; attribute dont_touch of G3737: signal is true;
	signal G3738: std_logic; attribute dont_touch of G3738: signal is true;
	signal G3742: std_logic; attribute dont_touch of G3742: signal is true;
	signal G3743: std_logic; attribute dont_touch of G3743: signal is true;
	signal G3744: std_logic; attribute dont_touch of G3744: signal is true;
	signal G3747: std_logic; attribute dont_touch of G3747: signal is true;
	signal G3748: std_logic; attribute dont_touch of G3748: signal is true;
	signal G3749: std_logic; attribute dont_touch of G3749: signal is true;
	signal G3750: std_logic; attribute dont_touch of G3750: signal is true;
	signal G3751: std_logic; attribute dont_touch of G3751: signal is true;
	signal G3752: std_logic; attribute dont_touch of G3752: signal is true;
	signal G3753: std_logic; attribute dont_touch of G3753: signal is true;
	signal G3756: std_logic; attribute dont_touch of G3756: signal is true;
	signal G3757: std_logic; attribute dont_touch of G3757: signal is true;
	signal G3758: std_logic; attribute dont_touch of G3758: signal is true;
	signal G3759: std_logic; attribute dont_touch of G3759: signal is true;
	signal G3760: std_logic; attribute dont_touch of G3760: signal is true;
	signal G3761: std_logic; attribute dont_touch of G3761: signal is true;
	signal G3762: std_logic; attribute dont_touch of G3762: signal is true;
	signal G3763: std_logic; attribute dont_touch of G3763: signal is true;
	signal G3764: std_logic; attribute dont_touch of G3764: signal is true;
	signal G3765: std_logic; attribute dont_touch of G3765: signal is true;
	signal G3766: std_logic; attribute dont_touch of G3766: signal is true;
	signal G3767: std_logic; attribute dont_touch of G3767: signal is true;
	signal G3768: std_logic; attribute dont_touch of G3768: signal is true;
	signal G3769: std_logic; attribute dont_touch of G3769: signal is true;
	signal G3770: std_logic; attribute dont_touch of G3770: signal is true;
	signal G3771: std_logic; attribute dont_touch of G3771: signal is true;
	signal G3772: std_logic; attribute dont_touch of G3772: signal is true;
	signal G3773: std_logic; attribute dont_touch of G3773: signal is true;
	signal G3774: std_logic; attribute dont_touch of G3774: signal is true;
	signal G3775: std_logic; attribute dont_touch of G3775: signal is true;
	signal G3776: std_logic; attribute dont_touch of G3776: signal is true;
	signal G3782: std_logic; attribute dont_touch of G3782: signal is true;
	signal G3783: std_logic; attribute dont_touch of G3783: signal is true;
	signal G3784: std_logic; attribute dont_touch of G3784: signal is true;
	signal G3790: std_logic; attribute dont_touch of G3790: signal is true;
	signal G3791: std_logic; attribute dont_touch of G3791: signal is true;
	signal G3792: std_logic; attribute dont_touch of G3792: signal is true;
	signal G3793: std_logic; attribute dont_touch of G3793: signal is true;
	signal G3798: std_logic; attribute dont_touch of G3798: signal is true;
	signal G3799: std_logic; attribute dont_touch of G3799: signal is true;
	signal G3800: std_logic; attribute dont_touch of G3800: signal is true;
	signal G3804: std_logic; attribute dont_touch of G3804: signal is true;
	signal G3807: std_logic; attribute dont_touch of G3807: signal is true;
	signal G3810: std_logic; attribute dont_touch of G3810: signal is true;
	signal G3811: std_logic; attribute dont_touch of G3811: signal is true;
	signal G3812: std_logic; attribute dont_touch of G3812: signal is true;
	signal G3813: std_logic; attribute dont_touch of G3813: signal is true;
	signal G3814: std_logic; attribute dont_touch of G3814: signal is true;
	signal G3815: std_logic; attribute dont_touch of G3815: signal is true;
	signal G3816: std_logic; attribute dont_touch of G3816: signal is true;
	signal G3817: std_logic; attribute dont_touch of G3817: signal is true;
	signal G3818: std_logic; attribute dont_touch of G3818: signal is true;
	signal G3819: std_logic; attribute dont_touch of G3819: signal is true;
	signal G3820: std_logic; attribute dont_touch of G3820: signal is true;
	signal G3828: std_logic; attribute dont_touch of G3828: signal is true;
	signal G3829: std_logic; attribute dont_touch of G3829: signal is true;
	signal G3860: std_logic; attribute dont_touch of G3860: signal is true;
	signal G3861: std_logic; attribute dont_touch of G3861: signal is true;
	signal G3862: std_logic; attribute dont_touch of G3862: signal is true;
	signal G3863: std_logic; attribute dont_touch of G3863: signal is true;
	signal G3874: std_logic; attribute dont_touch of G3874: signal is true;
	signal G3875: std_logic; attribute dont_touch of G3875: signal is true;
	signal G3876: std_logic; attribute dont_touch of G3876: signal is true;
	signal G3877: std_logic; attribute dont_touch of G3877: signal is true;
	signal G3878: std_logic; attribute dont_touch of G3878: signal is true;
	signal G3879: std_logic; attribute dont_touch of G3879: signal is true;
	signal G3880: std_logic; attribute dont_touch of G3880: signal is true;
	signal G3903: std_logic; attribute dont_touch of G3903: signal is true;
	signal G3904: std_logic; attribute dont_touch of G3904: signal is true;
	signal G3905: std_logic; attribute dont_touch of G3905: signal is true;
	signal G3906: std_logic; attribute dont_touch of G3906: signal is true;
	signal G3907: std_logic; attribute dont_touch of G3907: signal is true;
	signal G3908: std_logic; attribute dont_touch of G3908: signal is true;
	signal G3909: std_logic; attribute dont_touch of G3909: signal is true;
	signal G3910: std_logic; attribute dont_touch of G3910: signal is true;
	signal G3911: std_logic; attribute dont_touch of G3911: signal is true;
	signal G3912: std_logic; attribute dont_touch of G3912: signal is true;
	signal G3913: std_logic; attribute dont_touch of G3913: signal is true;
	signal G3914: std_logic; attribute dont_touch of G3914: signal is true;
	signal G3937: std_logic; attribute dont_touch of G3937: signal is true;
	signal G3938: std_logic; attribute dont_touch of G3938: signal is true;
	signal G3939: std_logic; attribute dont_touch of G3939: signal is true;
	signal G3940: std_logic; attribute dont_touch of G3940: signal is true;
	signal G3941: std_logic; attribute dont_touch of G3941: signal is true;
	signal G3942: std_logic; attribute dont_touch of G3942: signal is true;
	signal G3943: std_logic; attribute dont_touch of G3943: signal is true;
	signal G3944: std_logic; attribute dont_touch of G3944: signal is true;
	signal G3945: std_logic; attribute dont_touch of G3945: signal is true;
	signal G3946: std_logic; attribute dont_touch of G3946: signal is true;
	signal G3967: std_logic; attribute dont_touch of G3967: signal is true;
	signal G3970: std_logic; attribute dont_touch of G3970: signal is true;
	signal G3971: std_logic; attribute dont_touch of G3971: signal is true;
	signal G3974: std_logic; attribute dont_touch of G3974: signal is true;
	signal G3975: std_logic; attribute dont_touch of G3975: signal is true;
	signal G3976: std_logic; attribute dont_touch of G3976: signal is true;
	signal G3977: std_logic; attribute dont_touch of G3977: signal is true;
	signal G3978: std_logic; attribute dont_touch of G3978: signal is true;
	signal G3979: std_logic; attribute dont_touch of G3979: signal is true;
	signal G3980: std_logic; attribute dont_touch of G3980: signal is true;
	signal G3981: std_logic; attribute dont_touch of G3981: signal is true;
	signal G3982: std_logic; attribute dont_touch of G3982: signal is true;
	signal G3983: std_logic; attribute dont_touch of G3983: signal is true;
	signal G3987: std_logic; attribute dont_touch of G3987: signal is true;
	signal G3988: std_logic; attribute dont_touch of G3988: signal is true;
	signal G3989: std_logic; attribute dont_touch of G3989: signal is true;
	signal G3990: std_logic; attribute dont_touch of G3990: signal is true;
	signal G3991: std_logic; attribute dont_touch of G3991: signal is true;
	signal G3992: std_logic; attribute dont_touch of G3992: signal is true;
	signal G3995: std_logic; attribute dont_touch of G3995: signal is true;
	signal G3996: std_logic; attribute dont_touch of G3996: signal is true;
	signal G3997: std_logic; attribute dont_touch of G3997: signal is true;
	signal G3998: std_logic; attribute dont_touch of G3998: signal is true;
	signal G3999: std_logic; attribute dont_touch of G3999: signal is true;
	signal G4000: std_logic; attribute dont_touch of G4000: signal is true;
	signal G4001: std_logic; attribute dont_touch of G4001: signal is true;
	signal G4002: std_logic; attribute dont_touch of G4002: signal is true;
	signal G4003: std_logic; attribute dont_touch of G4003: signal is true;
	signal G4004: std_logic; attribute dont_touch of G4004: signal is true;
	signal G4005: std_logic; attribute dont_touch of G4005: signal is true;
	signal G4006: std_logic; attribute dont_touch of G4006: signal is true;
	signal G4007: std_logic; attribute dont_touch of G4007: signal is true;
	signal G4008: std_logic; attribute dont_touch of G4008: signal is true;
	signal G4009: std_logic; attribute dont_touch of G4009: signal is true;
	signal G4010: std_logic; attribute dont_touch of G4010: signal is true;
	signal G4011: std_logic; attribute dont_touch of G4011: signal is true;
	signal G4012: std_logic; attribute dont_touch of G4012: signal is true;
	signal G4013: std_logic; attribute dont_touch of G4013: signal is true;
	signal G4047: std_logic; attribute dont_touch of G4047: signal is true;
	signal G4048: std_logic; attribute dont_touch of G4048: signal is true;
	signal G4049: std_logic; attribute dont_touch of G4049: signal is true;
	signal G4050: std_logic; attribute dont_touch of G4050: signal is true;
	signal G4051: std_logic; attribute dont_touch of G4051: signal is true;
	signal G4052: std_logic; attribute dont_touch of G4052: signal is true;
	signal G4053: std_logic; attribute dont_touch of G4053: signal is true;
	signal G4054: std_logic; attribute dont_touch of G4054: signal is true;
	signal G4055: std_logic; attribute dont_touch of G4055: signal is true;
	signal G4056: std_logic; attribute dont_touch of G4056: signal is true;
	signal G4057: std_logic; attribute dont_touch of G4057: signal is true;
	signal G4058: std_logic; attribute dont_touch of G4058: signal is true;
	signal G4059: std_logic; attribute dont_touch of G4059: signal is true;
	signal G4060: std_logic; attribute dont_touch of G4060: signal is true;
	signal G4061: std_logic; attribute dont_touch of G4061: signal is true;
	signal G4062: std_logic; attribute dont_touch of G4062: signal is true;
	signal G4063: std_logic; attribute dont_touch of G4063: signal is true;
	signal G4064: std_logic; attribute dont_touch of G4064: signal is true;
	signal G4065: std_logic; attribute dont_touch of G4065: signal is true;
	signal G4066: std_logic; attribute dont_touch of G4066: signal is true;
	signal G4067: std_logic; attribute dont_touch of G4067: signal is true;
	signal G4068: std_logic; attribute dont_touch of G4068: signal is true;
	signal G4069: std_logic; attribute dont_touch of G4069: signal is true;
	signal G4070: std_logic; attribute dont_touch of G4070: signal is true;
	signal G4073: std_logic; attribute dont_touch of G4073: signal is true;
	signal G4076: std_logic; attribute dont_touch of G4076: signal is true;
	signal G4077: std_logic; attribute dont_touch of G4077: signal is true;
	signal G4078: std_logic; attribute dont_touch of G4078: signal is true;
	signal G4079: std_logic; attribute dont_touch of G4079: signal is true;
	signal G4080: std_logic; attribute dont_touch of G4080: signal is true;
	signal G4081: std_logic; attribute dont_touch of G4081: signal is true;
	signal G4082: std_logic; attribute dont_touch of G4082: signal is true;
	signal G4083: std_logic; attribute dont_touch of G4083: signal is true;
	signal G4084: std_logic; attribute dont_touch of G4084: signal is true;
	signal G4087: std_logic; attribute dont_touch of G4087: signal is true;
	signal G4088: std_logic; attribute dont_touch of G4088: signal is true;
	signal G4089: std_logic; attribute dont_touch of G4089: signal is true;
	signal G4093: std_logic; attribute dont_touch of G4093: signal is true;
	signal G4094: std_logic; attribute dont_touch of G4094: signal is true;
	signal G4095: std_logic; attribute dont_touch of G4095: signal is true;
	signal G4096: std_logic; attribute dont_touch of G4096: signal is true;
	signal G4097: std_logic; attribute dont_touch of G4097: signal is true;
	signal G4098: std_logic; attribute dont_touch of G4098: signal is true;
	signal G4099: std_logic; attribute dont_touch of G4099: signal is true;
	signal G4102: std_logic; attribute dont_touch of G4102: signal is true;
	signal G4103: std_logic; attribute dont_touch of G4103: signal is true;
	signal G4104: std_logic; attribute dont_touch of G4104: signal is true;
	signal G4105: std_logic; attribute dont_touch of G4105: signal is true;
	signal G4106: std_logic; attribute dont_touch of G4106: signal is true;
	signal G4109: std_logic; attribute dont_touch of G4109: signal is true;
	signal G4112: std_logic; attribute dont_touch of G4112: signal is true;
	signal G4113: std_logic; attribute dont_touch of G4113: signal is true;
	signal G4114: std_logic; attribute dont_touch of G4114: signal is true;
	signal G4115: std_logic; attribute dont_touch of G4115: signal is true;
	signal G4116: std_logic; attribute dont_touch of G4116: signal is true;
	signal G4117: std_logic; attribute dont_touch of G4117: signal is true;
	signal G4121: std_logic; attribute dont_touch of G4121: signal is true;
	signal G4122: std_logic; attribute dont_touch of G4122: signal is true;
	signal G4123: std_logic; attribute dont_touch of G4123: signal is true;
	signal G4124: std_logic; attribute dont_touch of G4124: signal is true;
	signal G4125: std_logic; attribute dont_touch of G4125: signal is true;
	signal G4126: std_logic; attribute dont_touch of G4126: signal is true;
	signal G4127: std_logic; attribute dont_touch of G4127: signal is true;
	signal G4128: std_logic; attribute dont_touch of G4128: signal is true;
	signal G4129: std_logic; attribute dont_touch of G4129: signal is true;
	signal G4130: std_logic; attribute dont_touch of G4130: signal is true;
	signal G4140: std_logic; attribute dont_touch of G4140: signal is true;
	signal G4141: std_logic; attribute dont_touch of G4141: signal is true;
	signal G4142: std_logic; attribute dont_touch of G4142: signal is true;
	signal G4143: std_logic; attribute dont_touch of G4143: signal is true;
	signal G4144: std_logic; attribute dont_touch of G4144: signal is true;
	signal G4156: std_logic; attribute dont_touch of G4156: signal is true;
	signal G4157: std_logic; attribute dont_touch of G4157: signal is true;
	signal G4158: std_logic; attribute dont_touch of G4158: signal is true;
	signal G4159: std_logic; attribute dont_touch of G4159: signal is true;
	signal G4160: std_logic; attribute dont_touch of G4160: signal is true;
	signal G4161: std_logic; attribute dont_touch of G4161: signal is true;
	signal G4162: std_logic; attribute dont_touch of G4162: signal is true;
	signal G4163: std_logic; attribute dont_touch of G4163: signal is true;
	signal G4164: std_logic; attribute dont_touch of G4164: signal is true;
	signal G4165: std_logic; attribute dont_touch of G4165: signal is true;
	signal G4166: std_logic; attribute dont_touch of G4166: signal is true;
	signal G4167: std_logic; attribute dont_touch of G4167: signal is true;
	signal G4168: std_logic; attribute dont_touch of G4168: signal is true;
	signal G4169: std_logic; attribute dont_touch of G4169: signal is true;
	signal G4170: std_logic; attribute dont_touch of G4170: signal is true;
	signal G4182: std_logic; attribute dont_touch of G4182: signal is true;
	signal G4183: std_logic; attribute dont_touch of G4183: signal is true;
	signal G4184: std_logic; attribute dont_touch of G4184: signal is true;
	signal G4185: std_logic; attribute dont_touch of G4185: signal is true;
	signal G4186: std_logic; attribute dont_touch of G4186: signal is true;
	signal G4187: std_logic; attribute dont_touch of G4187: signal is true;
	signal G4188: std_logic; attribute dont_touch of G4188: signal is true;
	signal G4189: std_logic; attribute dont_touch of G4189: signal is true;
	signal G4190: std_logic; attribute dont_touch of G4190: signal is true;
	signal G4217: std_logic; attribute dont_touch of G4217: signal is true;
	signal G4218: std_logic; attribute dont_touch of G4218: signal is true;
	signal G4219: std_logic; attribute dont_touch of G4219: signal is true;
	signal G4220: std_logic; attribute dont_touch of G4220: signal is true;
	signal G4221: std_logic; attribute dont_touch of G4221: signal is true;
	signal G4222: std_logic; attribute dont_touch of G4222: signal is true;
	signal G4223: std_logic; attribute dont_touch of G4223: signal is true;
	signal G4224: std_logic; attribute dont_touch of G4224: signal is true;
	signal G4225: std_logic; attribute dont_touch of G4225: signal is true;
	signal G4226: std_logic; attribute dont_touch of G4226: signal is true;
	signal G4227: std_logic; attribute dont_touch of G4227: signal is true;
	signal G4228: std_logic; attribute dont_touch of G4228: signal is true;
	signal G4229: std_logic; attribute dont_touch of G4229: signal is true;
	signal G4230: std_logic; attribute dont_touch of G4230: signal is true;
	signal G4231: std_logic; attribute dont_touch of G4231: signal is true;
	signal G4232: std_logic; attribute dont_touch of G4232: signal is true;
	signal G4233: std_logic; attribute dont_touch of G4233: signal is true;
	signal G4234: std_logic; attribute dont_touch of G4234: signal is true;
	signal G4235: std_logic; attribute dont_touch of G4235: signal is true;
	signal G4236: std_logic; attribute dont_touch of G4236: signal is true;
	signal G4237: std_logic; attribute dont_touch of G4237: signal is true;
	signal G4238: std_logic; attribute dont_touch of G4238: signal is true;
	signal G4239: std_logic; attribute dont_touch of G4239: signal is true;
	signal G4240: std_logic; attribute dont_touch of G4240: signal is true;
	signal G4241: std_logic; attribute dont_touch of G4241: signal is true;
	signal G4242: std_logic; attribute dont_touch of G4242: signal is true;
	signal G4243: std_logic; attribute dont_touch of G4243: signal is true;
	signal G4250: std_logic; attribute dont_touch of G4250: signal is true;
	signal G4251: std_logic; attribute dont_touch of G4251: signal is true;
	signal G4252: std_logic; attribute dont_touch of G4252: signal is true;
	signal G4253: std_logic; attribute dont_touch of G4253: signal is true;
	signal G4254: std_logic; attribute dont_touch of G4254: signal is true;
	signal G4255: std_logic; attribute dont_touch of G4255: signal is true;
	signal G4256: std_logic; attribute dont_touch of G4256: signal is true;
	signal G4257: std_logic; attribute dont_touch of G4257: signal is true;
	signal G4258: std_logic; attribute dont_touch of G4258: signal is true;
	signal G4259: std_logic; attribute dont_touch of G4259: signal is true;
	signal G4260: std_logic; attribute dont_touch of G4260: signal is true;
	signal G4261: std_logic; attribute dont_touch of G4261: signal is true;
	signal G4262: std_logic; attribute dont_touch of G4262: signal is true;
	signal G4263: std_logic; attribute dont_touch of G4263: signal is true;
	signal G4264: std_logic; attribute dont_touch of G4264: signal is true;
	signal G4265: std_logic; attribute dont_touch of G4265: signal is true;
	signal G4266: std_logic; attribute dont_touch of G4266: signal is true;
	signal G4267: std_logic; attribute dont_touch of G4267: signal is true;
	signal G4268: std_logic; attribute dont_touch of G4268: signal is true;
	signal G4269: std_logic; attribute dont_touch of G4269: signal is true;
	signal G4270: std_logic; attribute dont_touch of G4270: signal is true;
	signal G4271: std_logic; attribute dont_touch of G4271: signal is true;
	signal G4272: std_logic; attribute dont_touch of G4272: signal is true;
	signal G4273: std_logic; attribute dont_touch of G4273: signal is true;
	signal G4274: std_logic; attribute dont_touch of G4274: signal is true;
	signal G4275: std_logic; attribute dont_touch of G4275: signal is true;
	signal G4276: std_logic; attribute dont_touch of G4276: signal is true;
	signal G4277: std_logic; attribute dont_touch of G4277: signal is true;
	signal G4278: std_logic; attribute dont_touch of G4278: signal is true;
	signal G4279: std_logic; attribute dont_touch of G4279: signal is true;
	signal G4280: std_logic; attribute dont_touch of G4280: signal is true;
	signal G4281: std_logic; attribute dont_touch of G4281: signal is true;
	signal G4282: std_logic; attribute dont_touch of G4282: signal is true;
	signal G4283: std_logic; attribute dont_touch of G4283: signal is true;
	signal G4284: std_logic; attribute dont_touch of G4284: signal is true;
	signal G4285: std_logic; attribute dont_touch of G4285: signal is true;
	signal G4286: std_logic; attribute dont_touch of G4286: signal is true;
	signal G4287: std_logic; attribute dont_touch of G4287: signal is true;
	signal G4288: std_logic; attribute dont_touch of G4288: signal is true;
	signal G4289: std_logic; attribute dont_touch of G4289: signal is true;
	signal G4290: std_logic; attribute dont_touch of G4290: signal is true;
	signal G4291: std_logic; attribute dont_touch of G4291: signal is true;
	signal G4292: std_logic; attribute dont_touch of G4292: signal is true;
	signal G4293: std_logic; attribute dont_touch of G4293: signal is true;
	signal G4294: std_logic; attribute dont_touch of G4294: signal is true;
	signal G4295: std_logic; attribute dont_touch of G4295: signal is true;
	signal G4296: std_logic; attribute dont_touch of G4296: signal is true;
	signal G4297: std_logic; attribute dont_touch of G4297: signal is true;
	signal G4298: std_logic; attribute dont_touch of G4298: signal is true;
	signal G4299: std_logic; attribute dont_touch of G4299: signal is true;
	signal G4300: std_logic; attribute dont_touch of G4300: signal is true;
	signal G4305: std_logic; attribute dont_touch of G4305: signal is true;
	signal G4306: std_logic; attribute dont_touch of G4306: signal is true;
	signal G4307: std_logic; attribute dont_touch of G4307: signal is true;
	signal G4308: std_logic; attribute dont_touch of G4308: signal is true;
	signal G4309: std_logic; attribute dont_touch of G4309: signal is true;
	signal G4310: std_logic; attribute dont_touch of G4310: signal is true;
	signal G4311: std_logic; attribute dont_touch of G4311: signal is true;
	signal G4312: std_logic; attribute dont_touch of G4312: signal is true;
	signal G4313: std_logic; attribute dont_touch of G4313: signal is true;
	signal G4314: std_logic; attribute dont_touch of G4314: signal is true;
	signal G4315: std_logic; attribute dont_touch of G4315: signal is true;
	signal G4316: std_logic; attribute dont_touch of G4316: signal is true;
	signal G4317: std_logic; attribute dont_touch of G4317: signal is true;
	signal G4318: std_logic; attribute dont_touch of G4318: signal is true;
	signal G4319: std_logic; attribute dont_touch of G4319: signal is true;
	signal G4320: std_logic; attribute dont_touch of G4320: signal is true;
	signal G4321: std_logic; attribute dont_touch of G4321: signal is true;
	signal G4322: std_logic; attribute dont_touch of G4322: signal is true;
	signal G4323: std_logic; attribute dont_touch of G4323: signal is true;
	signal G4324: std_logic; attribute dont_touch of G4324: signal is true;
	signal G4325: std_logic; attribute dont_touch of G4325: signal is true;
	signal G4326: std_logic; attribute dont_touch of G4326: signal is true;
	signal G4327: std_logic; attribute dont_touch of G4327: signal is true;
	signal G4328: std_logic; attribute dont_touch of G4328: signal is true;
	signal G4329: std_logic; attribute dont_touch of G4329: signal is true;
	signal G4330: std_logic; attribute dont_touch of G4330: signal is true;
	signal G4331: std_logic; attribute dont_touch of G4331: signal is true;
	signal G4332: std_logic; attribute dont_touch of G4332: signal is true;
	signal G4333: std_logic; attribute dont_touch of G4333: signal is true;
	signal G4334: std_logic; attribute dont_touch of G4334: signal is true;
	signal G4335: std_logic; attribute dont_touch of G4335: signal is true;
	signal G4336: std_logic; attribute dont_touch of G4336: signal is true;
	signal G4337: std_logic; attribute dont_touch of G4337: signal is true;
	signal G4338: std_logic; attribute dont_touch of G4338: signal is true;
	signal G4339: std_logic; attribute dont_touch of G4339: signal is true;
	signal G4340: std_logic; attribute dont_touch of G4340: signal is true;
	signal G4341: std_logic; attribute dont_touch of G4341: signal is true;
	signal G4342: std_logic; attribute dont_touch of G4342: signal is true;
	signal G4343: std_logic; attribute dont_touch of G4343: signal is true;
	signal G4344: std_logic; attribute dont_touch of G4344: signal is true;
	signal G4345: std_logic; attribute dont_touch of G4345: signal is true;
	signal G4346: std_logic; attribute dont_touch of G4346: signal is true;
	signal G4347: std_logic; attribute dont_touch of G4347: signal is true;
	signal G4348: std_logic; attribute dont_touch of G4348: signal is true;
	signal G4351: std_logic; attribute dont_touch of G4351: signal is true;
	signal G4352: std_logic; attribute dont_touch of G4352: signal is true;
	signal G4353: std_logic; attribute dont_touch of G4353: signal is true;
	signal G4354: std_logic; attribute dont_touch of G4354: signal is true;
	signal G4355: std_logic; attribute dont_touch of G4355: signal is true;
	signal G4358: std_logic; attribute dont_touch of G4358: signal is true;
	signal G4359: std_logic; attribute dont_touch of G4359: signal is true;
	signal G4360: std_logic; attribute dont_touch of G4360: signal is true;
	signal G4361: std_logic; attribute dont_touch of G4361: signal is true;
	signal G4362: std_logic; attribute dont_touch of G4362: signal is true;
	signal G4363: std_logic; attribute dont_touch of G4363: signal is true;
	signal G4364: std_logic; attribute dont_touch of G4364: signal is true;
	signal G4365: std_logic; attribute dont_touch of G4365: signal is true;
	signal G4366: std_logic; attribute dont_touch of G4366: signal is true;
	signal G4367: std_logic; attribute dont_touch of G4367: signal is true;
	signal G4368: std_logic; attribute dont_touch of G4368: signal is true;
	signal G4369: std_logic; attribute dont_touch of G4369: signal is true;
	signal G4370: std_logic; attribute dont_touch of G4370: signal is true;
	signal G4371: std_logic; attribute dont_touch of G4371: signal is true;
	signal G4372: std_logic; attribute dont_touch of G4372: signal is true;
	signal G4373: std_logic; attribute dont_touch of G4373: signal is true;
	signal G4374: std_logic; attribute dont_touch of G4374: signal is true;
	signal G4375: std_logic; attribute dont_touch of G4375: signal is true;
	signal G4376: std_logic; attribute dont_touch of G4376: signal is true;
	signal G4377: std_logic; attribute dont_touch of G4377: signal is true;
	signal G4378: std_logic; attribute dont_touch of G4378: signal is true;
	signal G4379: std_logic; attribute dont_touch of G4379: signal is true;
	signal G4380: std_logic; attribute dont_touch of G4380: signal is true;
	signal G4381: std_logic; attribute dont_touch of G4381: signal is true;
	signal G4382: std_logic; attribute dont_touch of G4382: signal is true;
	signal G4383: std_logic; attribute dont_touch of G4383: signal is true;
	signal G4384: std_logic; attribute dont_touch of G4384: signal is true;
	signal G4385: std_logic; attribute dont_touch of G4385: signal is true;
	signal G4386: std_logic; attribute dont_touch of G4386: signal is true;
	signal G4387: std_logic; attribute dont_touch of G4387: signal is true;
	signal G4388: std_logic; attribute dont_touch of G4388: signal is true;
	signal G4389: std_logic; attribute dont_touch of G4389: signal is true;
	signal G4390: std_logic; attribute dont_touch of G4390: signal is true;
	signal G4391: std_logic; attribute dont_touch of G4391: signal is true;
	signal G4392: std_logic; attribute dont_touch of G4392: signal is true;
	signal G4393: std_logic; attribute dont_touch of G4393: signal is true;
	signal G4394: std_logic; attribute dont_touch of G4394: signal is true;
	signal G4395: std_logic; attribute dont_touch of G4395: signal is true;
	signal G4396: std_logic; attribute dont_touch of G4396: signal is true;
	signal G4397: std_logic; attribute dont_touch of G4397: signal is true;
	signal G4398: std_logic; attribute dont_touch of G4398: signal is true;
	signal G4399: std_logic; attribute dont_touch of G4399: signal is true;
	signal G4400: std_logic; attribute dont_touch of G4400: signal is true;
	signal G4401: std_logic; attribute dont_touch of G4401: signal is true;
	signal G4411: std_logic; attribute dont_touch of G4411: signal is true;
	signal G4412: std_logic; attribute dont_touch of G4412: signal is true;
	signal G4413: std_logic; attribute dont_touch of G4413: signal is true;
	signal G4414: std_logic; attribute dont_touch of G4414: signal is true;
	signal G4415: std_logic; attribute dont_touch of G4415: signal is true;
	signal G4416: std_logic; attribute dont_touch of G4416: signal is true;
	signal G4417: std_logic; attribute dont_touch of G4417: signal is true;
	signal G4418: std_logic; attribute dont_touch of G4418: signal is true;
	signal G4419: std_logic; attribute dont_touch of G4419: signal is true;
	signal G4420: std_logic; attribute dont_touch of G4420: signal is true;
	signal G4421: std_logic; attribute dont_touch of G4421: signal is true;
	signal G4424: std_logic; attribute dont_touch of G4424: signal is true;
	signal G4425: std_logic; attribute dont_touch of G4425: signal is true;
	signal G4426: std_logic; attribute dont_touch of G4426: signal is true;
	signal G4427: std_logic; attribute dont_touch of G4427: signal is true;
	signal G4428: std_logic; attribute dont_touch of G4428: signal is true;
	signal G4429: std_logic; attribute dont_touch of G4429: signal is true;
	signal G4430: std_logic; attribute dont_touch of G4430: signal is true;
	signal G4431: std_logic; attribute dont_touch of G4431: signal is true;
	signal G4432: std_logic; attribute dont_touch of G4432: signal is true;
	signal G4435: std_logic; attribute dont_touch of G4435: signal is true;
	signal G4436: std_logic; attribute dont_touch of G4436: signal is true;
	signal G4437: std_logic; attribute dont_touch of G4437: signal is true;
	signal G4438: std_logic; attribute dont_touch of G4438: signal is true;
	signal G4439: std_logic; attribute dont_touch of G4439: signal is true;
	signal G4440: std_logic; attribute dont_touch of G4440: signal is true;
	signal G4441: std_logic; attribute dont_touch of G4441: signal is true;
	signal G4442: std_logic; attribute dont_touch of G4442: signal is true;
	signal G4443: std_logic; attribute dont_touch of G4443: signal is true;
	signal G4444: std_logic; attribute dont_touch of G4444: signal is true;
	signal G4445: std_logic; attribute dont_touch of G4445: signal is true;
	signal G4449: std_logic; attribute dont_touch of G4449: signal is true;
	signal G4450: std_logic; attribute dont_touch of G4450: signal is true;
	signal G4451: std_logic; attribute dont_touch of G4451: signal is true;
	signal G4452: std_logic; attribute dont_touch of G4452: signal is true;
	signal G4453: std_logic; attribute dont_touch of G4453: signal is true;
	signal G4454: std_logic; attribute dont_touch of G4454: signal is true;
	signal G4455: std_logic; attribute dont_touch of G4455: signal is true;
	signal G4456: std_logic; attribute dont_touch of G4456: signal is true;
	signal G4457: std_logic; attribute dont_touch of G4457: signal is true;
	signal G4458: std_logic; attribute dont_touch of G4458: signal is true;
	signal G4459: std_logic; attribute dont_touch of G4459: signal is true;
	signal G4460: std_logic; attribute dont_touch of G4460: signal is true;
	signal G4461: std_logic; attribute dont_touch of G4461: signal is true;
	signal G4462: std_logic; attribute dont_touch of G4462: signal is true;
	signal G4463: std_logic; attribute dont_touch of G4463: signal is true;
	signal G4464: std_logic; attribute dont_touch of G4464: signal is true;
	signal G4465: std_logic; attribute dont_touch of G4465: signal is true;
	signal G4466: std_logic; attribute dont_touch of G4466: signal is true;
	signal G4467: std_logic; attribute dont_touch of G4467: signal is true;
	signal G4468: std_logic; attribute dont_touch of G4468: signal is true;
	signal G4469: std_logic; attribute dont_touch of G4469: signal is true;
	signal G4470: std_logic; attribute dont_touch of G4470: signal is true;
	signal G4471: std_logic; attribute dont_touch of G4471: signal is true;
	signal G4472: std_logic; attribute dont_touch of G4472: signal is true;
	signal G4473: std_logic; attribute dont_touch of G4473: signal is true;
	signal G4474: std_logic; attribute dont_touch of G4474: signal is true;
	signal G4475: std_logic; attribute dont_touch of G4475: signal is true;
	signal G4476: std_logic; attribute dont_touch of G4476: signal is true;
	signal G4477: std_logic; attribute dont_touch of G4477: signal is true;
	signal G4478: std_logic; attribute dont_touch of G4478: signal is true;
	signal G4479: std_logic; attribute dont_touch of G4479: signal is true;
	signal G4480: std_logic; attribute dont_touch of G4480: signal is true;
	signal G4481: std_logic; attribute dont_touch of G4481: signal is true;
	signal G4482: std_logic; attribute dont_touch of G4482: signal is true;
	signal G4483: std_logic; attribute dont_touch of G4483: signal is true;
	signal G4484: std_logic; attribute dont_touch of G4484: signal is true;
	signal G4485: std_logic; attribute dont_touch of G4485: signal is true;
	signal G4486: std_logic; attribute dont_touch of G4486: signal is true;
	signal G4487: std_logic; attribute dont_touch of G4487: signal is true;
	signal G4488: std_logic; attribute dont_touch of G4488: signal is true;
	signal G4489: std_logic; attribute dont_touch of G4489: signal is true;
	signal G4490: std_logic; attribute dont_touch of G4490: signal is true;
	signal G4491: std_logic; attribute dont_touch of G4491: signal is true;
	signal G4492: std_logic; attribute dont_touch of G4492: signal is true;
	signal G4495: std_logic; attribute dont_touch of G4495: signal is true;
	signal G4496: std_logic; attribute dont_touch of G4496: signal is true;
	signal G4497: std_logic; attribute dont_touch of G4497: signal is true;
	signal G4498: std_logic; attribute dont_touch of G4498: signal is true;
	signal G4499: std_logic; attribute dont_touch of G4499: signal is true;
	signal G4500: std_logic; attribute dont_touch of G4500: signal is true;
	signal G4501: std_logic; attribute dont_touch of G4501: signal is true;
	signal G4502: std_logic; attribute dont_touch of G4502: signal is true;
	signal G4503: std_logic; attribute dont_touch of G4503: signal is true;
	signal G4504: std_logic; attribute dont_touch of G4504: signal is true;
	signal G4505: std_logic; attribute dont_touch of G4505: signal is true;
	signal G4506: std_logic; attribute dont_touch of G4506: signal is true;
	signal G4507: std_logic; attribute dont_touch of G4507: signal is true;
	signal G4508: std_logic; attribute dont_touch of G4508: signal is true;
	signal G4509: std_logic; attribute dont_touch of G4509: signal is true;
	signal G4510: std_logic; attribute dont_touch of G4510: signal is true;
	signal G4511: std_logic; attribute dont_touch of G4511: signal is true;
	signal G4512: std_logic; attribute dont_touch of G4512: signal is true;
	signal G4513: std_logic; attribute dont_touch of G4513: signal is true;
	signal G4514: std_logic; attribute dont_touch of G4514: signal is true;
	signal G4515: std_logic; attribute dont_touch of G4515: signal is true;
	signal G4518: std_logic; attribute dont_touch of G4518: signal is true;
	signal G4519: std_logic; attribute dont_touch of G4519: signal is true;
	signal G4520: std_logic; attribute dont_touch of G4520: signal is true;
	signal G4521: std_logic; attribute dont_touch of G4521: signal is true;
	signal G4522: std_logic; attribute dont_touch of G4522: signal is true;
	signal G4523: std_logic; attribute dont_touch of G4523: signal is true;
	signal G4524: std_logic; attribute dont_touch of G4524: signal is true;
	signal G4525: std_logic; attribute dont_touch of G4525: signal is true;
	signal G4526: std_logic; attribute dont_touch of G4526: signal is true;
	signal G4529: std_logic; attribute dont_touch of G4529: signal is true;
	signal G4530: std_logic; attribute dont_touch of G4530: signal is true;
	signal G4533: std_logic; attribute dont_touch of G4533: signal is true;
	signal G4534: std_logic; attribute dont_touch of G4534: signal is true;
	signal G4535: std_logic; attribute dont_touch of G4535: signal is true;
	signal G4536: std_logic; attribute dont_touch of G4536: signal is true;
	signal G4537: std_logic; attribute dont_touch of G4537: signal is true;
	signal G4538: std_logic; attribute dont_touch of G4538: signal is true;
	signal G4541: std_logic; attribute dont_touch of G4541: signal is true;
	signal G4542: std_logic; attribute dont_touch of G4542: signal is true;
	signal G4543: std_logic; attribute dont_touch of G4543: signal is true;
	signal G4544: std_logic; attribute dont_touch of G4544: signal is true;
	signal G4545: std_logic; attribute dont_touch of G4545: signal is true;
	signal G4548: std_logic; attribute dont_touch of G4548: signal is true;
	signal G4549: std_logic; attribute dont_touch of G4549: signal is true;
	signal G4550: std_logic; attribute dont_touch of G4550: signal is true;
	signal G4551: std_logic; attribute dont_touch of G4551: signal is true;
	signal G4552: std_logic; attribute dont_touch of G4552: signal is true;
	signal G4553: std_logic; attribute dont_touch of G4553: signal is true;
	signal G4554: std_logic; attribute dont_touch of G4554: signal is true;
	signal G4555: std_logic; attribute dont_touch of G4555: signal is true;
	signal G4556: std_logic; attribute dont_touch of G4556: signal is true;
	signal G4557: std_logic; attribute dont_touch of G4557: signal is true;
	signal G4558: std_logic; attribute dont_touch of G4558: signal is true;
	signal G4559: std_logic; attribute dont_touch of G4559: signal is true;
	signal G4560: std_logic; attribute dont_touch of G4560: signal is true;
	signal G4561: std_logic; attribute dont_touch of G4561: signal is true;
	signal G4562: std_logic; attribute dont_touch of G4562: signal is true;
	signal G4563: std_logic; attribute dont_touch of G4563: signal is true;
	signal G4564: std_logic; attribute dont_touch of G4564: signal is true;
	signal G4565: std_logic; attribute dont_touch of G4565: signal is true;
	signal G4566: std_logic; attribute dont_touch of G4566: signal is true;
	signal G4567: std_logic; attribute dont_touch of G4567: signal is true;
	signal G4572: std_logic; attribute dont_touch of G4572: signal is true;
	signal G4575: std_logic; attribute dont_touch of G4575: signal is true;
	signal G4576: std_logic; attribute dont_touch of G4576: signal is true;
	signal G4577: std_logic; attribute dont_touch of G4577: signal is true;
	signal G4580: std_logic; attribute dont_touch of G4580: signal is true;
	signal G4581: std_logic; attribute dont_touch of G4581: signal is true;
	signal G4582: std_logic; attribute dont_touch of G4582: signal is true;
	signal G4583: std_logic; attribute dont_touch of G4583: signal is true;
	signal G4584: std_logic; attribute dont_touch of G4584: signal is true;
	signal G4585: std_logic; attribute dont_touch of G4585: signal is true;
	signal G4586: std_logic; attribute dont_touch of G4586: signal is true;
	signal G4587: std_logic; attribute dont_touch of G4587: signal is true;
	signal G4588: std_logic; attribute dont_touch of G4588: signal is true;
	signal G4589: std_logic; attribute dont_touch of G4589: signal is true;
	signal G4590: std_logic; attribute dont_touch of G4590: signal is true;
	signal G4591: std_logic; attribute dont_touch of G4591: signal is true;
	signal G4592: std_logic; attribute dont_touch of G4592: signal is true;
	signal G4593: std_logic; attribute dont_touch of G4593: signal is true;
	signal G4596: std_logic; attribute dont_touch of G4596: signal is true;
	signal G4601: std_logic; attribute dont_touch of G4601: signal is true;
	signal G4602: std_logic; attribute dont_touch of G4602: signal is true;
	signal G4603: std_logic; attribute dont_touch of G4603: signal is true;
	signal G4604: std_logic; attribute dont_touch of G4604: signal is true;
	signal G4605: std_logic; attribute dont_touch of G4605: signal is true;
	signal G4606: std_logic; attribute dont_touch of G4606: signal is true;
	signal G4607: std_logic; attribute dont_touch of G4607: signal is true;
	signal G4608: std_logic; attribute dont_touch of G4608: signal is true;
	signal G4609: std_logic; attribute dont_touch of G4609: signal is true;
	signal G4610: std_logic; attribute dont_touch of G4610: signal is true;
	signal G4613: std_logic; attribute dont_touch of G4613: signal is true;
	signal G4614: std_logic; attribute dont_touch of G4614: signal is true;
	signal G4615: std_logic; attribute dont_touch of G4615: signal is true;
	signal G4616: std_logic; attribute dont_touch of G4616: signal is true;
	signal G4617: std_logic; attribute dont_touch of G4617: signal is true;
	signal G4618: std_logic; attribute dont_touch of G4618: signal is true;
	signal G4619: std_logic; attribute dont_touch of G4619: signal is true;
	signal G4620: std_logic; attribute dont_touch of G4620: signal is true;
	signal G4630: std_logic; attribute dont_touch of G4630: signal is true;
	signal G4631: std_logic; attribute dont_touch of G4631: signal is true;
	signal G4636: std_logic; attribute dont_touch of G4636: signal is true;
	signal G4637: std_logic; attribute dont_touch of G4637: signal is true;
	signal G4638: std_logic; attribute dont_touch of G4638: signal is true;
	signal G4639: std_logic; attribute dont_touch of G4639: signal is true;
	signal G4640: std_logic; attribute dont_touch of G4640: signal is true;
	signal G4669: std_logic; attribute dont_touch of G4669: signal is true;
	signal G4670: std_logic; attribute dont_touch of G4670: signal is true;
	signal G4671: std_logic; attribute dont_touch of G4671: signal is true;
	signal G4672: std_logic; attribute dont_touch of G4672: signal is true;
	signal G4673: std_logic; attribute dont_touch of G4673: signal is true;
	signal G4674: std_logic; attribute dont_touch of G4674: signal is true;
	signal G4675: std_logic; attribute dont_touch of G4675: signal is true;
	signal G4676: std_logic; attribute dont_touch of G4676: signal is true;
	signal G4677: std_logic; attribute dont_touch of G4677: signal is true;
	signal G4678: std_logic; attribute dont_touch of G4678: signal is true;
	signal G4679: std_logic; attribute dont_touch of G4679: signal is true;
	signal G4680: std_logic; attribute dont_touch of G4680: signal is true;
	signal G4681: std_logic; attribute dont_touch of G4681: signal is true;
	signal G4682: std_logic; attribute dont_touch of G4682: signal is true;
	signal G4711: std_logic; attribute dont_touch of G4711: signal is true;
	signal G4712: std_logic; attribute dont_touch of G4712: signal is true;
	signal G4713: std_logic; attribute dont_touch of G4713: signal is true;
	signal G4714: std_logic; attribute dont_touch of G4714: signal is true;
	signal G4715: std_logic; attribute dont_touch of G4715: signal is true;
	signal G4716: std_logic; attribute dont_touch of G4716: signal is true;
	signal G4717: std_logic; attribute dont_touch of G4717: signal is true;
	signal G4718: std_logic; attribute dont_touch of G4718: signal is true;
	signal G4719: std_logic; attribute dont_touch of G4719: signal is true;
	signal G4720: std_logic; attribute dont_touch of G4720: signal is true;
	signal G4721: std_logic; attribute dont_touch of G4721: signal is true;
	signal G4722: std_logic; attribute dont_touch of G4722: signal is true;
	signal G4723: std_logic; attribute dont_touch of G4723: signal is true;
	signal G4724: std_logic; attribute dont_touch of G4724: signal is true;
	signal G4725: std_logic; attribute dont_touch of G4725: signal is true;
	signal G4726: std_logic; attribute dont_touch of G4726: signal is true;
	signal G4727: std_logic; attribute dont_touch of G4727: signal is true;
	signal G4728: std_logic; attribute dont_touch of G4728: signal is true;
	signal G4729: std_logic; attribute dont_touch of G4729: signal is true;
	signal G4730: std_logic; attribute dont_touch of G4730: signal is true;
	signal G4731: std_logic; attribute dont_touch of G4731: signal is true;
	signal G4732: std_logic; attribute dont_touch of G4732: signal is true;
	signal G4733: std_logic; attribute dont_touch of G4733: signal is true;
	signal G4734: std_logic; attribute dont_touch of G4734: signal is true;
	signal G4735: std_logic; attribute dont_touch of G4735: signal is true;
	signal G4736: std_logic; attribute dont_touch of G4736: signal is true;
	signal G4737: std_logic; attribute dont_touch of G4737: signal is true;
	signal G4738: std_logic; attribute dont_touch of G4738: signal is true;
	signal G4739: std_logic; attribute dont_touch of G4739: signal is true;
	signal G4746: std_logic; attribute dont_touch of G4746: signal is true;
	signal G4747: std_logic; attribute dont_touch of G4747: signal is true;
	signal G4748: std_logic; attribute dont_touch of G4748: signal is true;
	signal G4749: std_logic; attribute dont_touch of G4749: signal is true;
	signal G4752: std_logic; attribute dont_touch of G4752: signal is true;
	signal G4753: std_logic; attribute dont_touch of G4753: signal is true;
	signal G4754: std_logic; attribute dont_touch of G4754: signal is true;
	signal G4755: std_logic; attribute dont_touch of G4755: signal is true;
	signal G4756: std_logic; attribute dont_touch of G4756: signal is true;
	signal G4757: std_logic; attribute dont_touch of G4757: signal is true;
	signal G4758: std_logic; attribute dont_touch of G4758: signal is true;
	signal G4759: std_logic; attribute dont_touch of G4759: signal is true;
	signal G4760: std_logic; attribute dont_touch of G4760: signal is true;
	signal G4761: std_logic; attribute dont_touch of G4761: signal is true;
	signal G4762: std_logic; attribute dont_touch of G4762: signal is true;
	signal G4763: std_logic; attribute dont_touch of G4763: signal is true;
	signal G4764: std_logic; attribute dont_touch of G4764: signal is true;
	signal G4765: std_logic; attribute dont_touch of G4765: signal is true;
	signal G4766: std_logic; attribute dont_touch of G4766: signal is true;
	signal G4767: std_logic; attribute dont_touch of G4767: signal is true;
	signal G4768: std_logic; attribute dont_touch of G4768: signal is true;
	signal G4769: std_logic; attribute dont_touch of G4769: signal is true;
	signal G4770: std_logic; attribute dont_touch of G4770: signal is true;
	signal G4771: std_logic; attribute dont_touch of G4771: signal is true;
	signal G4772: std_logic; attribute dont_touch of G4772: signal is true;
	signal G4773: std_logic; attribute dont_touch of G4773: signal is true;
	signal G4774: std_logic; attribute dont_touch of G4774: signal is true;
	signal G4775: std_logic; attribute dont_touch of G4775: signal is true;
	signal G4776: std_logic; attribute dont_touch of G4776: signal is true;
	signal G4777: std_logic; attribute dont_touch of G4777: signal is true;
	signal G4778: std_logic; attribute dont_touch of G4778: signal is true;
	signal G4779: std_logic; attribute dont_touch of G4779: signal is true;
	signal G4780: std_logic; attribute dont_touch of G4780: signal is true;
	signal G4781: std_logic; attribute dont_touch of G4781: signal is true;
	signal G4782: std_logic; attribute dont_touch of G4782: signal is true;
	signal G4783: std_logic; attribute dont_touch of G4783: signal is true;
	signal G4784: std_logic; attribute dont_touch of G4784: signal is true;
	signal G4785: std_logic; attribute dont_touch of G4785: signal is true;
	signal G4786: std_logic; attribute dont_touch of G4786: signal is true;
	signal G4787: std_logic; attribute dont_touch of G4787: signal is true;
	signal G4788: std_logic; attribute dont_touch of G4788: signal is true;
	signal G4789: std_logic; attribute dont_touch of G4789: signal is true;
	signal G4790: std_logic; attribute dont_touch of G4790: signal is true;
	signal G4791: std_logic; attribute dont_touch of G4791: signal is true;
	signal G4794: std_logic; attribute dont_touch of G4794: signal is true;
	signal G4801: std_logic; attribute dont_touch of G4801: signal is true;
	signal G4802: std_logic; attribute dont_touch of G4802: signal is true;
	signal G4803: std_logic; attribute dont_touch of G4803: signal is true;
	signal G4804: std_logic; attribute dont_touch of G4804: signal is true;
	signal G4805: std_logic; attribute dont_touch of G4805: signal is true;
	signal G4806: std_logic; attribute dont_touch of G4806: signal is true;
	signal G4807: std_logic; attribute dont_touch of G4807: signal is true;
	signal G4811: std_logic; attribute dont_touch of G4811: signal is true;
	signal G4816: std_logic; attribute dont_touch of G4816: signal is true;
	signal G4819: std_logic; attribute dont_touch of G4819: signal is true;
	signal G4820: std_logic; attribute dont_touch of G4820: signal is true;
	signal G4821: std_logic; attribute dont_touch of G4821: signal is true;
	signal G4822: std_logic; attribute dont_touch of G4822: signal is true;
	signal G4823: std_logic; attribute dont_touch of G4823: signal is true;
	signal G4824: std_logic; attribute dont_touch of G4824: signal is true;
	signal G4827: std_logic; attribute dont_touch of G4827: signal is true;
	signal G4828: std_logic; attribute dont_touch of G4828: signal is true;
	signal G4831: std_logic; attribute dont_touch of G4831: signal is true;
	signal G4834: std_logic; attribute dont_touch of G4834: signal is true;
	signal G4835: std_logic; attribute dont_touch of G4835: signal is true;
	signal G4836: std_logic; attribute dont_touch of G4836: signal is true;
	signal G4837: std_logic; attribute dont_touch of G4837: signal is true;
	signal G4838: std_logic; attribute dont_touch of G4838: signal is true;
	signal G4839: std_logic; attribute dont_touch of G4839: signal is true;
	signal G4840: std_logic; attribute dont_touch of G4840: signal is true;
	signal G4865: std_logic; attribute dont_touch of G4865: signal is true;
	signal G4866: std_logic; attribute dont_touch of G4866: signal is true;
	signal G4867: std_logic; attribute dont_touch of G4867: signal is true;
	signal G4868: std_logic; attribute dont_touch of G4868: signal is true;
	signal G4869: std_logic; attribute dont_touch of G4869: signal is true;
	signal G4870: std_logic; attribute dont_touch of G4870: signal is true;
	signal G4871: std_logic; attribute dont_touch of G4871: signal is true;
	signal G4872: std_logic; attribute dont_touch of G4872: signal is true;
	signal G4873: std_logic; attribute dont_touch of G4873: signal is true;
	signal G4874: std_logic; attribute dont_touch of G4874: signal is true;
	signal G4875: std_logic; attribute dont_touch of G4875: signal is true;
	signal G4876: std_logic; attribute dont_touch of G4876: signal is true;
	signal G4877: std_logic; attribute dont_touch of G4877: signal is true;
	signal G4878: std_logic; attribute dont_touch of G4878: signal is true;
	signal G4879: std_logic; attribute dont_touch of G4879: signal is true;
	signal G4880: std_logic; attribute dont_touch of G4880: signal is true;
	signal G4881: std_logic; attribute dont_touch of G4881: signal is true;
	signal G4882: std_logic; attribute dont_touch of G4882: signal is true;
	signal G4883: std_logic; attribute dont_touch of G4883: signal is true;
	signal G4884: std_logic; attribute dont_touch of G4884: signal is true;
	signal G4885: std_logic; attribute dont_touch of G4885: signal is true;
	signal G4886: std_logic; attribute dont_touch of G4886: signal is true;
	signal G4889: std_logic; attribute dont_touch of G4889: signal is true;
	signal G4890: std_logic; attribute dont_touch of G4890: signal is true;
	signal G4891: std_logic; attribute dont_touch of G4891: signal is true;
	signal G4892: std_logic; attribute dont_touch of G4892: signal is true;
	signal G4893: std_logic; attribute dont_touch of G4893: signal is true;
	signal G4894: std_logic; attribute dont_touch of G4894: signal is true;
	signal G4895: std_logic; attribute dont_touch of G4895: signal is true;
	signal G4896: std_logic; attribute dont_touch of G4896: signal is true;
	signal G4897: std_logic; attribute dont_touch of G4897: signal is true;
	signal G4898: std_logic; attribute dont_touch of G4898: signal is true;
	signal G4899: std_logic; attribute dont_touch of G4899: signal is true;
	signal G4900: std_logic; attribute dont_touch of G4900: signal is true;
	signal G4901: std_logic; attribute dont_touch of G4901: signal is true;
	signal G4902: std_logic; attribute dont_touch of G4902: signal is true;
	signal G4903: std_logic; attribute dont_touch of G4903: signal is true;
	signal G4904: std_logic; attribute dont_touch of G4904: signal is true;
	signal G4905: std_logic; attribute dont_touch of G4905: signal is true;
	signal G4906: std_logic; attribute dont_touch of G4906: signal is true;
	signal G4907: std_logic; attribute dont_touch of G4907: signal is true;
	signal G4908: std_logic; attribute dont_touch of G4908: signal is true;
	signal G4912: std_logic; attribute dont_touch of G4912: signal is true;
	signal G4913: std_logic; attribute dont_touch of G4913: signal is true;
	signal G4914: std_logic; attribute dont_touch of G4914: signal is true;
	signal G4915: std_logic; attribute dont_touch of G4915: signal is true;
	signal G4919: std_logic; attribute dont_touch of G4919: signal is true;
	signal G4920: std_logic; attribute dont_touch of G4920: signal is true;
	signal G4921: std_logic; attribute dont_touch of G4921: signal is true;
	signal G4932: std_logic; attribute dont_touch of G4932: signal is true;
	signal G4933: std_logic; attribute dont_touch of G4933: signal is true;
	signal G4934: std_logic; attribute dont_touch of G4934: signal is true;
	signal G4935: std_logic; attribute dont_touch of G4935: signal is true;
	signal G4939: std_logic; attribute dont_touch of G4939: signal is true;
	signal G4940: std_logic; attribute dont_touch of G4940: signal is true;
	signal G4941: std_logic; attribute dont_touch of G4941: signal is true;
	signal G4942: std_logic; attribute dont_touch of G4942: signal is true;
	signal G4943: std_logic; attribute dont_touch of G4943: signal is true;
	signal G4944: std_logic; attribute dont_touch of G4944: signal is true;
	signal G4948: std_logic; attribute dont_touch of G4948: signal is true;
	signal G4949: std_logic; attribute dont_touch of G4949: signal is true;
	signal G4950: std_logic; attribute dont_touch of G4950: signal is true;
	signal G4951: std_logic; attribute dont_touch of G4951: signal is true;
	signal G4952: std_logic; attribute dont_touch of G4952: signal is true;
	signal G4953: std_logic; attribute dont_touch of G4953: signal is true;
	signal G4954: std_logic; attribute dont_touch of G4954: signal is true;
	signal G4958: std_logic; attribute dont_touch of G4958: signal is true;
	signal G4959: std_logic; attribute dont_touch of G4959: signal is true;
	signal G4960: std_logic; attribute dont_touch of G4960: signal is true;
	signal G4961: std_logic; attribute dont_touch of G4961: signal is true;
	signal G4962: std_logic; attribute dont_touch of G4962: signal is true;
	signal G4963: std_logic; attribute dont_touch of G4963: signal is true;
	signal G4966: std_logic; attribute dont_touch of G4966: signal is true;
	signal G4967: std_logic; attribute dont_touch of G4967: signal is true;
	signal G4968: std_logic; attribute dont_touch of G4968: signal is true;
	signal G4969: std_logic; attribute dont_touch of G4969: signal is true;
	signal G4970: std_logic; attribute dont_touch of G4970: signal is true;
	signal G4971: std_logic; attribute dont_touch of G4971: signal is true;
	signal G4972: std_logic; attribute dont_touch of G4972: signal is true;
	signal G4973: std_logic; attribute dont_touch of G4973: signal is true;
	signal G4974: std_logic; attribute dont_touch of G4974: signal is true;
	signal G4975: std_logic; attribute dont_touch of G4975: signal is true;
	signal G4976: std_logic; attribute dont_touch of G4976: signal is true;
	signal G4977: std_logic; attribute dont_touch of G4977: signal is true;
	signal G4986: std_logic; attribute dont_touch of G4986: signal is true;
	signal G4987: std_logic; attribute dont_touch of G4987: signal is true;
	signal G4988: std_logic; attribute dont_touch of G4988: signal is true;
	signal G4989: std_logic; attribute dont_touch of G4989: signal is true;
	signal G4990: std_logic; attribute dont_touch of G4990: signal is true;
	signal G4991: std_logic; attribute dont_touch of G4991: signal is true;
	signal G4992: std_logic; attribute dont_touch of G4992: signal is true;
	signal G4993: std_logic; attribute dont_touch of G4993: signal is true;
	signal G4994: std_logic; attribute dont_touch of G4994: signal is true;
	signal G4995: std_logic; attribute dont_touch of G4995: signal is true;
	signal G4996: std_logic; attribute dont_touch of G4996: signal is true;
	signal G4997: std_logic; attribute dont_touch of G4997: signal is true;
	signal G4998: std_logic; attribute dont_touch of G4998: signal is true;
	signal G4999: std_logic; attribute dont_touch of G4999: signal is true;
	signal G5000: std_logic; attribute dont_touch of G5000: signal is true;
	signal G5001: std_logic; attribute dont_touch of G5001: signal is true;
	signal G5002: std_logic; attribute dont_touch of G5002: signal is true;
	signal G5003: std_logic; attribute dont_touch of G5003: signal is true;
	signal G5004: std_logic; attribute dont_touch of G5004: signal is true;
	signal G5005: std_logic; attribute dont_touch of G5005: signal is true;
	signal G5006: std_logic; attribute dont_touch of G5006: signal is true;
	signal G5007: std_logic; attribute dont_touch of G5007: signal is true;
	signal G5008: std_logic; attribute dont_touch of G5008: signal is true;
	signal G5009: std_logic; attribute dont_touch of G5009: signal is true;
	signal G5010: std_logic; attribute dont_touch of G5010: signal is true;
	signal G5011: std_logic; attribute dont_touch of G5011: signal is true;
	signal G5012: std_logic; attribute dont_touch of G5012: signal is true;
	signal G5013: std_logic; attribute dont_touch of G5013: signal is true;
	signal G5023: std_logic; attribute dont_touch of G5023: signal is true;
	signal G5024: std_logic; attribute dont_touch of G5024: signal is true;
	signal G5025: std_logic; attribute dont_touch of G5025: signal is true;
	signal G5026: std_logic; attribute dont_touch of G5026: signal is true;
	signal G5027: std_logic; attribute dont_touch of G5027: signal is true;
	signal G5028: std_logic; attribute dont_touch of G5028: signal is true;
	signal G5029: std_logic; attribute dont_touch of G5029: signal is true;
	signal G5030: std_logic; attribute dont_touch of G5030: signal is true;
	signal G5031: std_logic; attribute dont_touch of G5031: signal is true;
	signal G5032: std_logic; attribute dont_touch of G5032: signal is true;
	signal G5033: std_logic; attribute dont_touch of G5033: signal is true;
	signal G5034: std_logic; attribute dont_touch of G5034: signal is true;
	signal G5035: std_logic; attribute dont_touch of G5035: signal is true;
	signal G5036: std_logic; attribute dont_touch of G5036: signal is true;
	signal G5037: std_logic; attribute dont_touch of G5037: signal is true;
	signal G5038: std_logic; attribute dont_touch of G5038: signal is true;
	signal G5039: std_logic; attribute dont_touch of G5039: signal is true;
	signal G5040: std_logic; attribute dont_touch of G5040: signal is true;
	signal G5041: std_logic; attribute dont_touch of G5041: signal is true;
	signal G5042: std_logic; attribute dont_touch of G5042: signal is true;
	signal G5043: std_logic; attribute dont_touch of G5043: signal is true;
	signal G5044: std_logic; attribute dont_touch of G5044: signal is true;
	signal G5047: std_logic; attribute dont_touch of G5047: signal is true;
	signal G5050: std_logic; attribute dont_touch of G5050: signal is true;
	signal G5051: std_logic; attribute dont_touch of G5051: signal is true;
	signal G5052: std_logic; attribute dont_touch of G5052: signal is true;
	signal G5062: std_logic; attribute dont_touch of G5062: signal is true;
	signal G5063: std_logic; attribute dont_touch of G5063: signal is true;
	signal G5066: std_logic; attribute dont_touch of G5066: signal is true;
	signal G5067: std_logic; attribute dont_touch of G5067: signal is true;
	signal G5068: std_logic; attribute dont_touch of G5068: signal is true;
	signal G5069: std_logic; attribute dont_touch of G5069: signal is true;
	signal G5072: std_logic; attribute dont_touch of G5072: signal is true;
	signal G5073: std_logic; attribute dont_touch of G5073: signal is true;
	signal G5074: std_logic; attribute dont_touch of G5074: signal is true;
	signal G5075: std_logic; attribute dont_touch of G5075: signal is true;
	signal G5078: std_logic; attribute dont_touch of G5078: signal is true;
	signal G5081: std_logic; attribute dont_touch of G5081: signal is true;
	signal G5082: std_logic; attribute dont_touch of G5082: signal is true;
	signal G5083: std_logic; attribute dont_touch of G5083: signal is true;
	signal G5084: std_logic; attribute dont_touch of G5084: signal is true;
	signal G5085: std_logic; attribute dont_touch of G5085: signal is true;
	signal G5088: std_logic; attribute dont_touch of G5088: signal is true;
	signal G5089: std_logic; attribute dont_touch of G5089: signal is true;
	signal G5090: std_logic; attribute dont_touch of G5090: signal is true;
	signal G5091: std_logic; attribute dont_touch of G5091: signal is true;
	signal G5094: std_logic; attribute dont_touch of G5094: signal is true;
	signal G5095: std_logic; attribute dont_touch of G5095: signal is true;
	signal G5096: std_logic; attribute dont_touch of G5096: signal is true;
	signal G5097: std_logic; attribute dont_touch of G5097: signal is true;
	signal G5098: std_logic; attribute dont_touch of G5098: signal is true;
	signal G5099: std_logic; attribute dont_touch of G5099: signal is true;
	signal G5100: std_logic; attribute dont_touch of G5100: signal is true;
	signal G5102: std_logic; attribute dont_touch of G5102: signal is true;
	signal G5103: std_logic; attribute dont_touch of G5103: signal is true;
	signal G5104: std_logic; attribute dont_touch of G5104: signal is true;
	signal G5106: std_logic; attribute dont_touch of G5106: signal is true;
	signal G5107: std_logic; attribute dont_touch of G5107: signal is true;
	signal G5108: std_logic; attribute dont_touch of G5108: signal is true;
	signal G5109: std_logic; attribute dont_touch of G5109: signal is true;
	signal G5110: std_logic; attribute dont_touch of G5110: signal is true;
	signal G5111: std_logic; attribute dont_touch of G5111: signal is true;
	signal G5112: std_logic; attribute dont_touch of G5112: signal is true;
	signal G5113: std_logic; attribute dont_touch of G5113: signal is true;
	signal G5114: std_logic; attribute dont_touch of G5114: signal is true;
	signal G5115: std_logic; attribute dont_touch of G5115: signal is true;
	signal G5116: std_logic; attribute dont_touch of G5116: signal is true;
	signal G5117: std_logic; attribute dont_touch of G5117: signal is true;
	signal G5118: std_logic; attribute dont_touch of G5118: signal is true;
	signal G5119: std_logic; attribute dont_touch of G5119: signal is true;
	signal G5120: std_logic; attribute dont_touch of G5120: signal is true;
	signal G5121: std_logic; attribute dont_touch of G5121: signal is true;
	signal G5122: std_logic; attribute dont_touch of G5122: signal is true;
	signal G5123: std_logic; attribute dont_touch of G5123: signal is true;
	signal G5124: std_logic; attribute dont_touch of G5124: signal is true;
	signal G5125: std_logic; attribute dont_touch of G5125: signal is true;
	signal G5126: std_logic; attribute dont_touch of G5126: signal is true;
	signal G5127: std_logic; attribute dont_touch of G5127: signal is true;
	signal G5128: std_logic; attribute dont_touch of G5128: signal is true;
	signal G5143: std_logic; attribute dont_touch of G5143: signal is true;
	signal G5144: std_logic; attribute dont_touch of G5144: signal is true;
	signal G5145: std_logic; attribute dont_touch of G5145: signal is true;
	signal G5146: std_logic; attribute dont_touch of G5146: signal is true;
	signal G5147: std_logic; attribute dont_touch of G5147: signal is true;
	signal G5148: std_logic; attribute dont_touch of G5148: signal is true;
	signal G5149: std_logic; attribute dont_touch of G5149: signal is true;
	signal G5150: std_logic; attribute dont_touch of G5150: signal is true;
	signal G5151: std_logic; attribute dont_touch of G5151: signal is true;
	signal G5166: std_logic; attribute dont_touch of G5166: signal is true;
	signal G5167: std_logic; attribute dont_touch of G5167: signal is true;
	signal G5168: std_logic; attribute dont_touch of G5168: signal is true;
	signal G5169: std_logic; attribute dont_touch of G5169: signal is true;
	signal G5170: std_logic; attribute dont_touch of G5170: signal is true;
	signal G5171: std_logic; attribute dont_touch of G5171: signal is true;
	signal G5172: std_logic; attribute dont_touch of G5172: signal is true;
	signal G5173: std_logic; attribute dont_touch of G5173: signal is true;
	signal G5174: std_logic; attribute dont_touch of G5174: signal is true;
	signal G5175: std_logic; attribute dont_touch of G5175: signal is true;
	signal G5176: std_logic; attribute dont_touch of G5176: signal is true;
	signal G5177: std_logic; attribute dont_touch of G5177: signal is true;
	signal G5178: std_logic; attribute dont_touch of G5178: signal is true;
	signal G5179: std_logic; attribute dont_touch of G5179: signal is true;
	signal G5180: std_logic; attribute dont_touch of G5180: signal is true;
	signal G5181: std_logic; attribute dont_touch of G5181: signal is true;
	signal G5182: std_logic; attribute dont_touch of G5182: signal is true;
	signal G5183: std_logic; attribute dont_touch of G5183: signal is true;
	signal G5184: std_logic; attribute dont_touch of G5184: signal is true;
	signal G5185: std_logic; attribute dont_touch of G5185: signal is true;
	signal G5186: std_logic; attribute dont_touch of G5186: signal is true;
	signal G5187: std_logic; attribute dont_touch of G5187: signal is true;
	signal G5188: std_logic; attribute dont_touch of G5188: signal is true;
	signal G5189: std_logic; attribute dont_touch of G5189: signal is true;
	signal G5190: std_logic; attribute dont_touch of G5190: signal is true;
	signal G5191: std_logic; attribute dont_touch of G5191: signal is true;
	signal G5192: std_logic; attribute dont_touch of G5192: signal is true;
	signal G5193: std_logic; attribute dont_touch of G5193: signal is true;
	signal G5194: std_logic; attribute dont_touch of G5194: signal is true;
	signal G5195: std_logic; attribute dont_touch of G5195: signal is true;
	signal G5196: std_logic; attribute dont_touch of G5196: signal is true;
	signal G5197: std_logic; attribute dont_touch of G5197: signal is true;
	signal G5198: std_logic; attribute dont_touch of G5198: signal is true;
	signal G5199: std_logic; attribute dont_touch of G5199: signal is true;
	signal G5200: std_logic; attribute dont_touch of G5200: signal is true;
	signal G5201: std_logic; attribute dont_touch of G5201: signal is true;
	signal G5202: std_logic; attribute dont_touch of G5202: signal is true;
	signal G5203: std_logic; attribute dont_touch of G5203: signal is true;
	signal G5204: std_logic; attribute dont_touch of G5204: signal is true;
	signal G5205: std_logic; attribute dont_touch of G5205: signal is true;
	signal G5209: std_logic; attribute dont_touch of G5209: signal is true;
	signal G5210: std_logic; attribute dont_touch of G5210: signal is true;
	signal G5211: std_logic; attribute dont_touch of G5211: signal is true;
	signal G5212: std_logic; attribute dont_touch of G5212: signal is true;
	signal G5213: std_logic; attribute dont_touch of G5213: signal is true;
	signal G5214: std_logic; attribute dont_touch of G5214: signal is true;
	signal G5215: std_logic; attribute dont_touch of G5215: signal is true;
	signal G5216: std_logic; attribute dont_touch of G5216: signal is true;
	signal G5217: std_logic; attribute dont_touch of G5217: signal is true;
	signal G5218: std_logic; attribute dont_touch of G5218: signal is true;
	signal G5219: std_logic; attribute dont_touch of G5219: signal is true;
	signal G5220: std_logic; attribute dont_touch of G5220: signal is true;
	signal G5221: std_logic; attribute dont_touch of G5221: signal is true;
	signal G5222: std_logic; attribute dont_touch of G5222: signal is true;
	signal G5223: std_logic; attribute dont_touch of G5223: signal is true;
	signal G5224: std_logic; attribute dont_touch of G5224: signal is true;
	signal G5225: std_logic; attribute dont_touch of G5225: signal is true;
	signal G5226: std_logic; attribute dont_touch of G5226: signal is true;
	signal G5227: std_logic; attribute dont_touch of G5227: signal is true;
	signal G5228: std_logic; attribute dont_touch of G5228: signal is true;
	signal G5229: std_logic; attribute dont_touch of G5229: signal is true;
	signal G5230: std_logic; attribute dont_touch of G5230: signal is true;
	signal G5231: std_logic; attribute dont_touch of G5231: signal is true;
	signal G5232: std_logic; attribute dont_touch of G5232: signal is true;
	signal G5233: std_logic; attribute dont_touch of G5233: signal is true;
	signal G5236: std_logic; attribute dont_touch of G5236: signal is true;
	signal G5241: std_logic; attribute dont_touch of G5241: signal is true;
	signal G5245: std_logic; attribute dont_touch of G5245: signal is true;
	signal G5248: std_logic; attribute dont_touch of G5248: signal is true;
	signal G5249: std_logic; attribute dont_touch of G5249: signal is true;
	signal G5250: std_logic; attribute dont_touch of G5250: signal is true;
	signal G5251: std_logic; attribute dont_touch of G5251: signal is true;
	signal G5252: std_logic; attribute dont_touch of G5252: signal is true;
	signal G5253: std_logic; attribute dont_touch of G5253: signal is true;
	signal G5254: std_logic; attribute dont_touch of G5254: signal is true;
	signal G5255: std_logic; attribute dont_touch of G5255: signal is true;
	signal G5256: std_logic; attribute dont_touch of G5256: signal is true;
	signal G5257: std_logic; attribute dont_touch of G5257: signal is true;
	signal G5258: std_logic; attribute dont_touch of G5258: signal is true;
	signal G5259: std_logic; attribute dont_touch of G5259: signal is true;
	signal G5260: std_logic; attribute dont_touch of G5260: signal is true;
	signal G5261: std_logic; attribute dont_touch of G5261: signal is true;
	signal G5262: std_logic; attribute dont_touch of G5262: signal is true;
	signal G5263: std_logic; attribute dont_touch of G5263: signal is true;
	signal G5264: std_logic; attribute dont_touch of G5264: signal is true;
	signal G5265: std_logic; attribute dont_touch of G5265: signal is true;
	signal G5266: std_logic; attribute dont_touch of G5266: signal is true;
	signal G5267: std_logic; attribute dont_touch of G5267: signal is true;
	signal G5268: std_logic; attribute dont_touch of G5268: signal is true;
	signal G5269: std_logic; attribute dont_touch of G5269: signal is true;
	signal G5270: std_logic; attribute dont_touch of G5270: signal is true;
	signal G5271: std_logic; attribute dont_touch of G5271: signal is true;
	signal G5272: std_logic; attribute dont_touch of G5272: signal is true;
	signal G5273: std_logic; attribute dont_touch of G5273: signal is true;
	signal G5274: std_logic; attribute dont_touch of G5274: signal is true;
	signal G5275: std_logic; attribute dont_touch of G5275: signal is true;
	signal G5276: std_logic; attribute dont_touch of G5276: signal is true;
	signal G5277: std_logic; attribute dont_touch of G5277: signal is true;
	signal G5278: std_logic; attribute dont_touch of G5278: signal is true;
	signal G5279: std_logic; attribute dont_touch of G5279: signal is true;
	signal G5280: std_logic; attribute dont_touch of G5280: signal is true;
	signal G5281: std_logic; attribute dont_touch of G5281: signal is true;
	signal G5284: std_logic; attribute dont_touch of G5284: signal is true;
	signal G5285: std_logic; attribute dont_touch of G5285: signal is true;
	signal G5286: std_logic; attribute dont_touch of G5286: signal is true;
	signal G5287: std_logic; attribute dont_touch of G5287: signal is true;
	signal G5288: std_logic; attribute dont_touch of G5288: signal is true;
	signal G5291: std_logic; attribute dont_touch of G5291: signal is true;
	signal G5292: std_logic; attribute dont_touch of G5292: signal is true;
	signal G5295: std_logic; attribute dont_touch of G5295: signal is true;
	signal G5296: std_logic; attribute dont_touch of G5296: signal is true;
	signal G5299: std_logic; attribute dont_touch of G5299: signal is true;
	signal G5300: std_logic; attribute dont_touch of G5300: signal is true;
	signal G5301: std_logic; attribute dont_touch of G5301: signal is true;
	signal G5304: std_logic; attribute dont_touch of G5304: signal is true;
	signal G5305: std_logic; attribute dont_touch of G5305: signal is true;
	signal G5308: std_logic; attribute dont_touch of G5308: signal is true;
	signal G5309: std_logic; attribute dont_touch of G5309: signal is true;
	signal G5314: std_logic; attribute dont_touch of G5314: signal is true;
	signal G5317: std_logic; attribute dont_touch of G5317: signal is true;
	signal G5318: std_logic; attribute dont_touch of G5318: signal is true;
	signal G5319: std_logic; attribute dont_touch of G5319: signal is true;
	signal G5320: std_logic; attribute dont_touch of G5320: signal is true;
	signal G5344: std_logic; attribute dont_touch of G5344: signal is true;
	signal G5345: std_logic; attribute dont_touch of G5345: signal is true;
	signal G5348: std_logic; attribute dont_touch of G5348: signal is true;
	signal G5349: std_logic; attribute dont_touch of G5349: signal is true;
	signal G5350: std_logic; attribute dont_touch of G5350: signal is true;
	signal G5353: std_logic; attribute dont_touch of G5353: signal is true;
	signal G5354: std_logic; attribute dont_touch of G5354: signal is true;
	signal G5360: std_logic; attribute dont_touch of G5360: signal is true;
	signal G5361: std_logic; attribute dont_touch of G5361: signal is true;
	signal G5390: std_logic; attribute dont_touch of G5390: signal is true;
	signal G5391: std_logic; attribute dont_touch of G5391: signal is true;
	signal G5392: std_logic; attribute dont_touch of G5392: signal is true;
	signal G5395: std_logic; attribute dont_touch of G5395: signal is true;
	signal G5396: std_logic; attribute dont_touch of G5396: signal is true;
	signal G5397: std_logic; attribute dont_touch of G5397: signal is true;
	signal G5398: std_logic; attribute dont_touch of G5398: signal is true;
	signal G5401: std_logic; attribute dont_touch of G5401: signal is true;
	signal G5402: std_logic; attribute dont_touch of G5402: signal is true;
	signal G5403: std_logic; attribute dont_touch of G5403: signal is true;
	signal G5404: std_logic; attribute dont_touch of G5404: signal is true;
	signal G5405: std_logic; attribute dont_touch of G5405: signal is true;
	signal G5415: std_logic; attribute dont_touch of G5415: signal is true;
	signal G5416: std_logic; attribute dont_touch of G5416: signal is true;
	signal G5417: std_logic; attribute dont_touch of G5417: signal is true;
	signal G5418: std_logic; attribute dont_touch of G5418: signal is true;
	signal G5419: std_logic; attribute dont_touch of G5419: signal is true;
	signal G5420: std_logic; attribute dont_touch of G5420: signal is true;
	signal G5421: std_logic; attribute dont_touch of G5421: signal is true;
	signal G5422: std_logic; attribute dont_touch of G5422: signal is true;
	signal G5423: std_logic; attribute dont_touch of G5423: signal is true;
	signal G5424: std_logic; attribute dont_touch of G5424: signal is true;
	signal G5425: std_logic; attribute dont_touch of G5425: signal is true;
	signal G5426: std_logic; attribute dont_touch of G5426: signal is true;
	signal G5443: std_logic; attribute dont_touch of G5443: signal is true;
	signal G5444: std_logic; attribute dont_touch of G5444: signal is true;
	signal G5445: std_logic; attribute dont_touch of G5445: signal is true;
	signal G5446: std_logic; attribute dont_touch of G5446: signal is true;
	signal G5469: std_logic; attribute dont_touch of G5469: signal is true;
	signal G5470: std_logic; attribute dont_touch of G5470: signal is true;
	signal G5471: std_logic; attribute dont_touch of G5471: signal is true;
	signal G5472: std_logic; attribute dont_touch of G5472: signal is true;
	signal G5473: std_logic; attribute dont_touch of G5473: signal is true;
	signal G5474: std_logic; attribute dont_touch of G5474: signal is true;
	signal G5475: std_logic; attribute dont_touch of G5475: signal is true;
	signal G5476: std_logic; attribute dont_touch of G5476: signal is true;
	signal G5477: std_logic; attribute dont_touch of G5477: signal is true;
	signal G5478: std_logic; attribute dont_touch of G5478: signal is true;
	signal G5479: std_logic; attribute dont_touch of G5479: signal is true;
	signal G5480: std_logic; attribute dont_touch of G5480: signal is true;
	signal G5481: std_logic; attribute dont_touch of G5481: signal is true;
	signal G5482: std_logic; attribute dont_touch of G5482: signal is true;
	signal G5483: std_logic; attribute dont_touch of G5483: signal is true;
	signal G5484: std_logic; attribute dont_touch of G5484: signal is true;
	signal G5485: std_logic; attribute dont_touch of G5485: signal is true;
	signal G5486: std_logic; attribute dont_touch of G5486: signal is true;
	signal G5489: std_logic; attribute dont_touch of G5489: signal is true;
	signal G5490: std_logic; attribute dont_touch of G5490: signal is true;
	signal G5491: std_logic; attribute dont_touch of G5491: signal is true;
	signal G5492: std_logic; attribute dont_touch of G5492: signal is true;
	signal G5493: std_logic; attribute dont_touch of G5493: signal is true;
	signal G5494: std_logic; attribute dont_touch of G5494: signal is true;
	signal G5497: std_logic; attribute dont_touch of G5497: signal is true;
	signal G5498: std_logic; attribute dont_touch of G5498: signal is true;
	signal G5499: std_logic; attribute dont_touch of G5499: signal is true;
	signal G5500: std_logic; attribute dont_touch of G5500: signal is true;
	signal G5501: std_logic; attribute dont_touch of G5501: signal is true;
	signal G5502: std_logic; attribute dont_touch of G5502: signal is true;
	signal G5503: std_logic; attribute dont_touch of G5503: signal is true;
	signal G5504: std_logic; attribute dont_touch of G5504: signal is true;
	signal G5507: std_logic; attribute dont_touch of G5507: signal is true;
	signal G5508: std_logic; attribute dont_touch of G5508: signal is true;
	signal G5509: std_logic; attribute dont_touch of G5509: signal is true;
	signal G5510: std_logic; attribute dont_touch of G5510: signal is true;
	signal G5511: std_logic; attribute dont_touch of G5511: signal is true;
	signal G5512: std_logic; attribute dont_touch of G5512: signal is true;
	signal G5513: std_logic; attribute dont_touch of G5513: signal is true;
	signal G5514: std_logic; attribute dont_touch of G5514: signal is true;
	signal G5515: std_logic; attribute dont_touch of G5515: signal is true;
	signal G5518: std_logic; attribute dont_touch of G5518: signal is true;
	signal G5519: std_logic; attribute dont_touch of G5519: signal is true;
	signal G5520: std_logic; attribute dont_touch of G5520: signal is true;
	signal G5521: std_logic; attribute dont_touch of G5521: signal is true;
	signal G5522: std_logic; attribute dont_touch of G5522: signal is true;
	signal G5523: std_logic; attribute dont_touch of G5523: signal is true;
	signal G5524: std_logic; attribute dont_touch of G5524: signal is true;
	signal G5525: std_logic; attribute dont_touch of G5525: signal is true;
	signal G5526: std_logic; attribute dont_touch of G5526: signal is true;
	signal G5527: std_logic; attribute dont_touch of G5527: signal is true;
	signal G5528: std_logic; attribute dont_touch of G5528: signal is true;
	signal G5529: std_logic; attribute dont_touch of G5529: signal is true;
	signal G5530: std_logic; attribute dont_touch of G5530: signal is true;
	signal G5531: std_logic; attribute dont_touch of G5531: signal is true;
	signal G5532: std_logic; attribute dont_touch of G5532: signal is true;
	signal G5533: std_logic; attribute dont_touch of G5533: signal is true;
	signal G5534: std_logic; attribute dont_touch of G5534: signal is true;
	signal G5535: std_logic; attribute dont_touch of G5535: signal is true;
	signal G5536: std_logic; attribute dont_touch of G5536: signal is true;
	signal G5537: std_logic; attribute dont_touch of G5537: signal is true;
	signal G5538: std_logic; attribute dont_touch of G5538: signal is true;
	signal G5539: std_logic; attribute dont_touch of G5539: signal is true;
	signal G5540: std_logic; attribute dont_touch of G5540: signal is true;
	signal G5541: std_logic; attribute dont_touch of G5541: signal is true;
	signal G5542: std_logic; attribute dont_touch of G5542: signal is true;
	signal G5543: std_logic; attribute dont_touch of G5543: signal is true;
	signal G5544: std_logic; attribute dont_touch of G5544: signal is true;
	signal G5545: std_logic; attribute dont_touch of G5545: signal is true;
	signal G5546: std_logic; attribute dont_touch of G5546: signal is true;
	signal G5547: std_logic; attribute dont_touch of G5547: signal is true;
	signal G5548: std_logic; attribute dont_touch of G5548: signal is true;
	signal G5552: std_logic; attribute dont_touch of G5552: signal is true;
	signal G5555: std_logic; attribute dont_touch of G5555: signal is true;
	signal G5556: std_logic; attribute dont_touch of G5556: signal is true;
	signal G5557: std_logic; attribute dont_touch of G5557: signal is true;
	signal G5567: std_logic; attribute dont_touch of G5567: signal is true;
	signal G5568: std_logic; attribute dont_touch of G5568: signal is true;
	signal G5569: std_logic; attribute dont_touch of G5569: signal is true;
	signal G5572: std_logic; attribute dont_touch of G5572: signal is true;
	signal G5573: std_logic; attribute dont_touch of G5573: signal is true;
	signal G5574: std_logic; attribute dont_touch of G5574: signal is true;
	signal G5575: std_logic; attribute dont_touch of G5575: signal is true;
	signal G5576: std_logic; attribute dont_touch of G5576: signal is true;
	signal G5586: std_logic; attribute dont_touch of G5586: signal is true;
	signal G5587: std_logic; attribute dont_touch of G5587: signal is true;
	signal G5588: std_logic; attribute dont_touch of G5588: signal is true;
	signal G5589: std_logic; attribute dont_touch of G5589: signal is true;
	signal G5590: std_logic; attribute dont_touch of G5590: signal is true;
	signal G5591: std_logic; attribute dont_touch of G5591: signal is true;
	signal G5592: std_logic; attribute dont_touch of G5592: signal is true;
	signal G5593: std_logic; attribute dont_touch of G5593: signal is true;
	signal G5594: std_logic; attribute dont_touch of G5594: signal is true;
	signal G5595: std_logic; attribute dont_touch of G5595: signal is true;
	signal G5596: std_logic; attribute dont_touch of G5596: signal is true;
	signal G5597: std_logic; attribute dont_touch of G5597: signal is true;
	signal G5598: std_logic; attribute dont_touch of G5598: signal is true;
	signal G5601: std_logic; attribute dont_touch of G5601: signal is true;
	signal G5602: std_logic; attribute dont_touch of G5602: signal is true;
	signal G5603: std_logic; attribute dont_touch of G5603: signal is true;
	signal G5604: std_logic; attribute dont_touch of G5604: signal is true;
	signal G5605: std_logic; attribute dont_touch of G5605: signal is true;
	signal G5608: std_logic; attribute dont_touch of G5608: signal is true;
	signal G5611: std_logic; attribute dont_touch of G5611: signal is true;
	signal G5612: std_logic; attribute dont_touch of G5612: signal is true;
	signal G5613: std_logic; attribute dont_touch of G5613: signal is true;
	signal G5614: std_logic; attribute dont_touch of G5614: signal is true;
	signal G5615: std_logic; attribute dont_touch of G5615: signal is true;
	signal G5616: std_logic; attribute dont_touch of G5616: signal is true;
	signal G5617: std_logic; attribute dont_touch of G5617: signal is true;
	signal G5618: std_logic; attribute dont_touch of G5618: signal is true;
	signal G5619: std_logic; attribute dont_touch of G5619: signal is true;
	signal G5620: std_logic; attribute dont_touch of G5620: signal is true;
	signal G5623: std_logic; attribute dont_touch of G5623: signal is true;
	signal G5624: std_logic; attribute dont_touch of G5624: signal is true;
	signal G5625: std_logic; attribute dont_touch of G5625: signal is true;
	signal G5626: std_logic; attribute dont_touch of G5626: signal is true;
	signal G5627: std_logic; attribute dont_touch of G5627: signal is true;
	signal G5628: std_logic; attribute dont_touch of G5628: signal is true;
	signal G5629: std_logic; attribute dont_touch of G5629: signal is true;
	signal G5630: std_logic; attribute dont_touch of G5630: signal is true;
	signal G5631: std_logic; attribute dont_touch of G5631: signal is true;
	signal G5632: std_logic; attribute dont_touch of G5632: signal is true;
	signal G5633: std_logic; attribute dont_touch of G5633: signal is true;
	signal G5637: std_logic; attribute dont_touch of G5637: signal is true;
	signal G5638: std_logic; attribute dont_touch of G5638: signal is true;
	signal G5639: std_logic; attribute dont_touch of G5639: signal is true;
	signal G5640: std_logic; attribute dont_touch of G5640: signal is true;
	signal G5641: std_logic; attribute dont_touch of G5641: signal is true;
	signal G5642: std_logic; attribute dont_touch of G5642: signal is true;
	signal G5643: std_logic; attribute dont_touch of G5643: signal is true;
	signal G5644: std_logic; attribute dont_touch of G5644: signal is true;
	signal G5645: std_logic; attribute dont_touch of G5645: signal is true;
	signal G5646: std_logic; attribute dont_touch of G5646: signal is true;
	signal G5647: std_logic; attribute dont_touch of G5647: signal is true;
	signal G5648: std_logic; attribute dont_touch of G5648: signal is true;
	signal G5649: std_logic; attribute dont_touch of G5649: signal is true;
	signal G5650: std_logic; attribute dont_touch of G5650: signal is true;
	signal G5651: std_logic; attribute dont_touch of G5651: signal is true;
	signal G5652: std_logic; attribute dont_touch of G5652: signal is true;
	signal G5653: std_logic; attribute dont_touch of G5653: signal is true;
	signal G5654: std_logic; attribute dont_touch of G5654: signal is true;
	signal G5655: std_logic; attribute dont_touch of G5655: signal is true;
	signal G5656: std_logic; attribute dont_touch of G5656: signal is true;
	signal G5657: std_logic; attribute dont_touch of G5657: signal is true;
	signal G5660: std_logic; attribute dont_touch of G5660: signal is true;
	signal G5661: std_logic; attribute dont_touch of G5661: signal is true;
	signal G5662: std_logic; attribute dont_touch of G5662: signal is true;
	signal G5663: std_logic; attribute dont_touch of G5663: signal is true;
	signal G5664: std_logic; attribute dont_touch of G5664: signal is true;
	signal G5665: std_logic; attribute dont_touch of G5665: signal is true;
	signal G5666: std_logic; attribute dont_touch of G5666: signal is true;
	signal G5667: std_logic; attribute dont_touch of G5667: signal is true;
	signal G5668: std_logic; attribute dont_touch of G5668: signal is true;
	signal G5669: std_logic; attribute dont_touch of G5669: signal is true;
	signal G5670: std_logic; attribute dont_touch of G5670: signal is true;
	signal G5671: std_logic; attribute dont_touch of G5671: signal is true;
	signal G5672: std_logic; attribute dont_touch of G5672: signal is true;
	signal G5673: std_logic; attribute dont_touch of G5673: signal is true;
	signal G5674: std_logic; attribute dont_touch of G5674: signal is true;
	signal G5675: std_logic; attribute dont_touch of G5675: signal is true;
	signal G5676: std_logic; attribute dont_touch of G5676: signal is true;
	signal G5677: std_logic; attribute dont_touch of G5677: signal is true;
	signal G5678: std_logic; attribute dont_touch of G5678: signal is true;
	signal G5679: std_logic; attribute dont_touch of G5679: signal is true;
	signal G5680: std_logic; attribute dont_touch of G5680: signal is true;
	signal G5681: std_logic; attribute dont_touch of G5681: signal is true;
	signal G5682: std_logic; attribute dont_touch of G5682: signal is true;
	signal G5683: std_logic; attribute dont_touch of G5683: signal is true;
	signal G5684: std_logic; attribute dont_touch of G5684: signal is true;
	signal G5685: std_logic; attribute dont_touch of G5685: signal is true;
	signal G5686: std_logic; attribute dont_touch of G5686: signal is true;
	signal G5687: std_logic; attribute dont_touch of G5687: signal is true;
	signal G5688: std_logic; attribute dont_touch of G5688: signal is true;
	signal G5689: std_logic; attribute dont_touch of G5689: signal is true;
	signal G5690: std_logic; attribute dont_touch of G5690: signal is true;
	signal G5691: std_logic; attribute dont_touch of G5691: signal is true;
	signal G5692: std_logic; attribute dont_touch of G5692: signal is true;
	signal G5693: std_logic; attribute dont_touch of G5693: signal is true;
	signal G5694: std_logic; attribute dont_touch of G5694: signal is true;
	signal G5695: std_logic; attribute dont_touch of G5695: signal is true;
	signal G5696: std_logic; attribute dont_touch of G5696: signal is true;
	signal G5697: std_logic; attribute dont_touch of G5697: signal is true;
	signal G5698: std_logic; attribute dont_touch of G5698: signal is true;
	signal G5699: std_logic; attribute dont_touch of G5699: signal is true;
	signal G5700: std_logic; attribute dont_touch of G5700: signal is true;
	signal G5701: std_logic; attribute dont_touch of G5701: signal is true;
	signal G5702: std_logic; attribute dont_touch of G5702: signal is true;
	signal G5703: std_logic; attribute dont_touch of G5703: signal is true;
	signal G5704: std_logic; attribute dont_touch of G5704: signal is true;
	signal G5705: std_logic; attribute dont_touch of G5705: signal is true;
	signal G5706: std_logic; attribute dont_touch of G5706: signal is true;
	signal G5707: std_logic; attribute dont_touch of G5707: signal is true;
	signal G5708: std_logic; attribute dont_touch of G5708: signal is true;
	signal G5718: std_logic; attribute dont_touch of G5718: signal is true;
	signal G5719: std_logic; attribute dont_touch of G5719: signal is true;
	signal G5720: std_logic; attribute dont_touch of G5720: signal is true;
	signal G5721: std_logic; attribute dont_touch of G5721: signal is true;
	signal G5722: std_logic; attribute dont_touch of G5722: signal is true;
	signal G5723: std_logic; attribute dont_touch of G5723: signal is true;
	signal G5724: std_logic; attribute dont_touch of G5724: signal is true;
	signal G5725: std_logic; attribute dont_touch of G5725: signal is true;
	signal G5726: std_logic; attribute dont_touch of G5726: signal is true;
	signal G5727: std_logic; attribute dont_touch of G5727: signal is true;
	signal G5728: std_logic; attribute dont_touch of G5728: signal is true;
	signal G5729: std_logic; attribute dont_touch of G5729: signal is true;
	signal G5730: std_logic; attribute dont_touch of G5730: signal is true;
	signal G5731: std_logic; attribute dont_touch of G5731: signal is true;
	signal G5732: std_logic; attribute dont_touch of G5732: signal is true;
	signal G5733: std_logic; attribute dont_touch of G5733: signal is true;
	signal G5734: std_logic; attribute dont_touch of G5734: signal is true;
	signal G5735: std_logic; attribute dont_touch of G5735: signal is true;
	signal G5736: std_logic; attribute dont_touch of G5736: signal is true;
	signal G5737: std_logic; attribute dont_touch of G5737: signal is true;
	signal G5738: std_logic; attribute dont_touch of G5738: signal is true;
	signal G5739: std_logic; attribute dont_touch of G5739: signal is true;
	signal G5740: std_logic; attribute dont_touch of G5740: signal is true;
	signal G5741: std_logic; attribute dont_touch of G5741: signal is true;
	signal G5742: std_logic; attribute dont_touch of G5742: signal is true;
	signal G5743: std_logic; attribute dont_touch of G5743: signal is true;
	signal G5744: std_logic; attribute dont_touch of G5744: signal is true;
	signal G5745: std_logic; attribute dont_touch of G5745: signal is true;
	signal G5746: std_logic; attribute dont_touch of G5746: signal is true;
	signal G5747: std_logic; attribute dont_touch of G5747: signal is true;
	signal G5748: std_logic; attribute dont_touch of G5748: signal is true;
	signal G5751: std_logic; attribute dont_touch of G5751: signal is true;
	signal G5752: std_logic; attribute dont_touch of G5752: signal is true;
	signal G5753: std_logic; attribute dont_touch of G5753: signal is true;
	signal G5754: std_logic; attribute dont_touch of G5754: signal is true;
	signal G5755: std_logic; attribute dont_touch of G5755: signal is true;
	signal G5756: std_logic; attribute dont_touch of G5756: signal is true;
	signal G5757: std_logic; attribute dont_touch of G5757: signal is true;
	signal G5758: std_logic; attribute dont_touch of G5758: signal is true;
	signal G5759: std_logic; attribute dont_touch of G5759: signal is true;
	signal G5762: std_logic; attribute dont_touch of G5762: signal is true;
	signal G5763: std_logic; attribute dont_touch of G5763: signal is true;
	signal G5766: std_logic; attribute dont_touch of G5766: signal is true;
	signal G5767: std_logic; attribute dont_touch of G5767: signal is true;
	signal G5768: std_logic; attribute dont_touch of G5768: signal is true;
	signal G5769: std_logic; attribute dont_touch of G5769: signal is true;
	signal G5770: std_logic; attribute dont_touch of G5770: signal is true;
	signal G5771: std_logic; attribute dont_touch of G5771: signal is true;
	signal G5772: std_logic; attribute dont_touch of G5772: signal is true;
	signal G5773: std_logic; attribute dont_touch of G5773: signal is true;
	signal G5774: std_logic; attribute dont_touch of G5774: signal is true;
	signal G5777: std_logic; attribute dont_touch of G5777: signal is true;
	signal G5778: std_logic; attribute dont_touch of G5778: signal is true;
	signal G5779: std_logic; attribute dont_touch of G5779: signal is true;
	signal G5780: std_logic; attribute dont_touch of G5780: signal is true;
	signal G5781: std_logic; attribute dont_touch of G5781: signal is true;
	signal G5782: std_logic; attribute dont_touch of G5782: signal is true;
	signal G5783: std_logic; attribute dont_touch of G5783: signal is true;
	signal G5784: std_logic; attribute dont_touch of G5784: signal is true;
	signal G5787: std_logic; attribute dont_touch of G5787: signal is true;
	signal G5788: std_logic; attribute dont_touch of G5788: signal is true;
	signal G5789: std_logic; attribute dont_touch of G5789: signal is true;
	signal G5790: std_logic; attribute dont_touch of G5790: signal is true;
	signal G5791: std_logic; attribute dont_touch of G5791: signal is true;
	signal G5794: std_logic; attribute dont_touch of G5794: signal is true;
	signal G5795: std_logic; attribute dont_touch of G5795: signal is true;
	signal G5796: std_logic; attribute dont_touch of G5796: signal is true;
	signal G5797: std_logic; attribute dont_touch of G5797: signal is true;
	signal G5800: std_logic; attribute dont_touch of G5800: signal is true;
	signal G5801: std_logic; attribute dont_touch of G5801: signal is true;
	signal G5802: std_logic; attribute dont_touch of G5802: signal is true;
	signal G5803: std_logic; attribute dont_touch of G5803: signal is true;
	signal G5804: std_logic; attribute dont_touch of G5804: signal is true;
	signal G5805: std_logic; attribute dont_touch of G5805: signal is true;
	signal G5808: std_logic; attribute dont_touch of G5808: signal is true;
	signal G5809: std_logic; attribute dont_touch of G5809: signal is true;
	signal G5810: std_logic; attribute dont_touch of G5810: signal is true;
	signal G5811: std_logic; attribute dont_touch of G5811: signal is true;
	signal G5812: std_logic; attribute dont_touch of G5812: signal is true;
	signal G5813: std_logic; attribute dont_touch of G5813: signal is true;
	signal G5814: std_logic; attribute dont_touch of G5814: signal is true;
	signal G5815: std_logic; attribute dont_touch of G5815: signal is true;
	signal G5817: std_logic; attribute dont_touch of G5817: signal is true;
	signal G5818: std_logic; attribute dont_touch of G5818: signal is true;
	signal G5819: std_logic; attribute dont_touch of G5819: signal is true;
	signal G5820: std_logic; attribute dont_touch of G5820: signal is true;
	signal G5821: std_logic; attribute dont_touch of G5821: signal is true;
	signal G5822: std_logic; attribute dont_touch of G5822: signal is true;
	signal G5823: std_logic; attribute dont_touch of G5823: signal is true;
	signal G5824: std_logic; attribute dont_touch of G5824: signal is true;
	signal G5825: std_logic; attribute dont_touch of G5825: signal is true;
	signal G5826: std_logic; attribute dont_touch of G5826: signal is true;
	signal G5827: std_logic; attribute dont_touch of G5827: signal is true;
	signal G5830: std_logic; attribute dont_touch of G5830: signal is true;
	signal G5836: std_logic; attribute dont_touch of G5836: signal is true;
	signal G5837: std_logic; attribute dont_touch of G5837: signal is true;
	signal G5838: std_logic; attribute dont_touch of G5838: signal is true;
	signal G5839: std_logic; attribute dont_touch of G5839: signal is true;
	signal G5840: std_logic; attribute dont_touch of G5840: signal is true;
	signal G5841: std_logic; attribute dont_touch of G5841: signal is true;
	signal G5842: std_logic; attribute dont_touch of G5842: signal is true;
	signal G5843: std_logic; attribute dont_touch of G5843: signal is true;
	signal G5844: std_logic; attribute dont_touch of G5844: signal is true;
	signal G5845: std_logic; attribute dont_touch of G5845: signal is true;
	signal G5846: std_logic; attribute dont_touch of G5846: signal is true;
	signal G5847: std_logic; attribute dont_touch of G5847: signal is true;
	signal G5848: std_logic; attribute dont_touch of G5848: signal is true;
	signal G5849: std_logic; attribute dont_touch of G5849: signal is true;
	signal G5850: std_logic; attribute dont_touch of G5850: signal is true;
	signal G5851: std_logic; attribute dont_touch of G5851: signal is true;
	signal G5852: std_logic; attribute dont_touch of G5852: signal is true;
	signal G5853: std_logic; attribute dont_touch of G5853: signal is true;
	signal G5856: std_logic; attribute dont_touch of G5856: signal is true;
	signal G5857: std_logic; attribute dont_touch of G5857: signal is true;
	signal G5858: std_logic; attribute dont_touch of G5858: signal is true;
	signal G5859: std_logic; attribute dont_touch of G5859: signal is true;
	signal G5862: std_logic; attribute dont_touch of G5862: signal is true;
	signal G5863: std_logic; attribute dont_touch of G5863: signal is true;
	signal G5864: std_logic; attribute dont_touch of G5864: signal is true;
	signal G5865: std_logic; attribute dont_touch of G5865: signal is true;
	signal G5866: std_logic; attribute dont_touch of G5866: signal is true;
	signal G5867: std_logic; attribute dont_touch of G5867: signal is true;
	signal G5874: std_logic; attribute dont_touch of G5874: signal is true;
	signal G5875: std_logic; attribute dont_touch of G5875: signal is true;
	signal G5876: std_logic; attribute dont_touch of G5876: signal is true;
	signal G5877: std_logic; attribute dont_touch of G5877: signal is true;
	signal G5878: std_logic; attribute dont_touch of G5878: signal is true;
	signal G5879: std_logic; attribute dont_touch of G5879: signal is true;
	signal G5880: std_logic; attribute dont_touch of G5880: signal is true;
	signal G5881: std_logic; attribute dont_touch of G5881: signal is true;
	signal G5882: std_logic; attribute dont_touch of G5882: signal is true;
	signal G5883: std_logic; attribute dont_touch of G5883: signal is true;
	signal G5884: std_logic; attribute dont_touch of G5884: signal is true;
	signal G5885: std_logic; attribute dont_touch of G5885: signal is true;
	signal G5886: std_logic; attribute dont_touch of G5886: signal is true;
	signal G5887: std_logic; attribute dont_touch of G5887: signal is true;
	signal G5888: std_logic; attribute dont_touch of G5888: signal is true;
	signal G5889: std_logic; attribute dont_touch of G5889: signal is true;
	signal G5890: std_logic; attribute dont_touch of G5890: signal is true;
	signal G5891: std_logic; attribute dont_touch of G5891: signal is true;
	signal G5892: std_logic; attribute dont_touch of G5892: signal is true;
	signal G5893: std_logic; attribute dont_touch of G5893: signal is true;
	signal G5894: std_logic; attribute dont_touch of G5894: signal is true;
	signal G5895: std_logic; attribute dont_touch of G5895: signal is true;
	signal G5896: std_logic; attribute dont_touch of G5896: signal is true;
	signal G5897: std_logic; attribute dont_touch of G5897: signal is true;
	signal G5898: std_logic; attribute dont_touch of G5898: signal is true;
	signal G5899: std_logic; attribute dont_touch of G5899: signal is true;
	signal G5900: std_logic; attribute dont_touch of G5900: signal is true;
	signal G5901: std_logic; attribute dont_touch of G5901: signal is true;
	signal G5902: std_logic; attribute dont_touch of G5902: signal is true;
	signal G5903: std_logic; attribute dont_touch of G5903: signal is true;
	signal G5904: std_logic; attribute dont_touch of G5904: signal is true;
	signal G5910: std_logic; attribute dont_touch of G5910: signal is true;
	signal G5911: std_logic; attribute dont_touch of G5911: signal is true;
	signal G5912: std_logic; attribute dont_touch of G5912: signal is true;
	signal G5913: std_logic; attribute dont_touch of G5913: signal is true;
	signal G5914: std_logic; attribute dont_touch of G5914: signal is true;
	signal G5915: std_logic; attribute dont_touch of G5915: signal is true;
	signal G5916: std_logic; attribute dont_touch of G5916: signal is true;
	signal G5917: std_logic; attribute dont_touch of G5917: signal is true;
	signal G5918: std_logic; attribute dont_touch of G5918: signal is true;
	signal G5919: std_logic; attribute dont_touch of G5919: signal is true;
	signal G5934: std_logic; attribute dont_touch of G5934: signal is true;
	signal G5935: std_logic; attribute dont_touch of G5935: signal is true;
	signal G5936: std_logic; attribute dont_touch of G5936: signal is true;
	signal G5937: std_logic; attribute dont_touch of G5937: signal is true;
	signal G5938: std_logic; attribute dont_touch of G5938: signal is true;
	signal G5941: std_logic; attribute dont_touch of G5941: signal is true;
	signal G5942: std_logic; attribute dont_touch of G5942: signal is true;
	signal G5943: std_logic; attribute dont_touch of G5943: signal is true;
	signal G5944: std_logic; attribute dont_touch of G5944: signal is true;
	signal G5947: std_logic; attribute dont_touch of G5947: signal is true;
	signal G5948: std_logic; attribute dont_touch of G5948: signal is true;
	signal G5949: std_logic; attribute dont_touch of G5949: signal is true;
	signal G5980: std_logic; attribute dont_touch of G5980: signal is true;
	signal G5981: std_logic; attribute dont_touch of G5981: signal is true;
	signal G5982: std_logic; attribute dont_touch of G5982: signal is true;
	signal G5983: std_logic; attribute dont_touch of G5983: signal is true;
	signal G5984: std_logic; attribute dont_touch of G5984: signal is true;
	signal G5987: std_logic; attribute dont_touch of G5987: signal is true;
	signal G5992: std_logic; attribute dont_touch of G5992: signal is true;
	signal G5993: std_logic; attribute dont_touch of G5993: signal is true;
	signal G5994: std_logic; attribute dont_touch of G5994: signal is true;
	signal G5995: std_logic; attribute dont_touch of G5995: signal is true;
	signal G5996: std_logic; attribute dont_touch of G5996: signal is true;
	signal G5997: std_logic; attribute dont_touch of G5997: signal is true;
	signal G5998: std_logic; attribute dont_touch of G5998: signal is true;
	signal G5999: std_logic; attribute dont_touch of G5999: signal is true;
	signal G6000: std_logic; attribute dont_touch of G6000: signal is true;
	signal G6001: std_logic; attribute dont_touch of G6001: signal is true;
	signal G6002: std_logic; attribute dont_touch of G6002: signal is true;
	signal G6003: std_logic; attribute dont_touch of G6003: signal is true;
	signal G6014: std_logic; attribute dont_touch of G6014: signal is true;
	signal G6015: std_logic; attribute dont_touch of G6015: signal is true;
	signal G6016: std_logic; attribute dont_touch of G6016: signal is true;
	signal G6019: std_logic; attribute dont_touch of G6019: signal is true;
	signal G6023: std_logic; attribute dont_touch of G6023: signal is true;
	signal G6026: std_logic; attribute dont_touch of G6026: signal is true;
	signal G6027: std_logic; attribute dont_touch of G6027: signal is true;
	signal G6030: std_logic; attribute dont_touch of G6030: signal is true;
	signal G6031: std_logic; attribute dont_touch of G6031: signal is true;
	signal G6032: std_logic; attribute dont_touch of G6032: signal is true;
	signal G6035: std_logic; attribute dont_touch of G6035: signal is true;
	signal G6036: std_logic; attribute dont_touch of G6036: signal is true;
	signal G6037: std_logic; attribute dont_touch of G6037: signal is true;
	signal G6038: std_logic; attribute dont_touch of G6038: signal is true;
	signal G6039: std_logic; attribute dont_touch of G6039: signal is true;
	signal G6040: std_logic; attribute dont_touch of G6040: signal is true;
	signal G6041: std_logic; attribute dont_touch of G6041: signal is true;
	signal G6042: std_logic; attribute dont_touch of G6042: signal is true;
	signal G6043: std_logic; attribute dont_touch of G6043: signal is true;
	signal G6044: std_logic; attribute dont_touch of G6044: signal is true;
	signal G6045: std_logic; attribute dont_touch of G6045: signal is true;
	signal G6046: std_logic; attribute dont_touch of G6046: signal is true;
	signal G6047: std_logic; attribute dont_touch of G6047: signal is true;
	signal G6048: std_logic; attribute dont_touch of G6048: signal is true;
	signal G6049: std_logic; attribute dont_touch of G6049: signal is true;
	signal G6050: std_logic; attribute dont_touch of G6050: signal is true;
	signal G6051: std_logic; attribute dont_touch of G6051: signal is true;
	signal G6052: std_logic; attribute dont_touch of G6052: signal is true;
	signal G6053: std_logic; attribute dont_touch of G6053: signal is true;
	signal G6054: std_logic; attribute dont_touch of G6054: signal is true;
	signal G6055: std_logic; attribute dont_touch of G6055: signal is true;
	signal G6056: std_logic; attribute dont_touch of G6056: signal is true;
	signal G6057: std_logic; attribute dont_touch of G6057: signal is true;
	signal G6058: std_logic; attribute dont_touch of G6058: signal is true;
	signal G6059: std_logic; attribute dont_touch of G6059: signal is true;
	signal G6060: std_logic; attribute dont_touch of G6060: signal is true;
	signal G6061: std_logic; attribute dont_touch of G6061: signal is true;
	signal G6062: std_logic; attribute dont_touch of G6062: signal is true;
	signal G6063: std_logic; attribute dont_touch of G6063: signal is true;
	signal G6064: std_logic; attribute dont_touch of G6064: signal is true;
	signal G6067: std_logic; attribute dont_touch of G6067: signal is true;
	signal G6068: std_logic; attribute dont_touch of G6068: signal is true;
	signal G6069: std_logic; attribute dont_touch of G6069: signal is true;
	signal G6070: std_logic; attribute dont_touch of G6070: signal is true;
	signal G6071: std_logic; attribute dont_touch of G6071: signal is true;
	signal G6072: std_logic; attribute dont_touch of G6072: signal is true;
	signal G6073: std_logic; attribute dont_touch of G6073: signal is true;
	signal G6074: std_logic; attribute dont_touch of G6074: signal is true;
	signal G6075: std_logic; attribute dont_touch of G6075: signal is true;
	signal G6076: std_logic; attribute dont_touch of G6076: signal is true;
	signal G6077: std_logic; attribute dont_touch of G6077: signal is true;
	signal G6078: std_logic; attribute dont_touch of G6078: signal is true;
	signal G6079: std_logic; attribute dont_touch of G6079: signal is true;
	signal G6080: std_logic; attribute dont_touch of G6080: signal is true;
	signal G6081: std_logic; attribute dont_touch of G6081: signal is true;
	signal G6082: std_logic; attribute dont_touch of G6082: signal is true;
	signal G6083: std_logic; attribute dont_touch of G6083: signal is true;
	signal G6084: std_logic; attribute dont_touch of G6084: signal is true;
	signal G6085: std_logic; attribute dont_touch of G6085: signal is true;
	signal G6086: std_logic; attribute dont_touch of G6086: signal is true;
	signal G6087: std_logic; attribute dont_touch of G6087: signal is true;
	signal G6088: std_logic; attribute dont_touch of G6088: signal is true;
	signal G6089: std_logic; attribute dont_touch of G6089: signal is true;
	signal G6090: std_logic; attribute dont_touch of G6090: signal is true;
	signal G6091: std_logic; attribute dont_touch of G6091: signal is true;
	signal G6092: std_logic; attribute dont_touch of G6092: signal is true;
	signal G6093: std_logic; attribute dont_touch of G6093: signal is true;
	signal G6094: std_logic; attribute dont_touch of G6094: signal is true;
	signal G6095: std_logic; attribute dont_touch of G6095: signal is true;
	signal G6096: std_logic; attribute dont_touch of G6096: signal is true;
	signal G6097: std_logic; attribute dont_touch of G6097: signal is true;
	signal G6098: std_logic; attribute dont_touch of G6098: signal is true;
	signal G6099: std_logic; attribute dont_touch of G6099: signal is true;
	signal G6100: std_logic; attribute dont_touch of G6100: signal is true;
	signal G6101: std_logic; attribute dont_touch of G6101: signal is true;
	signal G6102: std_logic; attribute dont_touch of G6102: signal is true;
	signal G6103: std_logic; attribute dont_touch of G6103: signal is true;
	signal G6104: std_logic; attribute dont_touch of G6104: signal is true;
	signal G6105: std_logic; attribute dont_touch of G6105: signal is true;
	signal G6106: std_logic; attribute dont_touch of G6106: signal is true;
	signal G6107: std_logic; attribute dont_touch of G6107: signal is true;
	signal G6108: std_logic; attribute dont_touch of G6108: signal is true;
	signal G6109: std_logic; attribute dont_touch of G6109: signal is true;
	signal G6110: std_logic; attribute dont_touch of G6110: signal is true;
	signal G6111: std_logic; attribute dont_touch of G6111: signal is true;
	signal G6112: std_logic; attribute dont_touch of G6112: signal is true;
	signal G6113: std_logic; attribute dont_touch of G6113: signal is true;
	signal G6114: std_logic; attribute dont_touch of G6114: signal is true;
	signal G6115: std_logic; attribute dont_touch of G6115: signal is true;
	signal G6116: std_logic; attribute dont_touch of G6116: signal is true;
	signal G6117: std_logic; attribute dont_touch of G6117: signal is true;
	signal G6118: std_logic; attribute dont_touch of G6118: signal is true;
	signal G6119: std_logic; attribute dont_touch of G6119: signal is true;
	signal G6120: std_logic; attribute dont_touch of G6120: signal is true;
	signal G6121: std_logic; attribute dont_touch of G6121: signal is true;
	signal G6122: std_logic; attribute dont_touch of G6122: signal is true;
	signal G6123: std_logic; attribute dont_touch of G6123: signal is true;
	signal G6124: std_logic; attribute dont_touch of G6124: signal is true;
	signal G6125: std_logic; attribute dont_touch of G6125: signal is true;
	signal G6126: std_logic; attribute dont_touch of G6126: signal is true;
	signal G6127: std_logic; attribute dont_touch of G6127: signal is true;
	signal G6128: std_logic; attribute dont_touch of G6128: signal is true;
	signal G6131: std_logic; attribute dont_touch of G6131: signal is true;
	signal G6132: std_logic; attribute dont_touch of G6132: signal is true;
	signal G6133: std_logic; attribute dont_touch of G6133: signal is true;
	signal G6134: std_logic; attribute dont_touch of G6134: signal is true;
	signal G6135: std_logic; attribute dont_touch of G6135: signal is true;
	signal G6136: std_logic; attribute dont_touch of G6136: signal is true;
	signal G6137: std_logic; attribute dont_touch of G6137: signal is true;
	signal G6140: std_logic; attribute dont_touch of G6140: signal is true;
	signal G6141: std_logic; attribute dont_touch of G6141: signal is true;
	signal G6144: std_logic; attribute dont_touch of G6144: signal is true;
	signal G6145: std_logic; attribute dont_touch of G6145: signal is true;
	signal G6146: std_logic; attribute dont_touch of G6146: signal is true;
	signal G6149: std_logic; attribute dont_touch of G6149: signal is true;
	signal G6150: std_logic; attribute dont_touch of G6150: signal is true;
	signal G6151: std_logic; attribute dont_touch of G6151: signal is true;
	signal G6154: std_logic; attribute dont_touch of G6154: signal is true;
	signal G6155: std_logic; attribute dont_touch of G6155: signal is true;
	signal G6156: std_logic; attribute dont_touch of G6156: signal is true;
	signal G6157: std_logic; attribute dont_touch of G6157: signal is true;
	signal G6158: std_logic; attribute dont_touch of G6158: signal is true;
	signal G6161: std_logic; attribute dont_touch of G6161: signal is true;
	signal G6162: std_logic; attribute dont_touch of G6162: signal is true;
	signal G6163: std_logic; attribute dont_touch of G6163: signal is true;
	signal G6164: std_logic; attribute dont_touch of G6164: signal is true;
	signal G6165: std_logic; attribute dont_touch of G6165: signal is true;
	signal G6166: std_logic; attribute dont_touch of G6166: signal is true;
	signal G6169: std_logic; attribute dont_touch of G6169: signal is true;
	signal G6170: std_logic; attribute dont_touch of G6170: signal is true;
	signal G6171: std_logic; attribute dont_touch of G6171: signal is true;
	signal G6172: std_logic; attribute dont_touch of G6172: signal is true;
	signal G6175: std_logic; attribute dont_touch of G6175: signal is true;
	signal G6176: std_logic; attribute dont_touch of G6176: signal is true;
	signal G6177: std_logic; attribute dont_touch of G6177: signal is true;
	signal G6178: std_logic; attribute dont_touch of G6178: signal is true;
	signal G6179: std_logic; attribute dont_touch of G6179: signal is true;
	signal G6180: std_logic; attribute dont_touch of G6180: signal is true;
	signal G6181: std_logic; attribute dont_touch of G6181: signal is true;
	signal G6182: std_logic; attribute dont_touch of G6182: signal is true;
	signal G6183: std_logic; attribute dont_touch of G6183: signal is true;
	signal G6184: std_logic; attribute dont_touch of G6184: signal is true;
	signal G6185: std_logic; attribute dont_touch of G6185: signal is true;
	signal G6186: std_logic; attribute dont_touch of G6186: signal is true;
	signal G6187: std_logic; attribute dont_touch of G6187: signal is true;
	signal G6190: std_logic; attribute dont_touch of G6190: signal is true;
	signal G6191: std_logic; attribute dont_touch of G6191: signal is true;
	signal G6192: std_logic; attribute dont_touch of G6192: signal is true;
	signal G6193: std_logic; attribute dont_touch of G6193: signal is true;
	signal G6194: std_logic; attribute dont_touch of G6194: signal is true;
	signal G6195: std_logic; attribute dont_touch of G6195: signal is true;
	signal G6196: std_logic; attribute dont_touch of G6196: signal is true;
	signal G6197: std_logic; attribute dont_touch of G6197: signal is true;
	signal G6198: std_logic; attribute dont_touch of G6198: signal is true;
	signal G6199: std_logic; attribute dont_touch of G6199: signal is true;
	signal G6200: std_logic; attribute dont_touch of G6200: signal is true;
	signal G6201: std_logic; attribute dont_touch of G6201: signal is true;
	signal G6202: std_logic; attribute dont_touch of G6202: signal is true;
	signal G6203: std_logic; attribute dont_touch of G6203: signal is true;
	signal G6204: std_logic; attribute dont_touch of G6204: signal is true;
	signal G6205: std_logic; attribute dont_touch of G6205: signal is true;
	signal G6206: std_logic; attribute dont_touch of G6206: signal is true;
	signal G6207: std_logic; attribute dont_touch of G6207: signal is true;
	signal G6208: std_logic; attribute dont_touch of G6208: signal is true;
	signal G6209: std_logic; attribute dont_touch of G6209: signal is true;
	signal G6210: std_logic; attribute dont_touch of G6210: signal is true;
	signal G6213: std_logic; attribute dont_touch of G6213: signal is true;
	signal G6214: std_logic; attribute dont_touch of G6214: signal is true;
	signal G6215: std_logic; attribute dont_touch of G6215: signal is true;
	signal G6216: std_logic; attribute dont_touch of G6216: signal is true;
	signal G6217: std_logic; attribute dont_touch of G6217: signal is true;
	signal G6218: std_logic; attribute dont_touch of G6218: signal is true;
	signal G6219: std_logic; attribute dont_touch of G6219: signal is true;
	signal G6220: std_logic; attribute dont_touch of G6220: signal is true;
	signal G6221: std_logic; attribute dont_touch of G6221: signal is true;
	signal G6224: std_logic; attribute dont_touch of G6224: signal is true;
	signal G6225: std_logic; attribute dont_touch of G6225: signal is true;
	signal G6226: std_logic; attribute dont_touch of G6226: signal is true;
	signal G6227: std_logic; attribute dont_touch of G6227: signal is true;
	signal G6228: std_logic; attribute dont_touch of G6228: signal is true;
	signal G6231: std_logic; attribute dont_touch of G6231: signal is true;
	signal G6234: std_logic; attribute dont_touch of G6234: signal is true;
	signal G6235: std_logic; attribute dont_touch of G6235: signal is true;
	signal G6236: std_logic; attribute dont_touch of G6236: signal is true;
	signal G6237: std_logic; attribute dont_touch of G6237: signal is true;
	signal G6238: std_logic; attribute dont_touch of G6238: signal is true;
	signal G6239: std_logic; attribute dont_touch of G6239: signal is true;
	signal G6240: std_logic; attribute dont_touch of G6240: signal is true;
	signal G6241: std_logic; attribute dont_touch of G6241: signal is true;
	signal G6242: std_logic; attribute dont_touch of G6242: signal is true;
	signal G6243: std_logic; attribute dont_touch of G6243: signal is true;
	signal G6244: std_logic; attribute dont_touch of G6244: signal is true;
	signal G6245: std_logic; attribute dont_touch of G6245: signal is true;
	signal G6246: std_logic; attribute dont_touch of G6246: signal is true;
	signal G6247: std_logic; attribute dont_touch of G6247: signal is true;
	signal G6248: std_logic; attribute dont_touch of G6248: signal is true;
	signal G6249: std_logic; attribute dont_touch of G6249: signal is true;
	signal G6250: std_logic; attribute dont_touch of G6250: signal is true;
	signal G6251: std_logic; attribute dont_touch of G6251: signal is true;
	signal G6252: std_logic; attribute dont_touch of G6252: signal is true;
	signal G6286: std_logic; attribute dont_touch of G6286: signal is true;
	signal G6287: std_logic; attribute dont_touch of G6287: signal is true;
	signal G6288: std_logic; attribute dont_touch of G6288: signal is true;
	signal G6289: std_logic; attribute dont_touch of G6289: signal is true;
	signal G6290: std_logic; attribute dont_touch of G6290: signal is true;
	signal G6291: std_logic; attribute dont_touch of G6291: signal is true;
	signal G6292: std_logic; attribute dont_touch of G6292: signal is true;
	signal G6293: std_logic; attribute dont_touch of G6293: signal is true;
	signal G6294: std_logic; attribute dont_touch of G6294: signal is true;
	signal G6295: std_logic; attribute dont_touch of G6295: signal is true;
	signal G6296: std_logic; attribute dont_touch of G6296: signal is true;
	signal G6297: std_logic; attribute dont_touch of G6297: signal is true;
	signal G6298: std_logic; attribute dont_touch of G6298: signal is true;
	signal G6299: std_logic; attribute dont_touch of G6299: signal is true;
	signal G6300: std_logic; attribute dont_touch of G6300: signal is true;
	signal G6301: std_logic; attribute dont_touch of G6301: signal is true;
	signal G6302: std_logic; attribute dont_touch of G6302: signal is true;
	signal G6303: std_logic; attribute dont_touch of G6303: signal is true;
	signal G6304: std_logic; attribute dont_touch of G6304: signal is true;
	signal G6305: std_logic; attribute dont_touch of G6305: signal is true;
	signal G6306: std_logic; attribute dont_touch of G6306: signal is true;
	signal G6307: std_logic; attribute dont_touch of G6307: signal is true;
	signal G6308: std_logic; attribute dont_touch of G6308: signal is true;
	signal G6309: std_logic; attribute dont_touch of G6309: signal is true;
	signal G6310: std_logic; attribute dont_touch of G6310: signal is true;
	signal G6311: std_logic; attribute dont_touch of G6311: signal is true;
	signal G6312: std_logic; attribute dont_touch of G6312: signal is true;
	signal G6313: std_logic; attribute dont_touch of G6313: signal is true;
	signal G6314: std_logic; attribute dont_touch of G6314: signal is true;
	signal G6315: std_logic; attribute dont_touch of G6315: signal is true;
	signal G6316: std_logic; attribute dont_touch of G6316: signal is true;
	signal G6317: std_logic; attribute dont_touch of G6317: signal is true;
	signal G6318: std_logic; attribute dont_touch of G6318: signal is true;
	signal G6319: std_logic; attribute dont_touch of G6319: signal is true;
	signal G6320: std_logic; attribute dont_touch of G6320: signal is true;
	signal G6321: std_logic; attribute dont_touch of G6321: signal is true;
	signal G6322: std_logic; attribute dont_touch of G6322: signal is true;
	signal G6323: std_logic; attribute dont_touch of G6323: signal is true;
	signal G6324: std_logic; attribute dont_touch of G6324: signal is true;
	signal G6325: std_logic; attribute dont_touch of G6325: signal is true;
	signal G6326: std_logic; attribute dont_touch of G6326: signal is true;
	signal G6327: std_logic; attribute dont_touch of G6327: signal is true;
	signal G6328: std_logic; attribute dont_touch of G6328: signal is true;
	signal G6329: std_logic; attribute dont_touch of G6329: signal is true;
	signal G6330: std_logic; attribute dont_touch of G6330: signal is true;
	signal G6331: std_logic; attribute dont_touch of G6331: signal is true;
	signal G6332: std_logic; attribute dont_touch of G6332: signal is true;
	signal G6333: std_logic; attribute dont_touch of G6333: signal is true;
	signal G6334: std_logic; attribute dont_touch of G6334: signal is true;
	signal G6335: std_logic; attribute dont_touch of G6335: signal is true;
	signal G6336: std_logic; attribute dont_touch of G6336: signal is true;
	signal G6337: std_logic; attribute dont_touch of G6337: signal is true;
	signal G6338: std_logic; attribute dont_touch of G6338: signal is true;
	signal G6339: std_logic; attribute dont_touch of G6339: signal is true;
	signal G6340: std_logic; attribute dont_touch of G6340: signal is true;
	signal G6341: std_logic; attribute dont_touch of G6341: signal is true;
	signal G6342: std_logic; attribute dont_touch of G6342: signal is true;
	signal G6343: std_logic; attribute dont_touch of G6343: signal is true;
	signal G6344: std_logic; attribute dont_touch of G6344: signal is true;
	signal G6345: std_logic; attribute dont_touch of G6345: signal is true;
	signal G6346: std_logic; attribute dont_touch of G6346: signal is true;
	signal G6347: std_logic; attribute dont_touch of G6347: signal is true;
	signal G6348: std_logic; attribute dont_touch of G6348: signal is true;
	signal G6349: std_logic; attribute dont_touch of G6349: signal is true;
	signal G6350: std_logic; attribute dont_touch of G6350: signal is true;
	signal G6351: std_logic; attribute dont_touch of G6351: signal is true;
	signal G6352: std_logic; attribute dont_touch of G6352: signal is true;
	signal G6353: std_logic; attribute dont_touch of G6353: signal is true;
	signal G6354: std_logic; attribute dont_touch of G6354: signal is true;
	signal G6355: std_logic; attribute dont_touch of G6355: signal is true;
	signal G6358: std_logic; attribute dont_touch of G6358: signal is true;
	signal G6359: std_logic; attribute dont_touch of G6359: signal is true;
	signal G6360: std_logic; attribute dont_touch of G6360: signal is true;
	signal G6361: std_logic; attribute dont_touch of G6361: signal is true;
	signal G6362: std_logic; attribute dont_touch of G6362: signal is true;
	signal G6363: std_logic; attribute dont_touch of G6363: signal is true;
	signal G6364: std_logic; attribute dont_touch of G6364: signal is true;
	signal G6365: std_logic; attribute dont_touch of G6365: signal is true;
	signal G6368: std_logic; attribute dont_touch of G6368: signal is true;
	signal G6382: std_logic; attribute dont_touch of G6382: signal is true;
	signal G6385: std_logic; attribute dont_touch of G6385: signal is true;
	signal G6386: std_logic; attribute dont_touch of G6386: signal is true;
	signal G6387: std_logic; attribute dont_touch of G6387: signal is true;
	signal G6388: std_logic; attribute dont_touch of G6388: signal is true;
	signal G6389: std_logic; attribute dont_touch of G6389: signal is true;
	signal G6392: std_logic; attribute dont_touch of G6392: signal is true;
	signal G6395: std_logic; attribute dont_touch of G6395: signal is true;
	signal G6396: std_logic; attribute dont_touch of G6396: signal is true;
	signal G6397: std_logic; attribute dont_touch of G6397: signal is true;
	signal G6398: std_logic; attribute dont_touch of G6398: signal is true;
	signal G6399: std_logic; attribute dont_touch of G6399: signal is true;
	signal G6400: std_logic; attribute dont_touch of G6400: signal is true;
	signal G6403: std_logic; attribute dont_touch of G6403: signal is true;
	signal G6404: std_logic; attribute dont_touch of G6404: signal is true;
	signal G6405: std_logic; attribute dont_touch of G6405: signal is true;
	signal G6406: std_logic; attribute dont_touch of G6406: signal is true;
	signal G6407: std_logic; attribute dont_touch of G6407: signal is true;
	signal G6410: std_logic; attribute dont_touch of G6410: signal is true;
	signal G6411: std_logic; attribute dont_touch of G6411: signal is true;
	signal G6412: std_logic; attribute dont_touch of G6412: signal is true;
	signal G6413: std_logic; attribute dont_touch of G6413: signal is true;
	signal G6416: std_logic; attribute dont_touch of G6416: signal is true;
	signal G6417: std_logic; attribute dont_touch of G6417: signal is true;
	signal G6418: std_logic; attribute dont_touch of G6418: signal is true;
	signal G6419: std_logic; attribute dont_touch of G6419: signal is true;
	signal G6420: std_logic; attribute dont_touch of G6420: signal is true;
	signal G6423: std_logic; attribute dont_touch of G6423: signal is true;
	signal G6424: std_logic; attribute dont_touch of G6424: signal is true;
	signal G6425: std_logic; attribute dont_touch of G6425: signal is true;
	signal G6426: std_logic; attribute dont_touch of G6426: signal is true;
	signal G6427: std_logic; attribute dont_touch of G6427: signal is true;
	signal G6430: std_logic; attribute dont_touch of G6430: signal is true;
	signal G6431: std_logic; attribute dont_touch of G6431: signal is true;
	signal G6432: std_logic; attribute dont_touch of G6432: signal is true;
	signal G6433: std_logic; attribute dont_touch of G6433: signal is true;
	signal G6434: std_logic; attribute dont_touch of G6434: signal is true;
	signal G6435: std_logic; attribute dont_touch of G6435: signal is true;
	signal G6438: std_logic; attribute dont_touch of G6438: signal is true;
	signal G6439: std_logic; attribute dont_touch of G6439: signal is true;
	signal G6440: std_logic; attribute dont_touch of G6440: signal is true;
	signal G6441: std_logic; attribute dont_touch of G6441: signal is true;
	signal G6442: std_logic; attribute dont_touch of G6442: signal is true;
	signal G6443: std_logic; attribute dont_touch of G6443: signal is true;
	signal G6444: std_logic; attribute dont_touch of G6444: signal is true;
	signal G6445: std_logic; attribute dont_touch of G6445: signal is true;
	signal G6446: std_logic; attribute dont_touch of G6446: signal is true;
	signal G6447: std_logic; attribute dont_touch of G6447: signal is true;
	signal G6448: std_logic; attribute dont_touch of G6448: signal is true;
	signal G6449: std_logic; attribute dont_touch of G6449: signal is true;
	signal G6450: std_logic; attribute dont_touch of G6450: signal is true;
	signal G6451: std_logic; attribute dont_touch of G6451: signal is true;
	signal G6452: std_logic; attribute dont_touch of G6452: signal is true;
	signal G6453: std_logic; attribute dont_touch of G6453: signal is true;
	signal G6454: std_logic; attribute dont_touch of G6454: signal is true;
	signal G6461: std_logic; attribute dont_touch of G6461: signal is true;
	signal G6462: std_logic; attribute dont_touch of G6462: signal is true;
	signal G6463: std_logic; attribute dont_touch of G6463: signal is true;
	signal G6464: std_logic; attribute dont_touch of G6464: signal is true;
	signal G6465: std_logic; attribute dont_touch of G6465: signal is true;
	signal G6468: std_logic; attribute dont_touch of G6468: signal is true;
	signal G6469: std_logic; attribute dont_touch of G6469: signal is true;
	signal G6470: std_logic; attribute dont_touch of G6470: signal is true;
	signal G6471: std_logic; attribute dont_touch of G6471: signal is true;
	signal G6472: std_logic; attribute dont_touch of G6472: signal is true;
	signal G6475: std_logic; attribute dont_touch of G6475: signal is true;
	signal G6478: std_logic; attribute dont_touch of G6478: signal is true;
	signal G6479: std_logic; attribute dont_touch of G6479: signal is true;
	signal G6480: std_logic; attribute dont_touch of G6480: signal is true;
	signal G6481: std_logic; attribute dont_touch of G6481: signal is true;
	signal G6482: std_logic; attribute dont_touch of G6482: signal is true;
	signal G6485: std_logic; attribute dont_touch of G6485: signal is true;
	signal G6488: std_logic; attribute dont_touch of G6488: signal is true;
	signal G6499: std_logic; attribute dont_touch of G6499: signal is true;
	signal G6500: std_logic; attribute dont_touch of G6500: signal is true;
	signal G6501: std_logic; attribute dont_touch of G6501: signal is true;
	signal G6502: std_logic; attribute dont_touch of G6502: signal is true;
	signal G6503: std_logic; attribute dont_touch of G6503: signal is true;
	signal G6506: std_logic; attribute dont_touch of G6506: signal is true;
	signal G6507: std_logic; attribute dont_touch of G6507: signal is true;
	signal G6508: std_logic; attribute dont_touch of G6508: signal is true;
	signal G6509: std_logic; attribute dont_touch of G6509: signal is true;
	signal G6513: std_logic; attribute dont_touch of G6513: signal is true;
	signal G6514: std_logic; attribute dont_touch of G6514: signal is true;
	signal G6515: std_logic; attribute dont_touch of G6515: signal is true;
	signal G6516: std_logic; attribute dont_touch of G6516: signal is true;
	signal G6517: std_logic; attribute dont_touch of G6517: signal is true;
	signal G6521: std_logic; attribute dont_touch of G6521: signal is true;
	signal G6522: std_logic; attribute dont_touch of G6522: signal is true;
	signal G6523: std_logic; attribute dont_touch of G6523: signal is true;
	signal G6524: std_logic; attribute dont_touch of G6524: signal is true;
	signal G6525: std_logic; attribute dont_touch of G6525: signal is true;
	signal G6526: std_logic; attribute dont_touch of G6526: signal is true;
	signal G6527: std_logic; attribute dont_touch of G6527: signal is true;
	signal G6528: std_logic; attribute dont_touch of G6528: signal is true;
	signal G6529: std_logic; attribute dont_touch of G6529: signal is true;
	signal G6530: std_logic; attribute dont_touch of G6530: signal is true;
	signal G6531: std_logic; attribute dont_touch of G6531: signal is true;
	signal G6532: std_logic; attribute dont_touch of G6532: signal is true;
	signal G6533: std_logic; attribute dont_touch of G6533: signal is true;
	signal G6534: std_logic; attribute dont_touch of G6534: signal is true;
	signal G6535: std_logic; attribute dont_touch of G6535: signal is true;
	signal G6536: std_logic; attribute dont_touch of G6536: signal is true;
	signal G6537: std_logic; attribute dont_touch of G6537: signal is true;
	signal G6538: std_logic; attribute dont_touch of G6538: signal is true;
	signal G6539: std_logic; attribute dont_touch of G6539: signal is true;
	signal G6540: std_logic; attribute dont_touch of G6540: signal is true;
	signal G6541: std_logic; attribute dont_touch of G6541: signal is true;
	signal G6542: std_logic; attribute dont_touch of G6542: signal is true;
	signal G6543: std_logic; attribute dont_touch of G6543: signal is true;
	signal G6544: std_logic; attribute dont_touch of G6544: signal is true;
	signal G6545: std_logic; attribute dont_touch of G6545: signal is true;
	signal G6546: std_logic; attribute dont_touch of G6546: signal is true;
	signal G6547: std_logic; attribute dont_touch of G6547: signal is true;
	signal G6548: std_logic; attribute dont_touch of G6548: signal is true;
	signal G6549: std_logic; attribute dont_touch of G6549: signal is true;
	signal G6550: std_logic; attribute dont_touch of G6550: signal is true;
	signal G6551: std_logic; attribute dont_touch of G6551: signal is true;
	signal G6552: std_logic; attribute dont_touch of G6552: signal is true;
	signal G6553: std_logic; attribute dont_touch of G6553: signal is true;
	signal G6554: std_logic; attribute dont_touch of G6554: signal is true;
	signal G6555: std_logic; attribute dont_touch of G6555: signal is true;
	signal G6556: std_logic; attribute dont_touch of G6556: signal is true;
	signal G6557: std_logic; attribute dont_touch of G6557: signal is true;
	signal G6558: std_logic; attribute dont_touch of G6558: signal is true;
	signal G6559: std_logic; attribute dont_touch of G6559: signal is true;
	signal G6560: std_logic; attribute dont_touch of G6560: signal is true;
	signal G6561: std_logic; attribute dont_touch of G6561: signal is true;
	signal G6562: std_logic; attribute dont_touch of G6562: signal is true;
	signal G6563: std_logic; attribute dont_touch of G6563: signal is true;
	signal G6564: std_logic; attribute dont_touch of G6564: signal is true;
	signal G6565: std_logic; attribute dont_touch of G6565: signal is true;
	signal G6566: std_logic; attribute dont_touch of G6566: signal is true;
	signal G6567: std_logic; attribute dont_touch of G6567: signal is true;
	signal G6568: std_logic; attribute dont_touch of G6568: signal is true;
	signal G6569: std_logic; attribute dont_touch of G6569: signal is true;
	signal G6570: std_logic; attribute dont_touch of G6570: signal is true;
	signal G6571: std_logic; attribute dont_touch of G6571: signal is true;
	signal G6572: std_logic; attribute dont_touch of G6572: signal is true;
	signal G6573: std_logic; attribute dont_touch of G6573: signal is true;
	signal G6574: std_logic; attribute dont_touch of G6574: signal is true;
	signal G6575: std_logic; attribute dont_touch of G6575: signal is true;
	signal G6576: std_logic; attribute dont_touch of G6576: signal is true;
	signal G6577: std_logic; attribute dont_touch of G6577: signal is true;
	signal G6578: std_logic; attribute dont_touch of G6578: signal is true;
	signal G6579: std_logic; attribute dont_touch of G6579: signal is true;
	signal G6580: std_logic; attribute dont_touch of G6580: signal is true;
	signal G6581: std_logic; attribute dont_touch of G6581: signal is true;
	signal G6582: std_logic; attribute dont_touch of G6582: signal is true;
	signal G6583: std_logic; attribute dont_touch of G6583: signal is true;
	signal G6584: std_logic; attribute dont_touch of G6584: signal is true;
	signal G6585: std_logic; attribute dont_touch of G6585: signal is true;
	signal G6586: std_logic; attribute dont_touch of G6586: signal is true;
	signal G6587: std_logic; attribute dont_touch of G6587: signal is true;
	signal G6588: std_logic; attribute dont_touch of G6588: signal is true;
	signal G6589: std_logic; attribute dont_touch of G6589: signal is true;
	signal G6590: std_logic; attribute dont_touch of G6590: signal is true;
	signal G6591: std_logic; attribute dont_touch of G6591: signal is true;
	signal G6592: std_logic; attribute dont_touch of G6592: signal is true;
	signal G6593: std_logic; attribute dont_touch of G6593: signal is true;
	signal G6594: std_logic; attribute dont_touch of G6594: signal is true;
	signal G6595: std_logic; attribute dont_touch of G6595: signal is true;
	signal G6596: std_logic; attribute dont_touch of G6596: signal is true;
	signal G6616: std_logic; attribute dont_touch of G6616: signal is true;
	signal G6617: std_logic; attribute dont_touch of G6617: signal is true;
	signal G6618: std_logic; attribute dont_touch of G6618: signal is true;
	signal G6619: std_logic; attribute dont_touch of G6619: signal is true;
	signal G6620: std_logic; attribute dont_touch of G6620: signal is true;
	signal G6621: std_logic; attribute dont_touch of G6621: signal is true;
	signal G6622: std_logic; attribute dont_touch of G6622: signal is true;
	signal G6623: std_logic; attribute dont_touch of G6623: signal is true;
	signal G6624: std_logic; attribute dont_touch of G6624: signal is true;
	signal G6625: std_logic; attribute dont_touch of G6625: signal is true;
	signal G6626: std_logic; attribute dont_touch of G6626: signal is true;
	signal G6627: std_logic; attribute dont_touch of G6627: signal is true;
	signal G6628: std_logic; attribute dont_touch of G6628: signal is true;
	signal G6629: std_logic; attribute dont_touch of G6629: signal is true;
	signal G6632: std_logic; attribute dont_touch of G6632: signal is true;
	signal G6633: std_logic; attribute dont_touch of G6633: signal is true;
	signal G6634: std_logic; attribute dont_touch of G6634: signal is true;
	signal G6635: std_logic; attribute dont_touch of G6635: signal is true;
	signal G6638: std_logic; attribute dont_touch of G6638: signal is true;
	signal G6639: std_logic; attribute dont_touch of G6639: signal is true;
	signal G6640: std_logic; attribute dont_touch of G6640: signal is true;
	signal G6641: std_logic; attribute dont_touch of G6641: signal is true;
	signal G6644: std_logic; attribute dont_touch of G6644: signal is true;
	signal G6645: std_logic; attribute dont_touch of G6645: signal is true;
	signal G6646: std_logic; attribute dont_touch of G6646: signal is true;
	signal G6647: std_logic; attribute dont_touch of G6647: signal is true;
	signal G6648: std_logic; attribute dont_touch of G6648: signal is true;
	signal G6649: std_logic; attribute dont_touch of G6649: signal is true;
	signal G6652: std_logic; attribute dont_touch of G6652: signal is true;
	signal G6653: std_logic; attribute dont_touch of G6653: signal is true;
	signal G6654: std_logic; attribute dont_touch of G6654: signal is true;
	signal G6655: std_logic; attribute dont_touch of G6655: signal is true;
	signal G6656: std_logic; attribute dont_touch of G6656: signal is true;
	signal G6657: std_logic; attribute dont_touch of G6657: signal is true;
	signal G6660: std_logic; attribute dont_touch of G6660: signal is true;
	signal G6661: std_logic; attribute dont_touch of G6661: signal is true;
	signal G6662: std_logic; attribute dont_touch of G6662: signal is true;
	signal G6663: std_logic; attribute dont_touch of G6663: signal is true;
	signal G6666: std_logic; attribute dont_touch of G6666: signal is true;
	signal G6667: std_logic; attribute dont_touch of G6667: signal is true;
	signal G6670: std_logic; attribute dont_touch of G6670: signal is true;
	signal G6671: std_logic; attribute dont_touch of G6671: signal is true;
	signal G6672: std_logic; attribute dont_touch of G6672: signal is true;
	signal G6673: std_logic; attribute dont_touch of G6673: signal is true;
	signal G6674: std_logic; attribute dont_touch of G6674: signal is true;
	signal G6679: std_logic; attribute dont_touch of G6679: signal is true;
	signal G6680: std_logic; attribute dont_touch of G6680: signal is true;
	signal G6681: std_logic; attribute dont_touch of G6681: signal is true;
	signal G6684: std_logic; attribute dont_touch of G6684: signal is true;
	signal G6685: std_logic; attribute dont_touch of G6685: signal is true;
	signal G6686: std_logic; attribute dont_touch of G6686: signal is true;
	signal G6687: std_logic; attribute dont_touch of G6687: signal is true;
	signal G6688: std_logic; attribute dont_touch of G6688: signal is true;
	signal G6689: std_logic; attribute dont_touch of G6689: signal is true;
	signal G6692: std_logic; attribute dont_touch of G6692: signal is true;
	signal G6693: std_logic; attribute dont_touch of G6693: signal is true;
	signal G6694: std_logic; attribute dont_touch of G6694: signal is true;
	signal G6695: std_logic; attribute dont_touch of G6695: signal is true;
	signal G6696: std_logic; attribute dont_touch of G6696: signal is true;
	signal G6697: std_logic; attribute dont_touch of G6697: signal is true;
	signal G6698: std_logic; attribute dont_touch of G6698: signal is true;
	signal G6699: std_logic; attribute dont_touch of G6699: signal is true;
	signal G6700: std_logic; attribute dont_touch of G6700: signal is true;
	signal G6701: std_logic; attribute dont_touch of G6701: signal is true;
	signal G6702: std_logic; attribute dont_touch of G6702: signal is true;
	signal G6703: std_logic; attribute dont_touch of G6703: signal is true;
	signal G6704: std_logic; attribute dont_touch of G6704: signal is true;
	signal G6705: std_logic; attribute dont_touch of G6705: signal is true;
	signal G6706: std_logic; attribute dont_touch of G6706: signal is true;
	signal G6707: std_logic; attribute dont_touch of G6707: signal is true;
	signal G6708: std_logic; attribute dont_touch of G6708: signal is true;
	signal G6709: std_logic; attribute dont_touch of G6709: signal is true;
	signal G6710: std_logic; attribute dont_touch of G6710: signal is true;
	signal G6711: std_logic; attribute dont_touch of G6711: signal is true;
	signal G6712: std_logic; attribute dont_touch of G6712: signal is true;
	signal G6713: std_logic; attribute dont_touch of G6713: signal is true;
	signal G6714: std_logic; attribute dont_touch of G6714: signal is true;
	signal G6715: std_logic; attribute dont_touch of G6715: signal is true;
	signal G6716: std_logic; attribute dont_touch of G6716: signal is true;
	signal G6717: std_logic; attribute dont_touch of G6717: signal is true;
	signal G6718: std_logic; attribute dont_touch of G6718: signal is true;
	signal G6719: std_logic; attribute dont_touch of G6719: signal is true;
	signal G6720: std_logic; attribute dont_touch of G6720: signal is true;
	signal G6723: std_logic; attribute dont_touch of G6723: signal is true;
	signal G6724: std_logic; attribute dont_touch of G6724: signal is true;
	signal G6727: std_logic; attribute dont_touch of G6727: signal is true;
	signal G6728: std_logic; attribute dont_touch of G6728: signal is true;
	signal G6729: std_logic; attribute dont_touch of G6729: signal is true;
	signal G6730: std_logic; attribute dont_touch of G6730: signal is true;
	signal G6731: std_logic; attribute dont_touch of G6731: signal is true;
	signal G6732: std_logic; attribute dont_touch of G6732: signal is true;
	signal G6733: std_logic; attribute dont_touch of G6733: signal is true;
	signal G6734: std_logic; attribute dont_touch of G6734: signal is true;
	signal G6735: std_logic; attribute dont_touch of G6735: signal is true;
	signal G6736: std_logic; attribute dont_touch of G6736: signal is true;
	signal G6737: std_logic; attribute dont_touch of G6737: signal is true;
	signal G6738: std_logic; attribute dont_touch of G6738: signal is true;
	signal G6739: std_logic; attribute dont_touch of G6739: signal is true;
	signal G6740: std_logic; attribute dont_touch of G6740: signal is true;
	signal G6741: std_logic; attribute dont_touch of G6741: signal is true;
	signal G6742: std_logic; attribute dont_touch of G6742: signal is true;
	signal G6743: std_logic; attribute dont_touch of G6743: signal is true;
	signal G6744: std_logic; attribute dont_touch of G6744: signal is true;
	signal G6745: std_logic; attribute dont_touch of G6745: signal is true;
	signal G6746: std_logic; attribute dont_touch of G6746: signal is true;
	signal G6747: std_logic; attribute dont_touch of G6747: signal is true;
	signal G6748: std_logic; attribute dont_touch of G6748: signal is true;
	signal G6749: std_logic; attribute dont_touch of G6749: signal is true;
	signal G6750: std_logic; attribute dont_touch of G6750: signal is true;
	signal G6751: std_logic; attribute dont_touch of G6751: signal is true;
	signal G6752: std_logic; attribute dont_touch of G6752: signal is true;
	signal G6755: std_logic; attribute dont_touch of G6755: signal is true;
	signal G6756: std_logic; attribute dont_touch of G6756: signal is true;
	signal G6757: std_logic; attribute dont_touch of G6757: signal is true;
	signal G6758: std_logic; attribute dont_touch of G6758: signal is true;
	signal G6759: std_logic; attribute dont_touch of G6759: signal is true;
	signal G6760: std_logic; attribute dont_touch of G6760: signal is true;
	signal G6763: std_logic; attribute dont_touch of G6763: signal is true;
	signal G6764: std_logic; attribute dont_touch of G6764: signal is true;
	signal G6771: std_logic; attribute dont_touch of G6771: signal is true;
	signal G6772: std_logic; attribute dont_touch of G6772: signal is true;
	signal G6775: std_logic; attribute dont_touch of G6775: signal is true;
	signal G6776: std_logic; attribute dont_touch of G6776: signal is true;
	signal G6777: std_logic; attribute dont_touch of G6777: signal is true;
	signal G6778: std_logic; attribute dont_touch of G6778: signal is true;
	signal G6786: std_logic; attribute dont_touch of G6786: signal is true;
	signal G6787: std_logic; attribute dont_touch of G6787: signal is true;
	signal G6788: std_logic; attribute dont_touch of G6788: signal is true;
	signal G6789: std_logic; attribute dont_touch of G6789: signal is true;
	signal G6790: std_logic; attribute dont_touch of G6790: signal is true;
	signal G6791: std_logic; attribute dont_touch of G6791: signal is true;
	signal G6792: std_logic; attribute dont_touch of G6792: signal is true;
	signal G6793: std_logic; attribute dont_touch of G6793: signal is true;
	signal G6794: std_logic; attribute dont_touch of G6794: signal is true;
	signal G6795: std_logic; attribute dont_touch of G6795: signal is true;
	signal G6796: std_logic; attribute dont_touch of G6796: signal is true;
	signal G6797: std_logic; attribute dont_touch of G6797: signal is true;
	signal G6798: std_logic; attribute dont_touch of G6798: signal is true;
	signal G6799: std_logic; attribute dont_touch of G6799: signal is true;
	signal G6800: std_logic; attribute dont_touch of G6800: signal is true;
	signal G6801: std_logic; attribute dont_touch of G6801: signal is true;
	signal G6802: std_logic; attribute dont_touch of G6802: signal is true;
	signal G6803: std_logic; attribute dont_touch of G6803: signal is true;
	signal G6804: std_logic; attribute dont_touch of G6804: signal is true;
	signal G6805: std_logic; attribute dont_touch of G6805: signal is true;
	signal G6806: std_logic; attribute dont_touch of G6806: signal is true;
	signal G6807: std_logic; attribute dont_touch of G6807: signal is true;
	signal G6808: std_logic; attribute dont_touch of G6808: signal is true;
	signal G6809: std_logic; attribute dont_touch of G6809: signal is true;
	signal G6810: std_logic; attribute dont_touch of G6810: signal is true;
	signal G6811: std_logic; attribute dont_touch of G6811: signal is true;
	signal G6812: std_logic; attribute dont_touch of G6812: signal is true;
	signal G6813: std_logic; attribute dont_touch of G6813: signal is true;
	signal G6814: std_logic; attribute dont_touch of G6814: signal is true;
	signal G6815: std_logic; attribute dont_touch of G6815: signal is true;
	signal G6816: std_logic; attribute dont_touch of G6816: signal is true;
	signal G6817: std_logic; attribute dont_touch of G6817: signal is true;
	signal G6818: std_logic; attribute dont_touch of G6818: signal is true;
	signal G6819: std_logic; attribute dont_touch of G6819: signal is true;
	signal G6820: std_logic; attribute dont_touch of G6820: signal is true;
	signal G6821: std_logic; attribute dont_touch of G6821: signal is true;
	signal G6822: std_logic; attribute dont_touch of G6822: signal is true;
	signal G6823: std_logic; attribute dont_touch of G6823: signal is true;
	signal G6824: std_logic; attribute dont_touch of G6824: signal is true;
	signal G6825: std_logic; attribute dont_touch of G6825: signal is true;
	signal G6826: std_logic; attribute dont_touch of G6826: signal is true;
	signal G6827: std_logic; attribute dont_touch of G6827: signal is true;
	signal G6828: std_logic; attribute dont_touch of G6828: signal is true;
	signal G6829: std_logic; attribute dont_touch of G6829: signal is true;
	signal G6830: std_logic; attribute dont_touch of G6830: signal is true;
	signal G6831: std_logic; attribute dont_touch of G6831: signal is true;
	signal G6832: std_logic; attribute dont_touch of G6832: signal is true;
	signal G6833: std_logic; attribute dont_touch of G6833: signal is true;
	signal G6834: std_logic; attribute dont_touch of G6834: signal is true;
	signal G6835: std_logic; attribute dont_touch of G6835: signal is true;
	signal G6836: std_logic; attribute dont_touch of G6836: signal is true;
	signal G6837: std_logic; attribute dont_touch of G6837: signal is true;
	signal G6838: std_logic; attribute dont_touch of G6838: signal is true;
	signal G6839: std_logic; attribute dont_touch of G6839: signal is true;
	signal G6840: std_logic; attribute dont_touch of G6840: signal is true;
	signal G6841: std_logic; attribute dont_touch of G6841: signal is true;
	signal G6843: std_logic; attribute dont_touch of G6843: signal is true;
	signal G6844: std_logic; attribute dont_touch of G6844: signal is true;
	signal G6845: std_logic; attribute dont_touch of G6845: signal is true;
	signal G6846: std_logic; attribute dont_touch of G6846: signal is true;
	signal G6847: std_logic; attribute dont_touch of G6847: signal is true;
	signal G6852: std_logic; attribute dont_touch of G6852: signal is true;
	signal G6853: std_logic; attribute dont_touch of G6853: signal is true;
	signal G6854: std_logic; attribute dont_touch of G6854: signal is true;
	signal G6855: std_logic; attribute dont_touch of G6855: signal is true;
	signal G6856: std_logic; attribute dont_touch of G6856: signal is true;
	signal G6857: std_logic; attribute dont_touch of G6857: signal is true;
	signal G6858: std_logic; attribute dont_touch of G6858: signal is true;
	signal G6859: std_logic; attribute dont_touch of G6859: signal is true;
	signal G6860: std_logic; attribute dont_touch of G6860: signal is true;
	signal G6861: std_logic; attribute dont_touch of G6861: signal is true;
	signal G6862: std_logic; attribute dont_touch of G6862: signal is true;
	signal G6863: std_logic; attribute dont_touch of G6863: signal is true;
	signal G6868: std_logic; attribute dont_touch of G6868: signal is true;
	signal G6869: std_logic; attribute dont_touch of G6869: signal is true;
	signal G6870: std_logic; attribute dont_touch of G6870: signal is true;
	signal G6871: std_logic; attribute dont_touch of G6871: signal is true;
	signal G6872: std_logic; attribute dont_touch of G6872: signal is true;
	signal G6873: std_logic; attribute dont_touch of G6873: signal is true;
	signal G6874: std_logic; attribute dont_touch of G6874: signal is true;
	signal G6875: std_logic; attribute dont_touch of G6875: signal is true;
	signal G6876: std_logic; attribute dont_touch of G6876: signal is true;
	signal G6877: std_logic; attribute dont_touch of G6877: signal is true;
	signal G6878: std_logic; attribute dont_touch of G6878: signal is true;
	signal G6879: std_logic; attribute dont_touch of G6879: signal is true;
	signal G6880: std_logic; attribute dont_touch of G6880: signal is true;
	signal G6881: std_logic; attribute dont_touch of G6881: signal is true;
	signal G6882: std_logic; attribute dont_touch of G6882: signal is true;
	signal G6883: std_logic; attribute dont_touch of G6883: signal is true;
	signal G6884: std_logic; attribute dont_touch of G6884: signal is true;
	signal G6885: std_logic; attribute dont_touch of G6885: signal is true;
	signal G6886: std_logic; attribute dont_touch of G6886: signal is true;
	signal G6887: std_logic; attribute dont_touch of G6887: signal is true;
	signal G6888: std_logic; attribute dont_touch of G6888: signal is true;
	signal G6889: std_logic; attribute dont_touch of G6889: signal is true;
	signal G6890: std_logic; attribute dont_touch of G6890: signal is true;
	signal G6891: std_logic; attribute dont_touch of G6891: signal is true;
	signal G6892: std_logic; attribute dont_touch of G6892: signal is true;
	signal G6893: std_logic; attribute dont_touch of G6893: signal is true;
	signal G6894: std_logic; attribute dont_touch of G6894: signal is true;
	signal G6895: std_logic; attribute dont_touch of G6895: signal is true;
	signal G6896: std_logic; attribute dont_touch of G6896: signal is true;
	signal G6897: std_logic; attribute dont_touch of G6897: signal is true;
	signal G6898: std_logic; attribute dont_touch of G6898: signal is true;
	signal G6899: std_logic; attribute dont_touch of G6899: signal is true;
	signal G6900: std_logic; attribute dont_touch of G6900: signal is true;
	signal G6901: std_logic; attribute dont_touch of G6901: signal is true;
	signal G6902: std_logic; attribute dont_touch of G6902: signal is true;
	signal G6903: std_logic; attribute dont_touch of G6903: signal is true;
	signal G6904: std_logic; attribute dont_touch of G6904: signal is true;
	signal G6905: std_logic; attribute dont_touch of G6905: signal is true;
	signal G6906: std_logic; attribute dont_touch of G6906: signal is true;
	signal G6907: std_logic; attribute dont_touch of G6907: signal is true;
	signal G6908: std_logic; attribute dont_touch of G6908: signal is true;
	signal G6909: std_logic; attribute dont_touch of G6909: signal is true;
	signal G6910: std_logic; attribute dont_touch of G6910: signal is true;
	signal G6911: std_logic; attribute dont_touch of G6911: signal is true;
	signal G6912: std_logic; attribute dont_touch of G6912: signal is true;
	signal G6913: std_logic; attribute dont_touch of G6913: signal is true;
	signal G6914: std_logic; attribute dont_touch of G6914: signal is true;
	signal G6915: std_logic; attribute dont_touch of G6915: signal is true;
	signal G6916: std_logic; attribute dont_touch of G6916: signal is true;
	signal G6917: std_logic; attribute dont_touch of G6917: signal is true;
	signal G6918: std_logic; attribute dont_touch of G6918: signal is true;
	signal G6919: std_logic; attribute dont_touch of G6919: signal is true;
	signal G6921: std_logic; attribute dont_touch of G6921: signal is true;
	signal G6922: std_logic; attribute dont_touch of G6922: signal is true;
	signal G6923: std_logic; attribute dont_touch of G6923: signal is true;
	signal G6924: std_logic; attribute dont_touch of G6924: signal is true;
	signal G6925: std_logic; attribute dont_touch of G6925: signal is true;
	signal G6927: std_logic; attribute dont_touch of G6927: signal is true;
	signal G6928: std_logic; attribute dont_touch of G6928: signal is true;
	signal G6929: std_logic; attribute dont_touch of G6929: signal is true;
	signal G6930: std_logic; attribute dont_touch of G6930: signal is true;
	signal G6931: std_logic; attribute dont_touch of G6931: signal is true;
	signal G6933: std_logic; attribute dont_touch of G6933: signal is true;
	signal G6934: std_logic; attribute dont_touch of G6934: signal is true;
	signal G6935: std_logic; attribute dont_touch of G6935: signal is true;
	signal G6938: std_logic; attribute dont_touch of G6938: signal is true;
	signal G6939: std_logic; attribute dont_touch of G6939: signal is true;
	signal G6940: std_logic; attribute dont_touch of G6940: signal is true;
	signal G6941: std_logic; attribute dont_touch of G6941: signal is true;
	signal G6943: std_logic; attribute dont_touch of G6943: signal is true;
	signal G6944: std_logic; attribute dont_touch of G6944: signal is true;
	signal G6947: std_logic; attribute dont_touch of G6947: signal is true;
	signal G6948: std_logic; attribute dont_touch of G6948: signal is true;
	signal G6950: std_logic; attribute dont_touch of G6950: signal is true;
	signal G6951: std_logic; attribute dont_touch of G6951: signal is true;
	signal G6954: std_logic; attribute dont_touch of G6954: signal is true;
	signal G6956: std_logic; attribute dont_touch of G6956: signal is true;
	signal G6957: std_logic; attribute dont_touch of G6957: signal is true;
	signal G6960: std_logic; attribute dont_touch of G6960: signal is true;
	signal G6961: std_logic; attribute dont_touch of G6961: signal is true;
	signal G6964: std_logic; attribute dont_touch of G6964: signal is true;
	signal G6967: std_logic; attribute dont_touch of G6967: signal is true;
	signal G6970: std_logic; attribute dont_touch of G6970: signal is true;
	signal G6971: std_logic; attribute dont_touch of G6971: signal is true;
	signal G6974: std_logic; attribute dont_touch of G6974: signal is true;
	signal G6980: std_logic; attribute dont_touch of G6980: signal is true;
	signal G6983: std_logic; attribute dont_touch of G6983: signal is true;
	signal G6984: std_logic; attribute dont_touch of G6984: signal is true;
	signal G6990: std_logic; attribute dont_touch of G6990: signal is true;
	signal G6993: std_logic; attribute dont_touch of G6993: signal is true;
	signal G6994: std_logic; attribute dont_touch of G6994: signal is true;
	signal G6995: std_logic; attribute dont_touch of G6995: signal is true;
	signal G7001: std_logic; attribute dont_touch of G7001: signal is true;
	signal G7004: std_logic; attribute dont_touch of G7004: signal is true;
	signal G7007: std_logic; attribute dont_touch of G7007: signal is true;
	signal G7008: std_logic; attribute dont_touch of G7008: signal is true;
	signal G7009: std_logic; attribute dont_touch of G7009: signal is true;
	signal G7010: std_logic; attribute dont_touch of G7010: signal is true;
	signal G7011: std_logic; attribute dont_touch of G7011: signal is true;
	signal G7020: std_logic; attribute dont_touch of G7020: signal is true;
	signal G7021: std_logic; attribute dont_touch of G7021: signal is true;
	signal G7022: std_logic; attribute dont_touch of G7022: signal is true;
	signal G7023: std_logic; attribute dont_touch of G7023: signal is true;
	signal G7024: std_logic; attribute dont_touch of G7024: signal is true;
	signal G7025: std_logic; attribute dont_touch of G7025: signal is true;
	signal G7026: std_logic; attribute dont_touch of G7026: signal is true;
	signal G7027: std_logic; attribute dont_touch of G7027: signal is true;
	signal G7028: std_logic; attribute dont_touch of G7028: signal is true;
	signal G7029: std_logic; attribute dont_touch of G7029: signal is true;
	signal G7030: std_logic; attribute dont_touch of G7030: signal is true;
	signal G7031: std_logic; attribute dont_touch of G7031: signal is true;
	signal G7032: std_logic; attribute dont_touch of G7032: signal is true;
	signal G7033: std_logic; attribute dont_touch of G7033: signal is true;
	signal G7034: std_logic; attribute dont_touch of G7034: signal is true;
	signal G7035: std_logic; attribute dont_touch of G7035: signal is true;
	signal G7036: std_logic; attribute dont_touch of G7036: signal is true;
	signal G7037: std_logic; attribute dont_touch of G7037: signal is true;
	signal G7038: std_logic; attribute dont_touch of G7038: signal is true;
	signal G7039: std_logic; attribute dont_touch of G7039: signal is true;
	signal G7040: std_logic; attribute dont_touch of G7040: signal is true;
	signal G7041: std_logic; attribute dont_touch of G7041: signal is true;
	signal G7042: std_logic; attribute dont_touch of G7042: signal is true;
	signal G7043: std_logic; attribute dont_touch of G7043: signal is true;
	signal G7044: std_logic; attribute dont_touch of G7044: signal is true;
	signal G7045: std_logic; attribute dont_touch of G7045: signal is true;
	signal G7046: std_logic; attribute dont_touch of G7046: signal is true;
	signal G7047: std_logic; attribute dont_touch of G7047: signal is true;
	signal G7048: std_logic; attribute dont_touch of G7048: signal is true;
	signal G7049: std_logic; attribute dont_touch of G7049: signal is true;
	signal G7050: std_logic; attribute dont_touch of G7050: signal is true;
	signal G7051: std_logic; attribute dont_touch of G7051: signal is true;
	signal G7052: std_logic; attribute dont_touch of G7052: signal is true;
	signal G7053: std_logic; attribute dont_touch of G7053: signal is true;
	signal G7054: std_logic; attribute dont_touch of G7054: signal is true;
	signal G7055: std_logic; attribute dont_touch of G7055: signal is true;
	signal G7056: std_logic; attribute dont_touch of G7056: signal is true;
	signal G7057: std_logic; attribute dont_touch of G7057: signal is true;
	signal G7058: std_logic; attribute dont_touch of G7058: signal is true;
	signal G7059: std_logic; attribute dont_touch of G7059: signal is true;
	signal G7060: std_logic; attribute dont_touch of G7060: signal is true;
	signal G7061: std_logic; attribute dont_touch of G7061: signal is true;
	signal G7062: std_logic; attribute dont_touch of G7062: signal is true;
	signal G7063: std_logic; attribute dont_touch of G7063: signal is true;
	signal G7064: std_logic; attribute dont_touch of G7064: signal is true;
	signal G7065: std_logic; attribute dont_touch of G7065: signal is true;
	signal G7066: std_logic; attribute dont_touch of G7066: signal is true;
	signal G7067: std_logic; attribute dont_touch of G7067: signal is true;
	signal G7068: std_logic; attribute dont_touch of G7068: signal is true;
	signal G7069: std_logic; attribute dont_touch of G7069: signal is true;
	signal G7070: std_logic; attribute dont_touch of G7070: signal is true;
	signal G7071: std_logic; attribute dont_touch of G7071: signal is true;
	signal G7072: std_logic; attribute dont_touch of G7072: signal is true;
	signal G7073: std_logic; attribute dont_touch of G7073: signal is true;
	signal G7074: std_logic; attribute dont_touch of G7074: signal is true;
	signal G7075: std_logic; attribute dont_touch of G7075: signal is true;
	signal G7076: std_logic; attribute dont_touch of G7076: signal is true;
	signal G7077: std_logic; attribute dont_touch of G7077: signal is true;
	signal G7078: std_logic; attribute dont_touch of G7078: signal is true;
	signal G7079: std_logic; attribute dont_touch of G7079: signal is true;
	signal G7082: std_logic; attribute dont_touch of G7082: signal is true;
	signal G7085: std_logic; attribute dont_touch of G7085: signal is true;
	signal G7088: std_logic; attribute dont_touch of G7088: signal is true;
	signal G7089: std_logic; attribute dont_touch of G7089: signal is true;
	signal G7092: std_logic; attribute dont_touch of G7092: signal is true;
	signal G7093: std_logic; attribute dont_touch of G7093: signal is true;
	signal G7096: std_logic; attribute dont_touch of G7096: signal is true;
	signal G7097: std_logic; attribute dont_touch of G7097: signal is true;
	signal G7098: std_logic; attribute dont_touch of G7098: signal is true;
	signal G7101: std_logic; attribute dont_touch of G7101: signal is true;
	signal G7102: std_logic; attribute dont_touch of G7102: signal is true;
	signal G7103: std_logic; attribute dont_touch of G7103: signal is true;
	signal G7106: std_logic; attribute dont_touch of G7106: signal is true;
	signal G7107: std_logic; attribute dont_touch of G7107: signal is true;
	signal G7110: std_logic; attribute dont_touch of G7110: signal is true;
	signal G7113: std_logic; attribute dont_touch of G7113: signal is true;
	signal G7116: std_logic; attribute dont_touch of G7116: signal is true;
	signal G7119: std_logic; attribute dont_touch of G7119: signal is true;
	signal G7122: std_logic; attribute dont_touch of G7122: signal is true;
	signal G7123: std_logic; attribute dont_touch of G7123: signal is true;
	signal G7124: std_logic; attribute dont_touch of G7124: signal is true;
	signal G7125: std_logic; attribute dont_touch of G7125: signal is true;
	signal G7126: std_logic; attribute dont_touch of G7126: signal is true;
	signal G7127: std_logic; attribute dont_touch of G7127: signal is true;
	signal G7130: std_logic; attribute dont_touch of G7130: signal is true;
	signal G7131: std_logic; attribute dont_touch of G7131: signal is true;
	signal G7132: std_logic; attribute dont_touch of G7132: signal is true;
	signal G7133: std_logic; attribute dont_touch of G7133: signal is true;
	signal G7134: std_logic; attribute dont_touch of G7134: signal is true;
	signal G7135: std_logic; attribute dont_touch of G7135: signal is true;
	signal G7136: std_logic; attribute dont_touch of G7136: signal is true;
	signal G7137: std_logic; attribute dont_touch of G7137: signal is true;
	signal G7138: std_logic; attribute dont_touch of G7138: signal is true;
	signal G7139: std_logic; attribute dont_touch of G7139: signal is true;
	signal G7140: std_logic; attribute dont_touch of G7140: signal is true;
	signal G7141: std_logic; attribute dont_touch of G7141: signal is true;
	signal G7142: std_logic; attribute dont_touch of G7142: signal is true;
	signal G7143: std_logic; attribute dont_touch of G7143: signal is true;
	signal G7144: std_logic; attribute dont_touch of G7144: signal is true;
	signal G7145: std_logic; attribute dont_touch of G7145: signal is true;
	signal G7146: std_logic; attribute dont_touch of G7146: signal is true;
	signal G7147: std_logic; attribute dont_touch of G7147: signal is true;
	signal G7148: std_logic; attribute dont_touch of G7148: signal is true;
	signal G7182: std_logic; attribute dont_touch of G7182: signal is true;
	signal G7183: std_logic; attribute dont_touch of G7183: signal is true;
	signal G7184: std_logic; attribute dont_touch of G7184: signal is true;
	signal G7185: std_logic; attribute dont_touch of G7185: signal is true;
	signal G7186: std_logic; attribute dont_touch of G7186: signal is true;
	signal G7187: std_logic; attribute dont_touch of G7187: signal is true;
	signal G7188: std_logic; attribute dont_touch of G7188: signal is true;
	signal G7189: std_logic; attribute dont_touch of G7189: signal is true;
	signal G7190: std_logic; attribute dont_touch of G7190: signal is true;
	signal G7191: std_logic; attribute dont_touch of G7191: signal is true;
	signal G7192: std_logic; attribute dont_touch of G7192: signal is true;
	signal G7195: std_logic; attribute dont_touch of G7195: signal is true;
	signal G7196: std_logic; attribute dont_touch of G7196: signal is true;
	signal G7197: std_logic; attribute dont_touch of G7197: signal is true;
	signal G7200: std_logic; attribute dont_touch of G7200: signal is true;
	signal G7201: std_logic; attribute dont_touch of G7201: signal is true;
	signal G7202: std_logic; attribute dont_touch of G7202: signal is true;
	signal G7203: std_logic; attribute dont_touch of G7203: signal is true;
	signal G7204: std_logic; attribute dont_touch of G7204: signal is true;
	signal G7205: std_logic; attribute dont_touch of G7205: signal is true;
	signal G7206: std_logic; attribute dont_touch of G7206: signal is true;
	signal G7209: std_logic; attribute dont_touch of G7209: signal is true;
	signal G7210: std_logic; attribute dont_touch of G7210: signal is true;
	signal G7211: std_logic; attribute dont_touch of G7211: signal is true;
	signal G7212: std_logic; attribute dont_touch of G7212: signal is true;
	signal G7213: std_logic; attribute dont_touch of G7213: signal is true;
	signal G7214: std_logic; attribute dont_touch of G7214: signal is true;
	signal G7217: std_logic; attribute dont_touch of G7217: signal is true;
	signal G7218: std_logic; attribute dont_touch of G7218: signal is true;
	signal G7219: std_logic; attribute dont_touch of G7219: signal is true;
	signal G7220: std_logic; attribute dont_touch of G7220: signal is true;
	signal G7221: std_logic; attribute dont_touch of G7221: signal is true;
	signal G7224: std_logic; attribute dont_touch of G7224: signal is true;
	signal G7225: std_logic; attribute dont_touch of G7225: signal is true;
	signal G7226: std_logic; attribute dont_touch of G7226: signal is true;
	signal G7227: std_logic; attribute dont_touch of G7227: signal is true;
	signal G7230: std_logic; attribute dont_touch of G7230: signal is true;
	signal G7231: std_logic; attribute dont_touch of G7231: signal is true;
	signal G7232: std_logic; attribute dont_touch of G7232: signal is true;
	signal G7235: std_logic; attribute dont_touch of G7235: signal is true;
	signal G7236: std_logic; attribute dont_touch of G7236: signal is true;
	signal G7237: std_logic; attribute dont_touch of G7237: signal is true;
	signal G7240: std_logic; attribute dont_touch of G7240: signal is true;
	signal G7241: std_logic; attribute dont_touch of G7241: signal is true;
	signal G7242: std_logic; attribute dont_touch of G7242: signal is true;
	signal G7243: std_logic; attribute dont_touch of G7243: signal is true;
	signal G7244: std_logic; attribute dont_touch of G7244: signal is true;
	signal G7245: std_logic; attribute dont_touch of G7245: signal is true;
	signal G7246: std_logic; attribute dont_touch of G7246: signal is true;
	signal G7256: std_logic; attribute dont_touch of G7256: signal is true;
	signal G7257: std_logic; attribute dont_touch of G7257: signal is true;
	signal G7258: std_logic; attribute dont_touch of G7258: signal is true;
	signal G7259: std_logic; attribute dont_touch of G7259: signal is true;
	signal G7260: std_logic; attribute dont_touch of G7260: signal is true;
	signal G7263: std_logic; attribute dont_touch of G7263: signal is true;
	signal G7264: std_logic; attribute dont_touch of G7264: signal is true;
	signal G7265: std_logic; attribute dont_touch of G7265: signal is true;
	signal G7268: std_logic; attribute dont_touch of G7268: signal is true;
	signal G7269: std_logic; attribute dont_touch of G7269: signal is true;
	signal G7270: std_logic; attribute dont_touch of G7270: signal is true;
	signal G7271: std_logic; attribute dont_touch of G7271: signal is true;
	signal G7272: std_logic; attribute dont_touch of G7272: signal is true;
	signal G7273: std_logic; attribute dont_touch of G7273: signal is true;
	signal G7277: std_logic; attribute dont_touch of G7277: signal is true;
	signal G7278: std_logic; attribute dont_touch of G7278: signal is true;
	signal G7279: std_logic; attribute dont_touch of G7279: signal is true;
	signal G7284: std_logic; attribute dont_touch of G7284: signal is true;
	signal G7285: std_logic; attribute dont_touch of G7285: signal is true;
	signal G7286: std_logic; attribute dont_touch of G7286: signal is true;
	signal G7287: std_logic; attribute dont_touch of G7287: signal is true;
	signal G7288: std_logic; attribute dont_touch of G7288: signal is true;
	signal G7289: std_logic; attribute dont_touch of G7289: signal is true;
	signal G7290: std_logic; attribute dont_touch of G7290: signal is true;
	signal G7291: std_logic; attribute dont_touch of G7291: signal is true;
	signal G7292: std_logic; attribute dont_touch of G7292: signal is true;
	signal G7293: std_logic; attribute dont_touch of G7293: signal is true;
	signal G7294: std_logic; attribute dont_touch of G7294: signal is true;
	signal G7295: std_logic; attribute dont_touch of G7295: signal is true;
	signal G7296: std_logic; attribute dont_touch of G7296: signal is true;
	signal G7297: std_logic; attribute dont_touch of G7297: signal is true;
	signal G7298: std_logic; attribute dont_touch of G7298: signal is true;
	signal G7299: std_logic; attribute dont_touch of G7299: signal is true;
	signal G7300: std_logic; attribute dont_touch of G7300: signal is true;
	signal G7301: std_logic; attribute dont_touch of G7301: signal is true;
	signal G7302: std_logic; attribute dont_touch of G7302: signal is true;
	signal G7303: std_logic; attribute dont_touch of G7303: signal is true;
	signal G7304: std_logic; attribute dont_touch of G7304: signal is true;
	signal G7305: std_logic; attribute dont_touch of G7305: signal is true;
	signal G7306: std_logic; attribute dont_touch of G7306: signal is true;
	signal G7307: std_logic; attribute dont_touch of G7307: signal is true;
	signal G7308: std_logic; attribute dont_touch of G7308: signal is true;
	signal G7309: std_logic; attribute dont_touch of G7309: signal is true;
	signal G7310: std_logic; attribute dont_touch of G7310: signal is true;
	signal G7311: std_logic; attribute dont_touch of G7311: signal is true;
	signal G7312: std_logic; attribute dont_touch of G7312: signal is true;
	signal G7313: std_logic; attribute dont_touch of G7313: signal is true;
	signal G7314: std_logic; attribute dont_touch of G7314: signal is true;
	signal G7315: std_logic; attribute dont_touch of G7315: signal is true;
	signal G7316: std_logic; attribute dont_touch of G7316: signal is true;
	signal G7317: std_logic; attribute dont_touch of G7317: signal is true;
	signal G7318: std_logic; attribute dont_touch of G7318: signal is true;
	signal G7319: std_logic; attribute dont_touch of G7319: signal is true;
	signal G7320: std_logic; attribute dont_touch of G7320: signal is true;
	signal G7321: std_logic; attribute dont_touch of G7321: signal is true;
	signal G7322: std_logic; attribute dont_touch of G7322: signal is true;
	signal G7323: std_logic; attribute dont_touch of G7323: signal is true;
	signal G7324: std_logic; attribute dont_touch of G7324: signal is true;
	signal G7325: std_logic; attribute dont_touch of G7325: signal is true;
	signal G7326: std_logic; attribute dont_touch of G7326: signal is true;
	signal G7327: std_logic; attribute dont_touch of G7327: signal is true;
	signal G7328: std_logic; attribute dont_touch of G7328: signal is true;
	signal G7329: std_logic; attribute dont_touch of G7329: signal is true;
	signal G7330: std_logic; attribute dont_touch of G7330: signal is true;
	signal G7331: std_logic; attribute dont_touch of G7331: signal is true;
	signal G7332: std_logic; attribute dont_touch of G7332: signal is true;
	signal G7333: std_logic; attribute dont_touch of G7333: signal is true;
	signal G7334: std_logic; attribute dont_touch of G7334: signal is true;
	signal G7335: std_logic; attribute dont_touch of G7335: signal is true;
	signal G7336: std_logic; attribute dont_touch of G7336: signal is true;
	signal G7337: std_logic; attribute dont_touch of G7337: signal is true;
	signal G7338: std_logic; attribute dont_touch of G7338: signal is true;
	signal G7339: std_logic; attribute dont_touch of G7339: signal is true;
	signal G7340: std_logic; attribute dont_touch of G7340: signal is true;
	signal G7341: std_logic; attribute dont_touch of G7341: signal is true;
	signal G7342: std_logic; attribute dont_touch of G7342: signal is true;
	signal G7343: std_logic; attribute dont_touch of G7343: signal is true;
	signal G7344: std_logic; attribute dont_touch of G7344: signal is true;
	signal G7345: std_logic; attribute dont_touch of G7345: signal is true;
	signal G7346: std_logic; attribute dont_touch of G7346: signal is true;
	signal G7347: std_logic; attribute dont_touch of G7347: signal is true;
	signal G7348: std_logic; attribute dont_touch of G7348: signal is true;
	signal G7349: std_logic; attribute dont_touch of G7349: signal is true;
	signal G7350: std_logic; attribute dont_touch of G7350: signal is true;
	signal G7351: std_logic; attribute dont_touch of G7351: signal is true;
	signal G7352: std_logic; attribute dont_touch of G7352: signal is true;
	signal G7353: std_logic; attribute dont_touch of G7353: signal is true;
	signal G7354: std_logic; attribute dont_touch of G7354: signal is true;
	signal G7355: std_logic; attribute dont_touch of G7355: signal is true;
	signal G7356: std_logic; attribute dont_touch of G7356: signal is true;
	signal G7357: std_logic; attribute dont_touch of G7357: signal is true;
	signal G7358: std_logic; attribute dont_touch of G7358: signal is true;
	signal G7359: std_logic; attribute dont_touch of G7359: signal is true;
	signal G7360: std_logic; attribute dont_touch of G7360: signal is true;
	signal G7361: std_logic; attribute dont_touch of G7361: signal is true;
	signal G7362: std_logic; attribute dont_touch of G7362: signal is true;
	signal G7363: std_logic; attribute dont_touch of G7363: signal is true;
	signal G7364: std_logic; attribute dont_touch of G7364: signal is true;
	signal G7365: std_logic; attribute dont_touch of G7365: signal is true;
	signal G7366: std_logic; attribute dont_touch of G7366: signal is true;
	signal G7367: std_logic; attribute dont_touch of G7367: signal is true;
	signal G7368: std_logic; attribute dont_touch of G7368: signal is true;
	signal G7369: std_logic; attribute dont_touch of G7369: signal is true;
	signal G7374: std_logic; attribute dont_touch of G7374: signal is true;
	signal G7375: std_logic; attribute dont_touch of G7375: signal is true;
	signal G7376: std_logic; attribute dont_touch of G7376: signal is true;
	signal G7377: std_logic; attribute dont_touch of G7377: signal is true;
	signal G7378: std_logic; attribute dont_touch of G7378: signal is true;
	signal G7379: std_logic; attribute dont_touch of G7379: signal is true;
	signal G7380: std_logic; attribute dont_touch of G7380: signal is true;
	signal G7384: std_logic; attribute dont_touch of G7384: signal is true;
	signal G7385: std_logic; attribute dont_touch of G7385: signal is true;
	signal G7386: std_logic; attribute dont_touch of G7386: signal is true;
	signal G7387: std_logic; attribute dont_touch of G7387: signal is true;
	signal G7388: std_logic; attribute dont_touch of G7388: signal is true;
	signal G7389: std_logic; attribute dont_touch of G7389: signal is true;
	signal G7390: std_logic; attribute dont_touch of G7390: signal is true;
	signal G7394: std_logic; attribute dont_touch of G7394: signal is true;
	signal G7395: std_logic; attribute dont_touch of G7395: signal is true;
	signal G7402: std_logic; attribute dont_touch of G7402: signal is true;
	signal G7403: std_logic; attribute dont_touch of G7403: signal is true;
	signal G7406: std_logic; attribute dont_touch of G7406: signal is true;
	signal G7409: std_logic; attribute dont_touch of G7409: signal is true;
	signal G7410: std_logic; attribute dont_touch of G7410: signal is true;
	signal G7413: std_logic; attribute dont_touch of G7413: signal is true;
	signal G7414: std_logic; attribute dont_touch of G7414: signal is true;
	signal G7415: std_logic; attribute dont_touch of G7415: signal is true;
	signal G7416: std_logic; attribute dont_touch of G7416: signal is true;
	signal G7419: std_logic; attribute dont_touch of G7419: signal is true;
	signal G7420: std_logic; attribute dont_touch of G7420: signal is true;
	signal G7421: std_logic; attribute dont_touch of G7421: signal is true;
	signal G7422: std_logic; attribute dont_touch of G7422: signal is true;
	signal G7425: std_logic; attribute dont_touch of G7425: signal is true;
	signal G7426: std_logic; attribute dont_touch of G7426: signal is true;
	signal G7427: std_logic; attribute dont_touch of G7427: signal is true;
	signal G7430: std_logic; attribute dont_touch of G7430: signal is true;
	signal G7431: std_logic; attribute dont_touch of G7431: signal is true;
	signal G7432: std_logic; attribute dont_touch of G7432: signal is true;
	signal G7435: std_logic; attribute dont_touch of G7435: signal is true;
	signal G7436: std_logic; attribute dont_touch of G7436: signal is true;
	signal G7437: std_logic; attribute dont_touch of G7437: signal is true;
	signal G7438: std_logic; attribute dont_touch of G7438: signal is true;
	signal G7439: std_logic; attribute dont_touch of G7439: signal is true;
	signal G7440: std_logic; attribute dont_touch of G7440: signal is true;
	signal G7441: std_logic; attribute dont_touch of G7441: signal is true;
	signal G7442: std_logic; attribute dont_touch of G7442: signal is true;
	signal G7443: std_logic; attribute dont_touch of G7443: signal is true;
	signal G7444: std_logic; attribute dont_touch of G7444: signal is true;
	signal G7445: std_logic; attribute dont_touch of G7445: signal is true;
	signal G7446: std_logic; attribute dont_touch of G7446: signal is true;
	signal G7449: std_logic; attribute dont_touch of G7449: signal is true;
	signal G7450: std_logic; attribute dont_touch of G7450: signal is true;
	signal G7453: std_logic; attribute dont_touch of G7453: signal is true;
	signal G7454: std_logic; attribute dont_touch of G7454: signal is true;
	signal G7457: std_logic; attribute dont_touch of G7457: signal is true;
	signal G7458: std_logic; attribute dont_touch of G7458: signal is true;
	signal G7459: std_logic; attribute dont_touch of G7459: signal is true;
	signal G7460: std_logic; attribute dont_touch of G7460: signal is true;
	signal G7463: std_logic; attribute dont_touch of G7463: signal is true;
	signal G7464: std_logic; attribute dont_touch of G7464: signal is true;
	signal G7465: std_logic; attribute dont_touch of G7465: signal is true;
	signal G7466: std_logic; attribute dont_touch of G7466: signal is true;
	signal G7467: std_logic; attribute dont_touch of G7467: signal is true;
	signal G7470: std_logic; attribute dont_touch of G7470: signal is true;
	signal G7471: std_logic; attribute dont_touch of G7471: signal is true;
	signal G7472: std_logic; attribute dont_touch of G7472: signal is true;
	signal G7473: std_logic; attribute dont_touch of G7473: signal is true;
	signal G7476: std_logic; attribute dont_touch of G7476: signal is true;
	signal G7477: std_logic; attribute dont_touch of G7477: signal is true;
	signal G7478: std_logic; attribute dont_touch of G7478: signal is true;
	signal G7479: std_logic; attribute dont_touch of G7479: signal is true;
	signal G7496: std_logic; attribute dont_touch of G7496: signal is true;
	signal G7497: std_logic; attribute dont_touch of G7497: signal is true;
	signal G7500: std_logic; attribute dont_touch of G7500: signal is true;
	signal G7501: std_logic; attribute dont_touch of G7501: signal is true;
	signal G7502: std_logic; attribute dont_touch of G7502: signal is true;
	signal G7503: std_logic; attribute dont_touch of G7503: signal is true;
	signal G7504: std_logic; attribute dont_touch of G7504: signal is true;
	signal G7505: std_logic; attribute dont_touch of G7505: signal is true;
	signal G7508: std_logic; attribute dont_touch of G7508: signal is true;
	signal G7509: std_logic; attribute dont_touch of G7509: signal is true;
	signal G7510: std_logic; attribute dont_touch of G7510: signal is true;
	signal G7511: std_logic; attribute dont_touch of G7511: signal is true;
	signal G7512: std_logic; attribute dont_touch of G7512: signal is true;
	signal G7515: std_logic; attribute dont_touch of G7515: signal is true;
	signal G7516: std_logic; attribute dont_touch of G7516: signal is true;
	signal G7519: std_logic; attribute dont_touch of G7519: signal is true;
	signal G7520: std_logic; attribute dont_touch of G7520: signal is true;
	signal G7521: std_logic; attribute dont_touch of G7521: signal is true;
	signal G7522: std_logic; attribute dont_touch of G7522: signal is true;
	signal G7523: std_logic; attribute dont_touch of G7523: signal is true;
	signal G7524: std_logic; attribute dont_touch of G7524: signal is true;
	signal G7525: std_logic; attribute dont_touch of G7525: signal is true;
	signal G7526: std_logic; attribute dont_touch of G7526: signal is true;
	signal G7527: std_logic; attribute dont_touch of G7527: signal is true;
	signal G7530: std_logic; attribute dont_touch of G7530: signal is true;
	signal G7531: std_logic; attribute dont_touch of G7531: signal is true;
	signal G7532: std_logic; attribute dont_touch of G7532: signal is true;
	signal G7533: std_logic; attribute dont_touch of G7533: signal is true;
	signal G7534: std_logic; attribute dont_touch of G7534: signal is true;
	signal G7535: std_logic; attribute dont_touch of G7535: signal is true;
	signal G7536: std_logic; attribute dont_touch of G7536: signal is true;
	signal G7537: std_logic; attribute dont_touch of G7537: signal is true;
	signal G7538: std_logic; attribute dont_touch of G7538: signal is true;
	signal G7539: std_logic; attribute dont_touch of G7539: signal is true;
	signal G7540: std_logic; attribute dont_touch of G7540: signal is true;
	signal G7541: std_logic; attribute dont_touch of G7541: signal is true;
	signal G7542: std_logic; attribute dont_touch of G7542: signal is true;
	signal G7543: std_logic; attribute dont_touch of G7543: signal is true;
	signal G7544: std_logic; attribute dont_touch of G7544: signal is true;
	signal G7545: std_logic; attribute dont_touch of G7545: signal is true;
	signal G7546: std_logic; attribute dont_touch of G7546: signal is true;
	signal G7547: std_logic; attribute dont_touch of G7547: signal is true;
	signal G7548: std_logic; attribute dont_touch of G7548: signal is true;
	signal G7549: std_logic; attribute dont_touch of G7549: signal is true;
	signal G7550: std_logic; attribute dont_touch of G7550: signal is true;
	signal G7555: std_logic; attribute dont_touch of G7555: signal is true;
	signal G7556: std_logic; attribute dont_touch of G7556: signal is true;
	signal G7557: std_logic; attribute dont_touch of G7557: signal is true;
	signal G7558: std_logic; attribute dont_touch of G7558: signal is true;
	signal G7559: std_logic; attribute dont_touch of G7559: signal is true;
	signal G7560: std_logic; attribute dont_touch of G7560: signal is true;
	signal G7561: std_logic; attribute dont_touch of G7561: signal is true;
	signal G7562: std_logic; attribute dont_touch of G7562: signal is true;
	signal G7567: std_logic; attribute dont_touch of G7567: signal is true;
	signal G7568: std_logic; attribute dont_touch of G7568: signal is true;
	signal G7569: std_logic; attribute dont_touch of G7569: signal is true;
	signal G7570: std_logic; attribute dont_touch of G7570: signal is true;
	signal G7571: std_logic; attribute dont_touch of G7571: signal is true;
	signal G7572: std_logic; attribute dont_touch of G7572: signal is true;
	signal G7573: std_logic; attribute dont_touch of G7573: signal is true;
	signal G7574: std_logic; attribute dont_touch of G7574: signal is true;
	signal G7579: std_logic; attribute dont_touch of G7579: signal is true;
	signal G7580: std_logic; attribute dont_touch of G7580: signal is true;
	signal G7581: std_logic; attribute dont_touch of G7581: signal is true;
	signal G7582: std_logic; attribute dont_touch of G7582: signal is true;
	signal G7583: std_logic; attribute dont_touch of G7583: signal is true;
	signal G7584: std_logic; attribute dont_touch of G7584: signal is true;
	signal G7585: std_logic; attribute dont_touch of G7585: signal is true;
	signal G7586: std_logic; attribute dont_touch of G7586: signal is true;
	signal G7587: std_logic; attribute dont_touch of G7587: signal is true;
	signal G7588: std_logic; attribute dont_touch of G7588: signal is true;
	signal G7589: std_logic; attribute dont_touch of G7589: signal is true;
	signal G7590: std_logic; attribute dont_touch of G7590: signal is true;
	signal G7591: std_logic; attribute dont_touch of G7591: signal is true;
	signal G7592: std_logic; attribute dont_touch of G7592: signal is true;
	signal G7593: std_logic; attribute dont_touch of G7593: signal is true;
	signal G7594: std_logic; attribute dont_touch of G7594: signal is true;
	signal G7595: std_logic; attribute dont_touch of G7595: signal is true;
	signal G7596: std_logic; attribute dont_touch of G7596: signal is true;
	signal G7597: std_logic; attribute dont_touch of G7597: signal is true;
	signal G7598: std_logic; attribute dont_touch of G7598: signal is true;
	signal G7599: std_logic; attribute dont_touch of G7599: signal is true;
	signal G7600: std_logic; attribute dont_touch of G7600: signal is true;
	signal G7601: std_logic; attribute dont_touch of G7601: signal is true;
	signal G7602: std_logic; attribute dont_touch of G7602: signal is true;
	signal G7603: std_logic; attribute dont_touch of G7603: signal is true;
	signal G7604: std_logic; attribute dont_touch of G7604: signal is true;
	signal G7605: std_logic; attribute dont_touch of G7605: signal is true;
	signal G7606: std_logic; attribute dont_touch of G7606: signal is true;
	signal G7607: std_logic; attribute dont_touch of G7607: signal is true;
	signal G7608: std_logic; attribute dont_touch of G7608: signal is true;
	signal G7609: std_logic; attribute dont_touch of G7609: signal is true;
	signal G7610: std_logic; attribute dont_touch of G7610: signal is true;
	signal G7611: std_logic; attribute dont_touch of G7611: signal is true;
	signal G7612: std_logic; attribute dont_touch of G7612: signal is true;
	signal G7613: std_logic; attribute dont_touch of G7613: signal is true;
	signal G7614: std_logic; attribute dont_touch of G7614: signal is true;
	signal G7615: std_logic; attribute dont_touch of G7615: signal is true;
	signal G7616: std_logic; attribute dont_touch of G7616: signal is true;
	signal G7617: std_logic; attribute dont_touch of G7617: signal is true;
	signal G7618: std_logic; attribute dont_touch of G7618: signal is true;
	signal G7619: std_logic; attribute dont_touch of G7619: signal is true;
	signal G7620: std_logic; attribute dont_touch of G7620: signal is true;
	signal G7621: std_logic; attribute dont_touch of G7621: signal is true;
	signal G7622: std_logic; attribute dont_touch of G7622: signal is true;
	signal G7623: std_logic; attribute dont_touch of G7623: signal is true;
	signal G7624: std_logic; attribute dont_touch of G7624: signal is true;
	signal G7625: std_logic; attribute dont_touch of G7625: signal is true;
	signal G7626: std_logic; attribute dont_touch of G7626: signal is true;
	signal G7627: std_logic; attribute dont_touch of G7627: signal is true;
	signal G7628: std_logic; attribute dont_touch of G7628: signal is true;
	signal G7629: std_logic; attribute dont_touch of G7629: signal is true;
	signal G7630: std_logic; attribute dont_touch of G7630: signal is true;
	signal G7631: std_logic; attribute dont_touch of G7631: signal is true;
	signal G7632: std_logic; attribute dont_touch of G7632: signal is true;
	signal G7633: std_logic; attribute dont_touch of G7633: signal is true;
	signal G7634: std_logic; attribute dont_touch of G7634: signal is true;
	signal G7635: std_logic; attribute dont_touch of G7635: signal is true;
	signal G7636: std_logic; attribute dont_touch of G7636: signal is true;
	signal G7637: std_logic; attribute dont_touch of G7637: signal is true;
	signal G7638: std_logic; attribute dont_touch of G7638: signal is true;
	signal G7648: std_logic; attribute dont_touch of G7648: signal is true;
	signal G7649: std_logic; attribute dont_touch of G7649: signal is true;
	signal G7650: std_logic; attribute dont_touch of G7650: signal is true;
	signal G7651: std_logic; attribute dont_touch of G7651: signal is true;
	signal G7656: std_logic; attribute dont_touch of G7656: signal is true;
	signal G7657: std_logic; attribute dont_touch of G7657: signal is true;
	signal G7658: std_logic; attribute dont_touch of G7658: signal is true;
	signal G7659: std_logic; attribute dont_touch of G7659: signal is true;
	signal G7660: std_logic; attribute dont_touch of G7660: signal is true;
	signal G7661: std_logic; attribute dont_touch of G7661: signal is true;
	signal G7662: std_logic; attribute dont_touch of G7662: signal is true;
	signal G7663: std_logic; attribute dont_touch of G7663: signal is true;
	signal G7664: std_logic; attribute dont_touch of G7664: signal is true;
	signal G7669: std_logic; attribute dont_touch of G7669: signal is true;
	signal G7670: std_logic; attribute dont_touch of G7670: signal is true;
	signal G7671: std_logic; attribute dont_touch of G7671: signal is true;
	signal G7672: std_logic; attribute dont_touch of G7672: signal is true;
	signal G7673: std_logic; attribute dont_touch of G7673: signal is true;
	signal G7674: std_logic; attribute dont_touch of G7674: signal is true;
	signal G7675: std_logic; attribute dont_touch of G7675: signal is true;
	signal G7676: std_logic; attribute dont_touch of G7676: signal is true;
	signal G7677: std_logic; attribute dont_touch of G7677: signal is true;
	signal G7678: std_logic; attribute dont_touch of G7678: signal is true;
	signal G7679: std_logic; attribute dont_touch of G7679: signal is true;
	signal G7680: std_logic; attribute dont_touch of G7680: signal is true;
	signal G7681: std_logic; attribute dont_touch of G7681: signal is true;
	signal G7682: std_logic; attribute dont_touch of G7682: signal is true;
	signal G7683: std_logic; attribute dont_touch of G7683: signal is true;
	signal G7684: std_logic; attribute dont_touch of G7684: signal is true;
	signal G7685: std_logic; attribute dont_touch of G7685: signal is true;
	signal G7686: std_logic; attribute dont_touch of G7686: signal is true;
	signal G7687: std_logic; attribute dont_touch of G7687: signal is true;
	signal G7688: std_logic; attribute dont_touch of G7688: signal is true;
	signal G7689: std_logic; attribute dont_touch of G7689: signal is true;
	signal G7692: std_logic; attribute dont_touch of G7692: signal is true;
	signal G7693: std_logic; attribute dont_touch of G7693: signal is true;
	signal G7696: std_logic; attribute dont_touch of G7696: signal is true;
	signal G7697: std_logic; attribute dont_touch of G7697: signal is true;
	signal G7702: std_logic; attribute dont_touch of G7702: signal is true;
	signal G7703: std_logic; attribute dont_touch of G7703: signal is true;
	signal G7704: std_logic; attribute dont_touch of G7704: signal is true;
	signal G7705: std_logic; attribute dont_touch of G7705: signal is true;
	signal G7706: std_logic; attribute dont_touch of G7706: signal is true;
	signal G7707: std_logic; attribute dont_touch of G7707: signal is true;
	signal G7708: std_logic; attribute dont_touch of G7708: signal is true;
	signal G7709: std_logic; attribute dont_touch of G7709: signal is true;
	signal G7710: std_logic; attribute dont_touch of G7710: signal is true;
	signal G7711: std_logic; attribute dont_touch of G7711: signal is true;
	signal G7712: std_logic; attribute dont_touch of G7712: signal is true;
	signal G7717: std_logic; attribute dont_touch of G7717: signal is true;
	signal G7718: std_logic; attribute dont_touch of G7718: signal is true;
	signal G7719: std_logic; attribute dont_touch of G7719: signal is true;
	signal G7720: std_logic; attribute dont_touch of G7720: signal is true;
	signal G7721: std_logic; attribute dont_touch of G7721: signal is true;
	signal G7722: std_logic; attribute dont_touch of G7722: signal is true;
	signal G7723: std_logic; attribute dont_touch of G7723: signal is true;
	signal G7724: std_logic; attribute dont_touch of G7724: signal is true;
	signal G7725: std_logic; attribute dont_touch of G7725: signal is true;
	signal G7726: std_logic; attribute dont_touch of G7726: signal is true;
	signal G7727: std_logic; attribute dont_touch of G7727: signal is true;
	signal G7728: std_logic; attribute dont_touch of G7728: signal is true;
	signal G7729: std_logic; attribute dont_touch of G7729: signal is true;
	signal G7730: std_logic; attribute dont_touch of G7730: signal is true;
	signal G7731: std_logic; attribute dont_touch of G7731: signal is true;
	signal G7732: std_logic; attribute dont_touch of G7732: signal is true;
	signal G7733: std_logic; attribute dont_touch of G7733: signal is true;
	signal G7734: std_logic; attribute dont_touch of G7734: signal is true;
	signal G7735: std_logic; attribute dont_touch of G7735: signal is true;
	signal G7736: std_logic; attribute dont_touch of G7736: signal is true;
	signal G7737: std_logic; attribute dont_touch of G7737: signal is true;
	signal G7738: std_logic; attribute dont_touch of G7738: signal is true;
	signal G7739: std_logic; attribute dont_touch of G7739: signal is true;
	signal G7740: std_logic; attribute dont_touch of G7740: signal is true;
	signal G7741: std_logic; attribute dont_touch of G7741: signal is true;
	signal G7742: std_logic; attribute dont_touch of G7742: signal is true;
	signal G7743: std_logic; attribute dont_touch of G7743: signal is true;
	signal G7745: std_logic; attribute dont_touch of G7745: signal is true;
	signal G7746: std_logic; attribute dont_touch of G7746: signal is true;
	signal G7747: std_logic; attribute dont_touch of G7747: signal is true;
	signal G7748: std_logic; attribute dont_touch of G7748: signal is true;
	signal G7749: std_logic; attribute dont_touch of G7749: signal is true;
	signal G7750: std_logic; attribute dont_touch of G7750: signal is true;
	signal G7751: std_logic; attribute dont_touch of G7751: signal is true;
	signal G7752: std_logic; attribute dont_touch of G7752: signal is true;
	signal G7753: std_logic; attribute dont_touch of G7753: signal is true;
	signal G7754: std_logic; attribute dont_touch of G7754: signal is true;
	signal G7755: std_logic; attribute dont_touch of G7755: signal is true;
	signal G7756: std_logic; attribute dont_touch of G7756: signal is true;
	signal G7757: std_logic; attribute dont_touch of G7757: signal is true;
	signal G7758: std_logic; attribute dont_touch of G7758: signal is true;
	signal G7759: std_logic; attribute dont_touch of G7759: signal is true;
	signal G7760: std_logic; attribute dont_touch of G7760: signal is true;
	signal G7761: std_logic; attribute dont_touch of G7761: signal is true;
	signal G7762: std_logic; attribute dont_touch of G7762: signal is true;
	signal G7763: std_logic; attribute dont_touch of G7763: signal is true;
	signal G7764: std_logic; attribute dont_touch of G7764: signal is true;
	signal G7765: std_logic; attribute dont_touch of G7765: signal is true;
	signal G7766: std_logic; attribute dont_touch of G7766: signal is true;
	signal G7767: std_logic; attribute dont_touch of G7767: signal is true;
	signal G7768: std_logic; attribute dont_touch of G7768: signal is true;
	signal G7769: std_logic; attribute dont_touch of G7769: signal is true;
	signal G7770: std_logic; attribute dont_touch of G7770: signal is true;
	signal G7771: std_logic; attribute dont_touch of G7771: signal is true;
	signal G7772: std_logic; attribute dont_touch of G7772: signal is true;
	signal G7773: std_logic; attribute dont_touch of G7773: signal is true;
	signal G7774: std_logic; attribute dont_touch of G7774: signal is true;
	signal G7775: std_logic; attribute dont_touch of G7775: signal is true;
	signal G7776: std_logic; attribute dont_touch of G7776: signal is true;
	signal G7777: std_logic; attribute dont_touch of G7777: signal is true;
	signal G7778: std_logic; attribute dont_touch of G7778: signal is true;
	signal G7779: std_logic; attribute dont_touch of G7779: signal is true;
	signal G7780: std_logic; attribute dont_touch of G7780: signal is true;
	signal G7781: std_logic; attribute dont_touch of G7781: signal is true;
	signal G7782: std_logic; attribute dont_touch of G7782: signal is true;
	signal G7783: std_logic; attribute dont_touch of G7783: signal is true;
	signal G7784: std_logic; attribute dont_touch of G7784: signal is true;
	signal G7785: std_logic; attribute dont_touch of G7785: signal is true;
	signal G7786: std_logic; attribute dont_touch of G7786: signal is true;
	signal G7787: std_logic; attribute dont_touch of G7787: signal is true;
	signal G7788: std_logic; attribute dont_touch of G7788: signal is true;
	signal G7789: std_logic; attribute dont_touch of G7789: signal is true;
	signal G7790: std_logic; attribute dont_touch of G7790: signal is true;
	signal G7791: std_logic; attribute dont_touch of G7791: signal is true;
	signal G7792: std_logic; attribute dont_touch of G7792: signal is true;
	signal G7793: std_logic; attribute dont_touch of G7793: signal is true;
	signal G7794: std_logic; attribute dont_touch of G7794: signal is true;
	signal G7795: std_logic; attribute dont_touch of G7795: signal is true;
	signal G7796: std_logic; attribute dont_touch of G7796: signal is true;
	signal G7797: std_logic; attribute dont_touch of G7797: signal is true;
	signal G7798: std_logic; attribute dont_touch of G7798: signal is true;
	signal G7799: std_logic; attribute dont_touch of G7799: signal is true;
	signal G7800: std_logic; attribute dont_touch of G7800: signal is true;
	signal G7801: std_logic; attribute dont_touch of G7801: signal is true;
	signal G7802: std_logic; attribute dont_touch of G7802: signal is true;
	signal G7803: std_logic; attribute dont_touch of G7803: signal is true;
	signal G7804: std_logic; attribute dont_touch of G7804: signal is true;
	signal G7805: std_logic; attribute dont_touch of G7805: signal is true;
	signal G7806: std_logic; attribute dont_touch of G7806: signal is true;
	signal G7807: std_logic; attribute dont_touch of G7807: signal is true;
	signal G7808: std_logic; attribute dont_touch of G7808: signal is true;
	signal G7809: std_logic; attribute dont_touch of G7809: signal is true;
	signal G7810: std_logic; attribute dont_touch of G7810: signal is true;
	signal G7811: std_logic; attribute dont_touch of G7811: signal is true;
	signal G7812: std_logic; attribute dont_touch of G7812: signal is true;
	signal G7813: std_logic; attribute dont_touch of G7813: signal is true;
	signal G7814: std_logic; attribute dont_touch of G7814: signal is true;
	signal G7815: std_logic; attribute dont_touch of G7815: signal is true;
	signal G7816: std_logic; attribute dont_touch of G7816: signal is true;
	signal G7817: std_logic; attribute dont_touch of G7817: signal is true;
	signal G7818: std_logic; attribute dont_touch of G7818: signal is true;
	signal G7819: std_logic; attribute dont_touch of G7819: signal is true;
	signal G7820: std_logic; attribute dont_touch of G7820: signal is true;
	signal G7821: std_logic; attribute dont_touch of G7821: signal is true;
	signal G7822: std_logic; attribute dont_touch of G7822: signal is true;
	signal G7823: std_logic; attribute dont_touch of G7823: signal is true;
	signal G7824: std_logic; attribute dont_touch of G7824: signal is true;
	signal G7825: std_logic; attribute dont_touch of G7825: signal is true;
	signal G7826: std_logic; attribute dont_touch of G7826: signal is true;
	signal G7843: std_logic; attribute dont_touch of G7843: signal is true;
	signal G7844: std_logic; attribute dont_touch of G7844: signal is true;
	signal G7845: std_logic; attribute dont_touch of G7845: signal is true;
	signal G7846: std_logic; attribute dont_touch of G7846: signal is true;
	signal G7847: std_logic; attribute dont_touch of G7847: signal is true;
	signal G7848: std_logic; attribute dont_touch of G7848: signal is true;
	signal G7849: std_logic; attribute dont_touch of G7849: signal is true;
	signal G7850: std_logic; attribute dont_touch of G7850: signal is true;
	signal G7851: std_logic; attribute dont_touch of G7851: signal is true;
	signal G7852: std_logic; attribute dont_touch of G7852: signal is true;
	signal G7853: std_logic; attribute dont_touch of G7853: signal is true;
	signal G7872: std_logic; attribute dont_touch of G7872: signal is true;
	signal G7876: std_logic; attribute dont_touch of G7876: signal is true;
	signal G7877: std_logic; attribute dont_touch of G7877: signal is true;
	signal G7878: std_logic; attribute dont_touch of G7878: signal is true;
	signal G7879: std_logic; attribute dont_touch of G7879: signal is true;
	signal G7880: std_logic; attribute dont_touch of G7880: signal is true;
	signal G7881: std_logic; attribute dont_touch of G7881: signal is true;
	signal G7882: std_logic; attribute dont_touch of G7882: signal is true;
	signal G7883: std_logic; attribute dont_touch of G7883: signal is true;
	signal G7884: std_logic; attribute dont_touch of G7884: signal is true;
	signal G7885: std_logic; attribute dont_touch of G7885: signal is true;
	signal G7886: std_logic; attribute dont_touch of G7886: signal is true;
	signal G7887: std_logic; attribute dont_touch of G7887: signal is true;
	signal G7888: std_logic; attribute dont_touch of G7888: signal is true;
	signal G7889: std_logic; attribute dont_touch of G7889: signal is true;
	signal G7890: std_logic; attribute dont_touch of G7890: signal is true;
	signal G7891: std_logic; attribute dont_touch of G7891: signal is true;
	signal G7892: std_logic; attribute dont_touch of G7892: signal is true;
	signal G7893: std_logic; attribute dont_touch of G7893: signal is true;
	signal G7894: std_logic; attribute dont_touch of G7894: signal is true;
	signal G7895: std_logic; attribute dont_touch of G7895: signal is true;
	signal G7896: std_logic; attribute dont_touch of G7896: signal is true;
	signal G7897: std_logic; attribute dont_touch of G7897: signal is true;
	signal G7898: std_logic; attribute dont_touch of G7898: signal is true;
	signal G7899: std_logic; attribute dont_touch of G7899: signal is true;
	signal G7900: std_logic; attribute dont_touch of G7900: signal is true;
	signal G7901: std_logic; attribute dont_touch of G7901: signal is true;
	signal G7902: std_logic; attribute dont_touch of G7902: signal is true;
	signal G7903: std_logic; attribute dont_touch of G7903: signal is true;
	signal G7904: std_logic; attribute dont_touch of G7904: signal is true;
	signal G7905: std_logic; attribute dont_touch of G7905: signal is true;
	signal G7906: std_logic; attribute dont_touch of G7906: signal is true;
	signal G7907: std_logic; attribute dont_touch of G7907: signal is true;
	signal G7908: std_logic; attribute dont_touch of G7908: signal is true;
	signal G7909: std_logic; attribute dont_touch of G7909: signal is true;
	signal G7910: std_logic; attribute dont_touch of G7910: signal is true;
	signal G7911: std_logic; attribute dont_touch of G7911: signal is true;
	signal G7912: std_logic; attribute dont_touch of G7912: signal is true;
	signal G7913: std_logic; attribute dont_touch of G7913: signal is true;
	signal G7914: std_logic; attribute dont_touch of G7914: signal is true;
	signal G7915: std_logic; attribute dont_touch of G7915: signal is true;
	signal G7916: std_logic; attribute dont_touch of G7916: signal is true;
	signal G7917: std_logic; attribute dont_touch of G7917: signal is true;
	signal G7918: std_logic; attribute dont_touch of G7918: signal is true;
	signal G7919: std_logic; attribute dont_touch of G7919: signal is true;
	signal G7920: std_logic; attribute dont_touch of G7920: signal is true;
	signal G7921: std_logic; attribute dont_touch of G7921: signal is true;
	signal G7922: std_logic; attribute dont_touch of G7922: signal is true;
	signal G7923: std_logic; attribute dont_touch of G7923: signal is true;
	signal G7924: std_logic; attribute dont_touch of G7924: signal is true;
	signal G7925: std_logic; attribute dont_touch of G7925: signal is true;
	signal G7926: std_logic; attribute dont_touch of G7926: signal is true;
	signal G7927: std_logic; attribute dont_touch of G7927: signal is true;
	signal G7928: std_logic; attribute dont_touch of G7928: signal is true;
	signal G7929: std_logic; attribute dont_touch of G7929: signal is true;
	signal G7930: std_logic; attribute dont_touch of G7930: signal is true;
	signal G7931: std_logic; attribute dont_touch of G7931: signal is true;
	signal G7932: std_logic; attribute dont_touch of G7932: signal is true;
	signal G7933: std_logic; attribute dont_touch of G7933: signal is true;
	signal G7934: std_logic; attribute dont_touch of G7934: signal is true;
	signal G7935: std_logic; attribute dont_touch of G7935: signal is true;
	signal G7936: std_logic; attribute dont_touch of G7936: signal is true;
	signal G7937: std_logic; attribute dont_touch of G7937: signal is true;
	signal G7938: std_logic; attribute dont_touch of G7938: signal is true;
	signal G7939: std_logic; attribute dont_touch of G7939: signal is true;
	signal G7940: std_logic; attribute dont_touch of G7940: signal is true;
	signal G7941: std_logic; attribute dont_touch of G7941: signal is true;
	signal G7942: std_logic; attribute dont_touch of G7942: signal is true;
	signal G7943: std_logic; attribute dont_touch of G7943: signal is true;
	signal G7944: std_logic; attribute dont_touch of G7944: signal is true;
	signal G7945: std_logic; attribute dont_touch of G7945: signal is true;
	signal G7946: std_logic; attribute dont_touch of G7946: signal is true;
	signal G7947: std_logic; attribute dont_touch of G7947: signal is true;
	signal G7948: std_logic; attribute dont_touch of G7948: signal is true;
	signal G7949: std_logic; attribute dont_touch of G7949: signal is true;
	signal G7950: std_logic; attribute dont_touch of G7950: signal is true;
	signal G7951: std_logic; attribute dont_touch of G7951: signal is true;
	signal G7952: std_logic; attribute dont_touch of G7952: signal is true;
	signal G7953: std_logic; attribute dont_touch of G7953: signal is true;
	signal G7954: std_logic; attribute dont_touch of G7954: signal is true;
	signal G7955: std_logic; attribute dont_touch of G7955: signal is true;
	signal G7956: std_logic; attribute dont_touch of G7956: signal is true;
	signal G7957: std_logic; attribute dont_touch of G7957: signal is true;
	signal G7958: std_logic; attribute dont_touch of G7958: signal is true;
	signal G7959: std_logic; attribute dont_touch of G7959: signal is true;
	signal G7960: std_logic; attribute dont_touch of G7960: signal is true;
	signal G7961: std_logic; attribute dont_touch of G7961: signal is true;
	signal G7962: std_logic; attribute dont_touch of G7962: signal is true;
	signal G7963: std_logic; attribute dont_touch of G7963: signal is true;
	signal G7964: std_logic; attribute dont_touch of G7964: signal is true;
	signal G7965: std_logic; attribute dont_touch of G7965: signal is true;
	signal G7966: std_logic; attribute dont_touch of G7966: signal is true;
	signal G7967: std_logic; attribute dont_touch of G7967: signal is true;
	signal G7970: std_logic; attribute dont_touch of G7970: signal is true;
	signal G7971: std_logic; attribute dont_touch of G7971: signal is true;
	signal G7972: std_logic; attribute dont_touch of G7972: signal is true;
	signal G7975: std_logic; attribute dont_touch of G7975: signal is true;
	signal G7976: std_logic; attribute dont_touch of G7976: signal is true;
	signal G7977: std_logic; attribute dont_touch of G7977: signal is true;
	signal G7978: std_logic; attribute dont_touch of G7978: signal is true;
	signal G7979: std_logic; attribute dont_touch of G7979: signal is true;
	signal G7980: std_logic; attribute dont_touch of G7980: signal is true;
	signal G7981: std_logic; attribute dont_touch of G7981: signal is true;
	signal G7982: std_logic; attribute dont_touch of G7982: signal is true;
	signal G7983: std_logic; attribute dont_touch of G7983: signal is true;
	signal G7984: std_logic; attribute dont_touch of G7984: signal is true;
	signal G7985: std_logic; attribute dont_touch of G7985: signal is true;
	signal G7986: std_logic; attribute dont_touch of G7986: signal is true;
	signal G7987: std_logic; attribute dont_touch of G7987: signal is true;
	signal G7988: std_logic; attribute dont_touch of G7988: signal is true;
	signal G7989: std_logic; attribute dont_touch of G7989: signal is true;
	signal G7990: std_logic; attribute dont_touch of G7990: signal is true;
	signal G7991: std_logic; attribute dont_touch of G7991: signal is true;
	signal G7992: std_logic; attribute dont_touch of G7992: signal is true;
	signal G7993: std_logic; attribute dont_touch of G7993: signal is true;
	signal G7994: std_logic; attribute dont_touch of G7994: signal is true;
	signal G7995: std_logic; attribute dont_touch of G7995: signal is true;
	signal G7996: std_logic; attribute dont_touch of G7996: signal is true;
	signal G7997: std_logic; attribute dont_touch of G7997: signal is true;
	signal G7998: std_logic; attribute dont_touch of G7998: signal is true;
	signal G7999: std_logic; attribute dont_touch of G7999: signal is true;
	signal G8000: std_logic; attribute dont_touch of G8000: signal is true;
	signal G8001: std_logic; attribute dont_touch of G8001: signal is true;
	signal G8002: std_logic; attribute dont_touch of G8002: signal is true;
	signal G8003: std_logic; attribute dont_touch of G8003: signal is true;
	signal G8004: std_logic; attribute dont_touch of G8004: signal is true;
	signal G8005: std_logic; attribute dont_touch of G8005: signal is true;
	signal G8006: std_logic; attribute dont_touch of G8006: signal is true;
	signal G8007: std_logic; attribute dont_touch of G8007: signal is true;
	signal G8008: std_logic; attribute dont_touch of G8008: signal is true;
	signal G8009: std_logic; attribute dont_touch of G8009: signal is true;
	signal G8010: std_logic; attribute dont_touch of G8010: signal is true;
	signal G8011: std_logic; attribute dont_touch of G8011: signal is true;
	signal G8014: std_logic; attribute dont_touch of G8014: signal is true;
	signal G8015: std_logic; attribute dont_touch of G8015: signal is true;
	signal G8018: std_logic; attribute dont_touch of G8018: signal is true;
	signal G8019: std_logic; attribute dont_touch of G8019: signal is true;
	signal G8020: std_logic; attribute dont_touch of G8020: signal is true;
	signal G8023: std_logic; attribute dont_touch of G8023: signal is true;
	signal G8024: std_logic; attribute dont_touch of G8024: signal is true;
	signal G8025: std_logic; attribute dont_touch of G8025: signal is true;
	signal G8028: std_logic; attribute dont_touch of G8028: signal is true;
	signal G8029: std_logic; attribute dont_touch of G8029: signal is true;
	signal G8032: std_logic; attribute dont_touch of G8032: signal is true;
	signal G8033: std_logic; attribute dont_touch of G8033: signal is true;
	signal G8036: std_logic; attribute dont_touch of G8036: signal is true;
	signal G8039: std_logic; attribute dont_touch of G8039: signal is true;
	signal G8040: std_logic; attribute dont_touch of G8040: signal is true;
	signal G8041: std_logic; attribute dont_touch of G8041: signal is true;
	signal G8042: std_logic; attribute dont_touch of G8042: signal is true;
	signal G8043: std_logic; attribute dont_touch of G8043: signal is true;
	signal G8044: std_logic; attribute dont_touch of G8044: signal is true;
	signal G8045: std_logic; attribute dont_touch of G8045: signal is true;
	signal G8046: std_logic; attribute dont_touch of G8046: signal is true;
	signal G8047: std_logic; attribute dont_touch of G8047: signal is true;
	signal G8048: std_logic; attribute dont_touch of G8048: signal is true;
	signal G8049: std_logic; attribute dont_touch of G8049: signal is true;
	signal G8050: std_logic; attribute dont_touch of G8050: signal is true;
	signal G8051: std_logic; attribute dont_touch of G8051: signal is true;
	signal G8052: std_logic; attribute dont_touch of G8052: signal is true;
	signal G8053: std_logic; attribute dont_touch of G8053: signal is true;
	signal G8054: std_logic; attribute dont_touch of G8054: signal is true;
	signal G8055: std_logic; attribute dont_touch of G8055: signal is true;
	signal G8056: std_logic; attribute dont_touch of G8056: signal is true;
	signal G8059: std_logic; attribute dont_touch of G8059: signal is true;
	signal G8060: std_logic; attribute dont_touch of G8060: signal is true;
	signal G8063: std_logic; attribute dont_touch of G8063: signal is true;
	signal G8064: std_logic; attribute dont_touch of G8064: signal is true;
	signal G8065: std_logic; attribute dont_touch of G8065: signal is true;
	signal G8066: std_logic; attribute dont_touch of G8066: signal is true;
	signal G8067: std_logic; attribute dont_touch of G8067: signal is true;
	signal G8068: std_logic; attribute dont_touch of G8068: signal is true;
	signal G8069: std_logic; attribute dont_touch of G8069: signal is true;
	signal G8070: std_logic; attribute dont_touch of G8070: signal is true;
	signal G8071: std_logic; attribute dont_touch of G8071: signal is true;
	signal G8072: std_logic; attribute dont_touch of G8072: signal is true;
	signal G8073: std_logic; attribute dont_touch of G8073: signal is true;
	signal G8074: std_logic; attribute dont_touch of G8074: signal is true;
	signal G8075: std_logic; attribute dont_touch of G8075: signal is true;
	signal G8076: std_logic; attribute dont_touch of G8076: signal is true;
	signal G8077: std_logic; attribute dont_touch of G8077: signal is true;
	signal G8078: std_logic; attribute dont_touch of G8078: signal is true;
	signal G8079: std_logic; attribute dont_touch of G8079: signal is true;
	signal G8080: std_logic; attribute dont_touch of G8080: signal is true;
	signal G8081: std_logic; attribute dont_touch of G8081: signal is true;
	signal G8085: std_logic; attribute dont_touch of G8085: signal is true;
	signal G8089: std_logic; attribute dont_touch of G8089: signal is true;
	signal G8093: std_logic; attribute dont_touch of G8093: signal is true;
	signal G8094: std_logic; attribute dont_touch of G8094: signal is true;
	signal G8095: std_logic; attribute dont_touch of G8095: signal is true;
	signal G8096: std_logic; attribute dont_touch of G8096: signal is true;
	signal G8097: std_logic; attribute dont_touch of G8097: signal is true;
	signal G8098: std_logic; attribute dont_touch of G8098: signal is true;
	signal G8099: std_logic; attribute dont_touch of G8099: signal is true;
	signal G8100: std_logic; attribute dont_touch of G8100: signal is true;
	signal G8101: std_logic; attribute dont_touch of G8101: signal is true;
	signal G8102: std_logic; attribute dont_touch of G8102: signal is true;
	signal G8103: std_logic; attribute dont_touch of G8103: signal is true;
	signal G8104: std_logic; attribute dont_touch of G8104: signal is true;
	signal G8105: std_logic; attribute dont_touch of G8105: signal is true;
	signal G8106: std_logic; attribute dont_touch of G8106: signal is true;
	signal G8107: std_logic; attribute dont_touch of G8107: signal is true;
	signal G8108: std_logic; attribute dont_touch of G8108: signal is true;
	signal G8109: std_logic; attribute dont_touch of G8109: signal is true;
	signal G8110: std_logic; attribute dont_touch of G8110: signal is true;
	signal G8115: std_logic; attribute dont_touch of G8115: signal is true;
	signal G8116: std_logic; attribute dont_touch of G8116: signal is true;
	signal G8117: std_logic; attribute dont_touch of G8117: signal is true;
	signal G8118: std_logic; attribute dont_touch of G8118: signal is true;
	signal G8119: std_logic; attribute dont_touch of G8119: signal is true;
	signal G8120: std_logic; attribute dont_touch of G8120: signal is true;
	signal G8121: std_logic; attribute dont_touch of G8121: signal is true;
	signal G8122: std_logic; attribute dont_touch of G8122: signal is true;
	signal G8123: std_logic; attribute dont_touch of G8123: signal is true;
	signal G8124: std_logic; attribute dont_touch of G8124: signal is true;
	signal G8125: std_logic; attribute dont_touch of G8125: signal is true;
	signal G8126: std_logic; attribute dont_touch of G8126: signal is true;
	signal G8127: std_logic; attribute dont_touch of G8127: signal is true;
	signal G8128: std_logic; attribute dont_touch of G8128: signal is true;
	signal G8129: std_logic; attribute dont_touch of G8129: signal is true;
	signal G8130: std_logic; attribute dont_touch of G8130: signal is true;
	signal G8131: std_logic; attribute dont_touch of G8131: signal is true;
	signal G8132: std_logic; attribute dont_touch of G8132: signal is true;
	signal G8133: std_logic; attribute dont_touch of G8133: signal is true;
	signal G8134: std_logic; attribute dont_touch of G8134: signal is true;
	signal G8135: std_logic; attribute dont_touch of G8135: signal is true;
	signal G8136: std_logic; attribute dont_touch of G8136: signal is true;
	signal G8137: std_logic; attribute dont_touch of G8137: signal is true;
	signal G8138: std_logic; attribute dont_touch of G8138: signal is true;
	signal G8139: std_logic; attribute dont_touch of G8139: signal is true;
	signal G8140: std_logic; attribute dont_touch of G8140: signal is true;
	signal G8141: std_logic; attribute dont_touch of G8141: signal is true;
	signal G8142: std_logic; attribute dont_touch of G8142: signal is true;
	signal G8143: std_logic; attribute dont_touch of G8143: signal is true;
	signal G8144: std_logic; attribute dont_touch of G8144: signal is true;
	signal G8145: std_logic; attribute dont_touch of G8145: signal is true;
	signal G8146: std_logic; attribute dont_touch of G8146: signal is true;
	signal G8147: std_logic; attribute dont_touch of G8147: signal is true;
	signal G8148: std_logic; attribute dont_touch of G8148: signal is true;
	signal G8149: std_logic; attribute dont_touch of G8149: signal is true;
	signal G8150: std_logic; attribute dont_touch of G8150: signal is true;
	signal G8151: std_logic; attribute dont_touch of G8151: signal is true;
	signal G8152: std_logic; attribute dont_touch of G8152: signal is true;
	signal G8153: std_logic; attribute dont_touch of G8153: signal is true;
	signal G8154: std_logic; attribute dont_touch of G8154: signal is true;
	signal G8155: std_logic; attribute dont_touch of G8155: signal is true;
	signal G8156: std_logic; attribute dont_touch of G8156: signal is true;
	signal G8157: std_logic; attribute dont_touch of G8157: signal is true;
	signal G8158: std_logic; attribute dont_touch of G8158: signal is true;
	signal G8159: std_logic; attribute dont_touch of G8159: signal is true;
	signal G8160: std_logic; attribute dont_touch of G8160: signal is true;
	signal G8161: std_logic; attribute dont_touch of G8161: signal is true;
	signal G8162: std_logic; attribute dont_touch of G8162: signal is true;
	signal G8163: std_logic; attribute dont_touch of G8163: signal is true;
	signal G8164: std_logic; attribute dont_touch of G8164: signal is true;
	signal G8167: std_logic; attribute dont_touch of G8167: signal is true;
	signal G8168: std_logic; attribute dont_touch of G8168: signal is true;
	signal G8169: std_logic; attribute dont_touch of G8169: signal is true;
	signal G8170: std_logic; attribute dont_touch of G8170: signal is true;
	signal G8171: std_logic; attribute dont_touch of G8171: signal is true;
	signal G8172: std_logic; attribute dont_touch of G8172: signal is true;
	signal G8173: std_logic; attribute dont_touch of G8173: signal is true;
	signal G8174: std_logic; attribute dont_touch of G8174: signal is true;
	signal G8175: std_logic; attribute dont_touch of G8175: signal is true;
	signal G8176: std_logic; attribute dont_touch of G8176: signal is true;
	signal G8177: std_logic; attribute dont_touch of G8177: signal is true;
	signal G8178: std_logic; attribute dont_touch of G8178: signal is true;
	signal G8179: std_logic; attribute dont_touch of G8179: signal is true;
	signal G8180: std_logic; attribute dont_touch of G8180: signal is true;
	signal G8181: std_logic; attribute dont_touch of G8181: signal is true;
	signal G8182: std_logic; attribute dont_touch of G8182: signal is true;
	signal G8183: std_logic; attribute dont_touch of G8183: signal is true;
	signal G8184: std_logic; attribute dont_touch of G8184: signal is true;
	signal G8185: std_logic; attribute dont_touch of G8185: signal is true;
	signal G8186: std_logic; attribute dont_touch of G8186: signal is true;
	signal G8187: std_logic; attribute dont_touch of G8187: signal is true;
	signal G8190: std_logic; attribute dont_touch of G8190: signal is true;
	signal G8191: std_logic; attribute dont_touch of G8191: signal is true;
	signal G8192: std_logic; attribute dont_touch of G8192: signal is true;
	signal G8193: std_logic; attribute dont_touch of G8193: signal is true;
	signal G8194: std_logic; attribute dont_touch of G8194: signal is true;
	signal G8195: std_logic; attribute dont_touch of G8195: signal is true;
	signal G8196: std_logic; attribute dont_touch of G8196: signal is true;
	signal G8197: std_logic; attribute dont_touch of G8197: signal is true;
	signal G8198: std_logic; attribute dont_touch of G8198: signal is true;
	signal G8199: std_logic; attribute dont_touch of G8199: signal is true;
	signal G8200: std_logic; attribute dont_touch of G8200: signal is true;
	signal G8203: std_logic; attribute dont_touch of G8203: signal is true;
	signal G8206: std_logic; attribute dont_touch of G8206: signal is true;
	signal G8209: std_logic; attribute dont_touch of G8209: signal is true;
	signal G8210: std_logic; attribute dont_touch of G8210: signal is true;
	signal G8213: std_logic; attribute dont_touch of G8213: signal is true;
	signal G8214: std_logic; attribute dont_touch of G8214: signal is true;
	signal G8217: std_logic; attribute dont_touch of G8217: signal is true;
	signal G8218: std_logic; attribute dont_touch of G8218: signal is true;
	signal G8219: std_logic; attribute dont_touch of G8219: signal is true;
	signal G8220: std_logic; attribute dont_touch of G8220: signal is true;
	signal G8221: std_logic; attribute dont_touch of G8221: signal is true;
	signal G8224: std_logic; attribute dont_touch of G8224: signal is true;
	signal G8225: std_logic; attribute dont_touch of G8225: signal is true;
	signal G8226: std_logic; attribute dont_touch of G8226: signal is true;
	signal G8229: std_logic; attribute dont_touch of G8229: signal is true;
	signal G8230: std_logic; attribute dont_touch of G8230: signal is true;
	signal G8233: std_logic; attribute dont_touch of G8233: signal is true;
	signal G8234: std_logic; attribute dont_touch of G8234: signal is true;
	signal G8235: std_logic; attribute dont_touch of G8235: signal is true;
	signal G8236: std_logic; attribute dont_touch of G8236: signal is true;
	signal G8239: std_logic; attribute dont_touch of G8239: signal is true;
	signal G8240: std_logic; attribute dont_touch of G8240: signal is true;
	signal G8241: std_logic; attribute dont_touch of G8241: signal is true;
	signal G8244: std_logic; attribute dont_touch of G8244: signal is true;
	signal G8245: std_logic; attribute dont_touch of G8245: signal is true;
	signal G8246: std_logic; attribute dont_touch of G8246: signal is true;
	signal G8247: std_logic; attribute dont_touch of G8247: signal is true;
	signal G8248: std_logic; attribute dont_touch of G8248: signal is true;
	signal G8249: std_logic; attribute dont_touch of G8249: signal is true;
	signal G8250: std_logic; attribute dont_touch of G8250: signal is true;
	signal G8251: std_logic; attribute dont_touch of G8251: signal is true;
	signal G8252: std_logic; attribute dont_touch of G8252: signal is true;
	signal G8253: std_logic; attribute dont_touch of G8253: signal is true;
	signal G8254: std_logic; attribute dont_touch of G8254: signal is true;
	signal G8255: std_logic; attribute dont_touch of G8255: signal is true;
	signal G8259: std_logic; attribute dont_touch of G8259: signal is true;
	signal G8260: std_logic; attribute dont_touch of G8260: signal is true;
	signal G8261: std_logic; attribute dont_touch of G8261: signal is true;
	signal G8262: std_logic; attribute dont_touch of G8262: signal is true;
	signal G8263: std_logic; attribute dont_touch of G8263: signal is true;
	signal G8264: std_logic; attribute dont_touch of G8264: signal is true;
	signal G8265: std_logic; attribute dont_touch of G8265: signal is true;
	signal G8266: std_logic; attribute dont_touch of G8266: signal is true;
	signal G8267: std_logic; attribute dont_touch of G8267: signal is true;
	signal G8268: std_logic; attribute dont_touch of G8268: signal is true;
	signal G8269: std_logic; attribute dont_touch of G8269: signal is true;
	signal G8270: std_logic; attribute dont_touch of G8270: signal is true;
	signal G8272: std_logic; attribute dont_touch of G8272: signal is true;
	signal G8273: std_logic; attribute dont_touch of G8273: signal is true;
	signal G8274: std_logic; attribute dont_touch of G8274: signal is true;
	signal G8275: std_logic; attribute dont_touch of G8275: signal is true;
	signal G8276: std_logic; attribute dont_touch of G8276: signal is true;
	signal G8277: std_logic; attribute dont_touch of G8277: signal is true;
	signal G8278: std_logic; attribute dont_touch of G8278: signal is true;
	signal G8279: std_logic; attribute dont_touch of G8279: signal is true;
	signal G8280: std_logic; attribute dont_touch of G8280: signal is true;
	signal G8281: std_logic; attribute dont_touch of G8281: signal is true;
	signal G8282: std_logic; attribute dont_touch of G8282: signal is true;
	signal G8283: std_logic; attribute dont_touch of G8283: signal is true;
	signal G8284: std_logic; attribute dont_touch of G8284: signal is true;
	signal G8285: std_logic; attribute dont_touch of G8285: signal is true;
	signal G8286: std_logic; attribute dont_touch of G8286: signal is true;
	signal G8287: std_logic; attribute dont_touch of G8287: signal is true;
	signal G8288: std_logic; attribute dont_touch of G8288: signal is true;
	signal G8289: std_logic; attribute dont_touch of G8289: signal is true;
	signal G8290: std_logic; attribute dont_touch of G8290: signal is true;
	signal G8291: std_logic; attribute dont_touch of G8291: signal is true;
	signal G8292: std_logic; attribute dont_touch of G8292: signal is true;
	signal G8293: std_logic; attribute dont_touch of G8293: signal is true;
	signal G8294: std_logic; attribute dont_touch of G8294: signal is true;
	signal G8295: std_logic; attribute dont_touch of G8295: signal is true;
	signal G8296: std_logic; attribute dont_touch of G8296: signal is true;
	signal G8297: std_logic; attribute dont_touch of G8297: signal is true;
	signal G8298: std_logic; attribute dont_touch of G8298: signal is true;
	signal G8299: std_logic; attribute dont_touch of G8299: signal is true;
	signal G8300: std_logic; attribute dont_touch of G8300: signal is true;
	signal G8301: std_logic; attribute dont_touch of G8301: signal is true;
	signal G8302: std_logic; attribute dont_touch of G8302: signal is true;
	signal G8303: std_logic; attribute dont_touch of G8303: signal is true;
	signal G8304: std_logic; attribute dont_touch of G8304: signal is true;
	signal G8305: std_logic; attribute dont_touch of G8305: signal is true;
	signal G8306: std_logic; attribute dont_touch of G8306: signal is true;
	signal G8307: std_logic; attribute dont_touch of G8307: signal is true;
	signal G8308: std_logic; attribute dont_touch of G8308: signal is true;
	signal G8309: std_logic; attribute dont_touch of G8309: signal is true;
	signal G8310: std_logic; attribute dont_touch of G8310: signal is true;
	signal G8311: std_logic; attribute dont_touch of G8311: signal is true;
	signal G8312: std_logic; attribute dont_touch of G8312: signal is true;
	signal G8314: std_logic; attribute dont_touch of G8314: signal is true;
	signal G8315: std_logic; attribute dont_touch of G8315: signal is true;
	signal G8317: std_logic; attribute dont_touch of G8317: signal is true;
	signal G8319: std_logic; attribute dont_touch of G8319: signal is true;
	signal G8320: std_logic; attribute dont_touch of G8320: signal is true;
	signal G8321: std_logic; attribute dont_touch of G8321: signal is true;
	signal G8322: std_logic; attribute dont_touch of G8322: signal is true;
	signal G8324: std_logic; attribute dont_touch of G8324: signal is true;
	signal G8325: std_logic; attribute dont_touch of G8325: signal is true;
	signal G8326: std_logic; attribute dont_touch of G8326: signal is true;
	signal G8327: std_logic; attribute dont_touch of G8327: signal is true;
	signal G8329: std_logic; attribute dont_touch of G8329: signal is true;
	signal G8330: std_logic; attribute dont_touch of G8330: signal is true;
	signal G8332: std_logic; attribute dont_touch of G8332: signal is true;
	signal G8333: std_logic; attribute dont_touch of G8333: signal is true;
	signal G8334: std_logic; attribute dont_touch of G8334: signal is true;
	signal G8336: std_logic; attribute dont_touch of G8336: signal is true;
	signal G8337: std_logic; attribute dont_touch of G8337: signal is true;
	signal G8338: std_logic; attribute dont_touch of G8338: signal is true;
	signal G8339: std_logic; attribute dont_touch of G8339: signal is true;
	signal G8341: std_logic; attribute dont_touch of G8341: signal is true;
	signal G8342: std_logic; attribute dont_touch of G8342: signal is true;
	signal G8343: std_logic; attribute dont_touch of G8343: signal is true;
	signal G8344: std_logic; attribute dont_touch of G8344: signal is true;
	signal G8345: std_logic; attribute dont_touch of G8345: signal is true;
	signal G8346: std_logic; attribute dont_touch of G8346: signal is true;
	signal G8348: std_logic; attribute dont_touch of G8348: signal is true;
	signal G8350: std_logic; attribute dont_touch of G8350: signal is true;
	signal G8351: std_logic; attribute dont_touch of G8351: signal is true;
	signal G8353: std_logic; attribute dont_touch of G8353: signal is true;
	signal G8354: std_logic; attribute dont_touch of G8354: signal is true;
	signal G8355: std_logic; attribute dont_touch of G8355: signal is true;
	signal G8356: std_logic; attribute dont_touch of G8356: signal is true;
	signal G8357: std_logic; attribute dont_touch of G8357: signal is true;
	signal G8358: std_logic; attribute dont_touch of G8358: signal is true;
	signal G8359: std_logic; attribute dont_touch of G8359: signal is true;
	signal G8360: std_logic; attribute dont_touch of G8360: signal is true;
	signal G8361: std_logic; attribute dont_touch of G8361: signal is true;
	signal G8362: std_logic; attribute dont_touch of G8362: signal is true;
	signal G8363: std_logic; attribute dont_touch of G8363: signal is true;
	signal G8364: std_logic; attribute dont_touch of G8364: signal is true;
	signal G8365: std_logic; attribute dont_touch of G8365: signal is true;
	signal G8366: std_logic; attribute dont_touch of G8366: signal is true;
	signal G8375: std_logic; attribute dont_touch of G8375: signal is true;
	signal G8376: std_logic; attribute dont_touch of G8376: signal is true;
	signal G8377: std_logic; attribute dont_touch of G8377: signal is true;
	signal G8378: std_logic; attribute dont_touch of G8378: signal is true;
	signal G8379: std_logic; attribute dont_touch of G8379: signal is true;
	signal G8380: std_logic; attribute dont_touch of G8380: signal is true;
	signal G8381: std_logic; attribute dont_touch of G8381: signal is true;
	signal G8382: std_logic; attribute dont_touch of G8382: signal is true;
	signal G8383: std_logic; attribute dont_touch of G8383: signal is true;
	signal G8384: std_logic; attribute dont_touch of G8384: signal is true;
	signal G8385: std_logic; attribute dont_touch of G8385: signal is true;
	signal G8386: std_logic; attribute dont_touch of G8386: signal is true;
	signal G8387: std_logic; attribute dont_touch of G8387: signal is true;
	signal G8388: std_logic; attribute dont_touch of G8388: signal is true;
	signal G8389: std_logic; attribute dont_touch of G8389: signal is true;
	signal G8390: std_logic; attribute dont_touch of G8390: signal is true;
	signal G8399: std_logic; attribute dont_touch of G8399: signal is true;
	signal G8400: std_logic; attribute dont_touch of G8400: signal is true;
	signal G8401: std_logic; attribute dont_touch of G8401: signal is true;
	signal G8402: std_logic; attribute dont_touch of G8402: signal is true;
	signal G8403: std_logic; attribute dont_touch of G8403: signal is true;
	signal G8404: std_logic; attribute dont_touch of G8404: signal is true;
	signal G8405: std_logic; attribute dont_touch of G8405: signal is true;
	signal G8406: std_logic; attribute dont_touch of G8406: signal is true;
	signal G8407: std_logic; attribute dont_touch of G8407: signal is true;
	signal G8408: std_logic; attribute dont_touch of G8408: signal is true;
	signal G8409: std_logic; attribute dont_touch of G8409: signal is true;
	signal G8410: std_logic; attribute dont_touch of G8410: signal is true;
	signal G8411: std_logic; attribute dont_touch of G8411: signal is true;
	signal G8412: std_logic; attribute dont_touch of G8412: signal is true;
	signal G8413: std_logic; attribute dont_touch of G8413: signal is true;
	signal G8414: std_logic; attribute dont_touch of G8414: signal is true;
	signal G8415: std_logic; attribute dont_touch of G8415: signal is true;
	signal G8416: std_logic; attribute dont_touch of G8416: signal is true;
	signal G8417: std_logic; attribute dont_touch of G8417: signal is true;
	signal G8418: std_logic; attribute dont_touch of G8418: signal is true;
	signal G8419: std_logic; attribute dont_touch of G8419: signal is true;
	signal G8420: std_logic; attribute dont_touch of G8420: signal is true;
	signal G8421: std_logic; attribute dont_touch of G8421: signal is true;
	signal G8422: std_logic; attribute dont_touch of G8422: signal is true;
	signal G8423: std_logic; attribute dont_touch of G8423: signal is true;
	signal G8424: std_logic; attribute dont_touch of G8424: signal is true;
	signal G8425: std_logic; attribute dont_touch of G8425: signal is true;
	signal G8426: std_logic; attribute dont_touch of G8426: signal is true;
	signal G8427: std_logic; attribute dont_touch of G8427: signal is true;
	signal G8428: std_logic; attribute dont_touch of G8428: signal is true;
	signal G8429: std_logic; attribute dont_touch of G8429: signal is true;
	signal G8430: std_logic; attribute dont_touch of G8430: signal is true;
	signal G8431: std_logic; attribute dont_touch of G8431: signal is true;
	signal G8432: std_logic; attribute dont_touch of G8432: signal is true;
	signal G8433: std_logic; attribute dont_touch of G8433: signal is true;
	signal G8434: std_logic; attribute dont_touch of G8434: signal is true;
	signal G8435: std_logic; attribute dont_touch of G8435: signal is true;
	signal G8436: std_logic; attribute dont_touch of G8436: signal is true;
	signal G8437: std_logic; attribute dont_touch of G8437: signal is true;
	signal G8438: std_logic; attribute dont_touch of G8438: signal is true;
	signal G8439: std_logic; attribute dont_touch of G8439: signal is true;
	signal G8440: std_logic; attribute dont_touch of G8440: signal is true;
	signal G8441: std_logic; attribute dont_touch of G8441: signal is true;
	signal G8442: std_logic; attribute dont_touch of G8442: signal is true;
	signal G8443: std_logic; attribute dont_touch of G8443: signal is true;
	signal G8444: std_logic; attribute dont_touch of G8444: signal is true;
	signal G8445: std_logic; attribute dont_touch of G8445: signal is true;
	signal G8446: std_logic; attribute dont_touch of G8446: signal is true;
	signal G8447: std_logic; attribute dont_touch of G8447: signal is true;
	signal G8448: std_logic; attribute dont_touch of G8448: signal is true;
	signal G8449: std_logic; attribute dont_touch of G8449: signal is true;
	signal G8450: std_logic; attribute dont_touch of G8450: signal is true;
	signal G8451: std_logic; attribute dont_touch of G8451: signal is true;
	signal G8461: std_logic; attribute dont_touch of G8461: signal is true;
	signal G8462: std_logic; attribute dont_touch of G8462: signal is true;
	signal G8463: std_logic; attribute dont_touch of G8463: signal is true;
	signal G8464: std_logic; attribute dont_touch of G8464: signal is true;
	signal G8465: std_logic; attribute dont_touch of G8465: signal is true;
	signal G8469: std_logic; attribute dont_touch of G8469: signal is true;
	signal G8470: std_logic; attribute dont_touch of G8470: signal is true;
	signal G8471: std_logic; attribute dont_touch of G8471: signal is true;
	signal G8472: std_logic; attribute dont_touch of G8472: signal is true;
	signal G8473: std_logic; attribute dont_touch of G8473: signal is true;
	signal G8474: std_logic; attribute dont_touch of G8474: signal is true;
	signal G8475: std_logic; attribute dont_touch of G8475: signal is true;
	signal G8476: std_logic; attribute dont_touch of G8476: signal is true;
	signal G8477: std_logic; attribute dont_touch of G8477: signal is true;
	signal G8478: std_logic; attribute dont_touch of G8478: signal is true;
	signal G8479: std_logic; attribute dont_touch of G8479: signal is true;
	signal G8480: std_logic; attribute dont_touch of G8480: signal is true;
	signal G8481: std_logic; attribute dont_touch of G8481: signal is true;
	signal G8482: std_logic; attribute dont_touch of G8482: signal is true;
	signal G8483: std_logic; attribute dont_touch of G8483: signal is true;
	signal G8484: std_logic; attribute dont_touch of G8484: signal is true;
	signal G8485: std_logic; attribute dont_touch of G8485: signal is true;
	signal G8486: std_logic; attribute dont_touch of G8486: signal is true;
	signal G8487: std_logic; attribute dont_touch of G8487: signal is true;
	signal G8488: std_logic; attribute dont_touch of G8488: signal is true;
	signal G8498: std_logic; attribute dont_touch of G8498: signal is true;
	signal G8499: std_logic; attribute dont_touch of G8499: signal is true;
	signal G8500: std_logic; attribute dont_touch of G8500: signal is true;
	signal G8501: std_logic; attribute dont_touch of G8501: signal is true;
	signal G8502: std_logic; attribute dont_touch of G8502: signal is true;
	signal G8505: std_logic; attribute dont_touch of G8505: signal is true;
	signal G8506: std_logic; attribute dont_touch of G8506: signal is true;
	signal G8507: std_logic; attribute dont_touch of G8507: signal is true;
	signal G8508: std_logic; attribute dont_touch of G8508: signal is true;
	signal G8509: std_logic; attribute dont_touch of G8509: signal is true;
	signal G8510: std_logic; attribute dont_touch of G8510: signal is true;
	signal G8511: std_logic; attribute dont_touch of G8511: signal is true;
	signal G8512: std_logic; attribute dont_touch of G8512: signal is true;
	signal G8513: std_logic; attribute dont_touch of G8513: signal is true;
	signal G8514: std_logic; attribute dont_touch of G8514: signal is true;
	signal G8515: std_logic; attribute dont_touch of G8515: signal is true;
	signal G8516: std_logic; attribute dont_touch of G8516: signal is true;
	signal G8517: std_logic; attribute dont_touch of G8517: signal is true;
	signal G8518: std_logic; attribute dont_touch of G8518: signal is true;
	signal G8519: std_logic; attribute dont_touch of G8519: signal is true;
	signal G8520: std_logic; attribute dont_touch of G8520: signal is true;
	signal G8523: std_logic; attribute dont_touch of G8523: signal is true;
	signal G8526: std_logic; attribute dont_touch of G8526: signal is true;
	signal G8529: std_logic; attribute dont_touch of G8529: signal is true;
	signal G8532: std_logic; attribute dont_touch of G8532: signal is true;
	signal G8535: std_logic; attribute dont_touch of G8535: signal is true;
	signal G8538: std_logic; attribute dont_touch of G8538: signal is true;
	signal G8541: std_logic; attribute dont_touch of G8541: signal is true;
	signal G8542: std_logic; attribute dont_touch of G8542: signal is true;
	signal G8545: std_logic; attribute dont_touch of G8545: signal is true;
	signal G8546: std_logic; attribute dont_touch of G8546: signal is true;
	signal G8547: std_logic; attribute dont_touch of G8547: signal is true;
	signal G8548: std_logic; attribute dont_touch of G8548: signal is true;
	signal G8549: std_logic; attribute dont_touch of G8549: signal is true;
	signal G8550: std_logic; attribute dont_touch of G8550: signal is true;
	signal G8551: std_logic; attribute dont_touch of G8551: signal is true;
	signal G8552: std_logic; attribute dont_touch of G8552: signal is true;
	signal G8553: std_logic; attribute dont_touch of G8553: signal is true;
	signal G8554: std_logic; attribute dont_touch of G8554: signal is true;
	signal G8555: std_logic; attribute dont_touch of G8555: signal is true;
	signal G8556: std_logic; attribute dont_touch of G8556: signal is true;
	signal G8557: std_logic; attribute dont_touch of G8557: signal is true;
	signal G8558: std_logic; attribute dont_touch of G8558: signal is true;
	signal G8559: std_logic; attribute dont_touch of G8559: signal is true;
	signal G8560: std_logic; attribute dont_touch of G8560: signal is true;
	signal G8567: std_logic; attribute dont_touch of G8567: signal is true;
	signal G8568: std_logic; attribute dont_touch of G8568: signal is true;
	signal G8569: std_logic; attribute dont_touch of G8569: signal is true;
	signal G8570: std_logic; attribute dont_touch of G8570: signal is true;
	signal G8571: std_logic; attribute dont_touch of G8571: signal is true;
	signal G8572: std_logic; attribute dont_touch of G8572: signal is true;
	signal G8573: std_logic; attribute dont_touch of G8573: signal is true;
	signal G8574: std_logic; attribute dont_touch of G8574: signal is true;
	signal G8575: std_logic; attribute dont_touch of G8575: signal is true;
	signal G8576: std_logic; attribute dont_touch of G8576: signal is true;
	signal G8579: std_logic; attribute dont_touch of G8579: signal is true;
	signal G8582: std_logic; attribute dont_touch of G8582: signal is true;
	signal G8585: std_logic; attribute dont_touch of G8585: signal is true;
	signal G8588: std_logic; attribute dont_touch of G8588: signal is true;
	signal G8589: std_logic; attribute dont_touch of G8589: signal is true;
	signal G8592: std_logic; attribute dont_touch of G8592: signal is true;
	signal G8595: std_logic; attribute dont_touch of G8595: signal is true;
	signal G8598: std_logic; attribute dont_touch of G8598: signal is true;
	signal G8599: std_logic; attribute dont_touch of G8599: signal is true;
	signal G8600: std_logic; attribute dont_touch of G8600: signal is true;
	signal G8601: std_logic; attribute dont_touch of G8601: signal is true;
	signal G8602: std_logic; attribute dont_touch of G8602: signal is true;
	signal G8603: std_logic; attribute dont_touch of G8603: signal is true;
	signal G8604: std_logic; attribute dont_touch of G8604: signal is true;
	signal G8605: std_logic; attribute dont_touch of G8605: signal is true;
	signal G8606: std_logic; attribute dont_touch of G8606: signal is true;
	signal G8607: std_logic; attribute dont_touch of G8607: signal is true;
	signal G8608: std_logic; attribute dont_touch of G8608: signal is true;
	signal G8609: std_logic; attribute dont_touch of G8609: signal is true;
	signal G8610: std_logic; attribute dont_touch of G8610: signal is true;
	signal G8611: std_logic; attribute dont_touch of G8611: signal is true;
	signal G8612: std_logic; attribute dont_touch of G8612: signal is true;
	signal G8613: std_logic; attribute dont_touch of G8613: signal is true;
	signal G8614: std_logic; attribute dont_touch of G8614: signal is true;
	signal G8615: std_logic; attribute dont_touch of G8615: signal is true;
	signal G8616: std_logic; attribute dont_touch of G8616: signal is true;
	signal G8617: std_logic; attribute dont_touch of G8617: signal is true;
	signal G8622: std_logic; attribute dont_touch of G8622: signal is true;
	signal G8623: std_logic; attribute dont_touch of G8623: signal is true;
	signal G8624: std_logic; attribute dont_touch of G8624: signal is true;
	signal G8625: std_logic; attribute dont_touch of G8625: signal is true;
	signal G8626: std_logic; attribute dont_touch of G8626: signal is true;
	signal G8627: std_logic; attribute dont_touch of G8627: signal is true;
	signal G8628: std_logic; attribute dont_touch of G8628: signal is true;
	signal G8629: std_logic; attribute dont_touch of G8629: signal is true;
	signal G8630: std_logic; attribute dont_touch of G8630: signal is true;
	signal G8631: std_logic; attribute dont_touch of G8631: signal is true;
	signal G8632: std_logic; attribute dont_touch of G8632: signal is true;
	signal G8635: std_logic; attribute dont_touch of G8635: signal is true;
	signal G8638: std_logic; attribute dont_touch of G8638: signal is true;
	signal G8639: std_logic; attribute dont_touch of G8639: signal is true;
	signal G8640: std_logic; attribute dont_touch of G8640: signal is true;
	signal G8641: std_logic; attribute dont_touch of G8641: signal is true;
	signal G8642: std_logic; attribute dont_touch of G8642: signal is true;
	signal G8643: std_logic; attribute dont_touch of G8643: signal is true;
	signal G8644: std_logic; attribute dont_touch of G8644: signal is true;
	signal G8645: std_logic; attribute dont_touch of G8645: signal is true;
	signal G8646: std_logic; attribute dont_touch of G8646: signal is true;
	signal G8647: std_logic; attribute dont_touch of G8647: signal is true;
	signal G8648: std_logic; attribute dont_touch of G8648: signal is true;
	signal G8649: std_logic; attribute dont_touch of G8649: signal is true;
	signal G8650: std_logic; attribute dont_touch of G8650: signal is true;
	signal G8651: std_logic; attribute dont_touch of G8651: signal is true;
	signal G8652: std_logic; attribute dont_touch of G8652: signal is true;
	signal G8653: std_logic; attribute dont_touch of G8653: signal is true;
	signal G8654: std_logic; attribute dont_touch of G8654: signal is true;
	signal G8655: std_logic; attribute dont_touch of G8655: signal is true;
	signal G8656: std_logic; attribute dont_touch of G8656: signal is true;
	signal G8659: std_logic; attribute dont_touch of G8659: signal is true;
	signal G8660: std_logic; attribute dont_touch of G8660: signal is true;
	signal G8663: std_logic; attribute dont_touch of G8663: signal is true;
	signal G8664: std_logic; attribute dont_touch of G8664: signal is true;
	signal G8667: std_logic; attribute dont_touch of G8667: signal is true;
	signal G8670: std_logic; attribute dont_touch of G8670: signal is true;
	signal G8671: std_logic; attribute dont_touch of G8671: signal is true;
	signal G8674: std_logic; attribute dont_touch of G8674: signal is true;
	signal G8677: std_logic; attribute dont_touch of G8677: signal is true;
	signal G8680: std_logic; attribute dont_touch of G8680: signal is true;
	signal G8683: std_logic; attribute dont_touch of G8683: signal is true;
	signal G8684: std_logic; attribute dont_touch of G8684: signal is true;
	signal G8687: std_logic; attribute dont_touch of G8687: signal is true;
	signal G8688: std_logic; attribute dont_touch of G8688: signal is true;
	signal G8693: std_logic; attribute dont_touch of G8693: signal is true;
	signal G8694: std_logic; attribute dont_touch of G8694: signal is true;
	signal G8695: std_logic; attribute dont_touch of G8695: signal is true;
	signal G8696: std_logic; attribute dont_touch of G8696: signal is true;
	signal G8697: std_logic; attribute dont_touch of G8697: signal is true;
	signal G8698: std_logic; attribute dont_touch of G8698: signal is true;
	signal G8699: std_logic; attribute dont_touch of G8699: signal is true;
	signal G8700: std_logic; attribute dont_touch of G8700: signal is true;
	signal G8701: std_logic; attribute dont_touch of G8701: signal is true;
	signal G8702: std_logic; attribute dont_touch of G8702: signal is true;
	signal G8703: std_logic; attribute dont_touch of G8703: signal is true;
	signal G8704: std_logic; attribute dont_touch of G8704: signal is true;
	signal G8705: std_logic; attribute dont_touch of G8705: signal is true;
	signal G8706: std_logic; attribute dont_touch of G8706: signal is true;
	signal G8707: std_logic; attribute dont_touch of G8707: signal is true;
	signal G8708: std_logic; attribute dont_touch of G8708: signal is true;
	signal G8709: std_logic; attribute dont_touch of G8709: signal is true;
	signal G8710: std_logic; attribute dont_touch of G8710: signal is true;
	signal G8711: std_logic; attribute dont_touch of G8711: signal is true;
	signal G8712: std_logic; attribute dont_touch of G8712: signal is true;
	signal G8713: std_logic; attribute dont_touch of G8713: signal is true;
	signal G8714: std_logic; attribute dont_touch of G8714: signal is true;
	signal G8715: std_logic; attribute dont_touch of G8715: signal is true;
	signal G8716: std_logic; attribute dont_touch of G8716: signal is true;
	signal G8717: std_logic; attribute dont_touch of G8717: signal is true;
	signal G8718: std_logic; attribute dont_touch of G8718: signal is true;
	signal G8719: std_logic; attribute dont_touch of G8719: signal is true;
	signal G8720: std_logic; attribute dont_touch of G8720: signal is true;
	signal G8721: std_logic; attribute dont_touch of G8721: signal is true;
	signal G8722: std_logic; attribute dont_touch of G8722: signal is true;
	signal G8723: std_logic; attribute dont_touch of G8723: signal is true;
	signal G8724: std_logic; attribute dont_touch of G8724: signal is true;
	signal G8725: std_logic; attribute dont_touch of G8725: signal is true;
	signal G8726: std_logic; attribute dont_touch of G8726: signal is true;
	signal G8727: std_logic; attribute dont_touch of G8727: signal is true;
	signal G8728: std_logic; attribute dont_touch of G8728: signal is true;
	signal G8729: std_logic; attribute dont_touch of G8729: signal is true;
	signal G8730: std_logic; attribute dont_touch of G8730: signal is true;
	signal G8731: std_logic; attribute dont_touch of G8731: signal is true;
	signal G8732: std_logic; attribute dont_touch of G8732: signal is true;
	signal G8733: std_logic; attribute dont_touch of G8733: signal is true;
	signal G8734: std_logic; attribute dont_touch of G8734: signal is true;
	signal G8735: std_logic; attribute dont_touch of G8735: signal is true;
	signal G8736: std_logic; attribute dont_touch of G8736: signal is true;
	signal G8737: std_logic; attribute dont_touch of G8737: signal is true;
	signal G8738: std_logic; attribute dont_touch of G8738: signal is true;
	signal G8739: std_logic; attribute dont_touch of G8739: signal is true;
	signal G8742: std_logic; attribute dont_touch of G8742: signal is true;
	signal G8743: std_logic; attribute dont_touch of G8743: signal is true;
	signal G8744: std_logic; attribute dont_touch of G8744: signal is true;
	signal G8745: std_logic; attribute dont_touch of G8745: signal is true;
	signal G8746: std_logic; attribute dont_touch of G8746: signal is true;
	signal G8747: std_logic; attribute dont_touch of G8747: signal is true;
	signal G8748: std_logic; attribute dont_touch of G8748: signal is true;
	signal G8749: std_logic; attribute dont_touch of G8749: signal is true;
	signal G8750: std_logic; attribute dont_touch of G8750: signal is true;
	signal G8751: std_logic; attribute dont_touch of G8751: signal is true;
	signal G8752: std_logic; attribute dont_touch of G8752: signal is true;
	signal G8753: std_logic; attribute dont_touch of G8753: signal is true;
	signal G8754: std_logic; attribute dont_touch of G8754: signal is true;
	signal G8755: std_logic; attribute dont_touch of G8755: signal is true;
	signal G8756: std_logic; attribute dont_touch of G8756: signal is true;
	signal G8757: std_logic; attribute dont_touch of G8757: signal is true;
	signal G8758: std_logic; attribute dont_touch of G8758: signal is true;
	signal G8759: std_logic; attribute dont_touch of G8759: signal is true;
	signal G8760: std_logic; attribute dont_touch of G8760: signal is true;
	signal G8763: std_logic; attribute dont_touch of G8763: signal is true;
	signal G8764: std_logic; attribute dont_touch of G8764: signal is true;
	signal G8765: std_logic; attribute dont_touch of G8765: signal is true;
	signal G8766: std_logic; attribute dont_touch of G8766: signal is true;
	signal G8767: std_logic; attribute dont_touch of G8767: signal is true;
	signal G8768: std_logic; attribute dont_touch of G8768: signal is true;
	signal G8769: std_logic; attribute dont_touch of G8769: signal is true;
	signal G8770: std_logic; attribute dont_touch of G8770: signal is true;
	signal G8771: std_logic; attribute dont_touch of G8771: signal is true;
	signal G8772: std_logic; attribute dont_touch of G8772: signal is true;
	signal G8773: std_logic; attribute dont_touch of G8773: signal is true;
	signal G8774: std_logic; attribute dont_touch of G8774: signal is true;
	signal G8775: std_logic; attribute dont_touch of G8775: signal is true;
	signal G8776: std_logic; attribute dont_touch of G8776: signal is true;
	signal G8777: std_logic; attribute dont_touch of G8777: signal is true;
	signal G8778: std_logic; attribute dont_touch of G8778: signal is true;
	signal G8779: std_logic; attribute dont_touch of G8779: signal is true;
	signal G8780: std_logic; attribute dont_touch of G8780: signal is true;
	signal G8781: std_logic; attribute dont_touch of G8781: signal is true;
	signal G8782: std_logic; attribute dont_touch of G8782: signal is true;
	signal G8783: std_logic; attribute dont_touch of G8783: signal is true;
	signal G8784: std_logic; attribute dont_touch of G8784: signal is true;
	signal G8785: std_logic; attribute dont_touch of G8785: signal is true;
	signal G8786: std_logic; attribute dont_touch of G8786: signal is true;
	signal G8787: std_logic; attribute dont_touch of G8787: signal is true;
	signal G8788: std_logic; attribute dont_touch of G8788: signal is true;
	signal G8789: std_logic; attribute dont_touch of G8789: signal is true;
	signal G8790: std_logic; attribute dont_touch of G8790: signal is true;
	signal G8791: std_logic; attribute dont_touch of G8791: signal is true;
	signal G8792: std_logic; attribute dont_touch of G8792: signal is true;
	signal G8793: std_logic; attribute dont_touch of G8793: signal is true;
	signal G8794: std_logic; attribute dont_touch of G8794: signal is true;
	signal G8795: std_logic; attribute dont_touch of G8795: signal is true;
	signal G8796: std_logic; attribute dont_touch of G8796: signal is true;
	signal G8797: std_logic; attribute dont_touch of G8797: signal is true;
	signal G8798: std_logic; attribute dont_touch of G8798: signal is true;
	signal G8799: std_logic; attribute dont_touch of G8799: signal is true;
	signal G8800: std_logic; attribute dont_touch of G8800: signal is true;
	signal G8801: std_logic; attribute dont_touch of G8801: signal is true;
	signal G8802: std_logic; attribute dont_touch of G8802: signal is true;
	signal G8803: std_logic; attribute dont_touch of G8803: signal is true;
	signal G8804: std_logic; attribute dont_touch of G8804: signal is true;
	signal G8805: std_logic; attribute dont_touch of G8805: signal is true;
	signal G8806: std_logic; attribute dont_touch of G8806: signal is true;
	signal G8807: std_logic; attribute dont_touch of G8807: signal is true;
	signal G8810: std_logic; attribute dont_touch of G8810: signal is true;
	signal G8811: std_logic; attribute dont_touch of G8811: signal is true;
	signal G8812: std_logic; attribute dont_touch of G8812: signal is true;
	signal G8813: std_logic; attribute dont_touch of G8813: signal is true;
	signal G8814: std_logic; attribute dont_touch of G8814: signal is true;
	signal G8815: std_logic; attribute dont_touch of G8815: signal is true;
	signal G8816: std_logic; attribute dont_touch of G8816: signal is true;
	signal G8817: std_logic; attribute dont_touch of G8817: signal is true;
	signal G8818: std_logic; attribute dont_touch of G8818: signal is true;
	signal G8819: std_logic; attribute dont_touch of G8819: signal is true;
	signal G8820: std_logic; attribute dont_touch of G8820: signal is true;
	signal G8821: std_logic; attribute dont_touch of G8821: signal is true;
	signal G8822: std_logic; attribute dont_touch of G8822: signal is true;
	signal G8823: std_logic; attribute dont_touch of G8823: signal is true;
	signal G8824: std_logic; attribute dont_touch of G8824: signal is true;
	signal G8825: std_logic; attribute dont_touch of G8825: signal is true;
	signal G8826: std_logic; attribute dont_touch of G8826: signal is true;
	signal G8827: std_logic; attribute dont_touch of G8827: signal is true;
	signal G8828: std_logic; attribute dont_touch of G8828: signal is true;
	signal G8837: std_logic; attribute dont_touch of G8837: signal is true;
	signal G8838: std_logic; attribute dont_touch of G8838: signal is true;
	signal G8839: std_logic; attribute dont_touch of G8839: signal is true;
	signal G8840: std_logic; attribute dont_touch of G8840: signal is true;
	signal G8841: std_logic; attribute dont_touch of G8841: signal is true;
	signal G8842: std_logic; attribute dont_touch of G8842: signal is true;
	signal G8843: std_logic; attribute dont_touch of G8843: signal is true;
	signal G8844: std_logic; attribute dont_touch of G8844: signal is true;
	signal G8845: std_logic; attribute dont_touch of G8845: signal is true;
	signal G8846: std_logic; attribute dont_touch of G8846: signal is true;
	signal G8847: std_logic; attribute dont_touch of G8847: signal is true;
	signal G8848: std_logic; attribute dont_touch of G8848: signal is true;
	signal G8849: std_logic; attribute dont_touch of G8849: signal is true;
	signal G8858: std_logic; attribute dont_touch of G8858: signal is true;
	signal G8868: std_logic; attribute dont_touch of G8868: signal is true;
	signal G8869: std_logic; attribute dont_touch of G8869: signal is true;
	signal G8870: std_logic; attribute dont_touch of G8870: signal is true;
	signal G8871: std_logic; attribute dont_touch of G8871: signal is true;
	signal G8872: std_logic; attribute dont_touch of G8872: signal is true;
	signal G8873: std_logic; attribute dont_touch of G8873: signal is true;
	signal G8874: std_logic; attribute dont_touch of G8874: signal is true;
	signal G8875: std_logic; attribute dont_touch of G8875: signal is true;
	signal G8876: std_logic; attribute dont_touch of G8876: signal is true;
	signal G8877: std_logic; attribute dont_touch of G8877: signal is true;
	signal G8878: std_logic; attribute dont_touch of G8878: signal is true;
	signal G8879: std_logic; attribute dont_touch of G8879: signal is true;
	signal G8880: std_logic; attribute dont_touch of G8880: signal is true;
	signal G8881: std_logic; attribute dont_touch of G8881: signal is true;
	signal G8882: std_logic; attribute dont_touch of G8882: signal is true;
	signal G8883: std_logic; attribute dont_touch of G8883: signal is true;
	signal G8884: std_logic; attribute dont_touch of G8884: signal is true;
	signal G8885: std_logic; attribute dont_touch of G8885: signal is true;
	signal G8886: std_logic; attribute dont_touch of G8886: signal is true;
	signal G8887: std_logic; attribute dont_touch of G8887: signal is true;
	signal G8888: std_logic; attribute dont_touch of G8888: signal is true;
	signal G8889: std_logic; attribute dont_touch of G8889: signal is true;
	signal G8890: std_logic; attribute dont_touch of G8890: signal is true;
	signal G8891: std_logic; attribute dont_touch of G8891: signal is true;
	signal G8892: std_logic; attribute dont_touch of G8892: signal is true;
	signal G8920: std_logic; attribute dont_touch of G8920: signal is true;
	signal G8921: std_logic; attribute dont_touch of G8921: signal is true;
	signal G8922: std_logic; attribute dont_touch of G8922: signal is true;
	signal G8923: std_logic; attribute dont_touch of G8923: signal is true;
	signal G8924: std_logic; attribute dont_touch of G8924: signal is true;
	signal G8925: std_logic; attribute dont_touch of G8925: signal is true;
	signal G8926: std_logic; attribute dont_touch of G8926: signal is true;
	signal G8927: std_logic; attribute dont_touch of G8927: signal is true;
	signal G8928: std_logic; attribute dont_touch of G8928: signal is true;
	signal G8929: std_logic; attribute dont_touch of G8929: signal is true;
	signal G8930: std_logic; attribute dont_touch of G8930: signal is true;
	signal G8931: std_logic; attribute dont_touch of G8931: signal is true;
	signal G8932: std_logic; attribute dont_touch of G8932: signal is true;
	signal G8933: std_logic; attribute dont_touch of G8933: signal is true;
	signal G8934: std_logic; attribute dont_touch of G8934: signal is true;
	signal G8935: std_logic; attribute dont_touch of G8935: signal is true;
	signal G8936: std_logic; attribute dont_touch of G8936: signal is true;
	signal G8937: std_logic; attribute dont_touch of G8937: signal is true;
	signal G8938: std_logic; attribute dont_touch of G8938: signal is true;
	signal G8939: std_logic; attribute dont_touch of G8939: signal is true;
	signal G8940: std_logic; attribute dont_touch of G8940: signal is true;
	signal G8941: std_logic; attribute dont_touch of G8941: signal is true;
	signal G8942: std_logic; attribute dont_touch of G8942: signal is true;
	signal G8943: std_logic; attribute dont_touch of G8943: signal is true;
	signal G8944: std_logic; attribute dont_touch of G8944: signal is true;
	signal G8945: std_logic; attribute dont_touch of G8945: signal is true;
	signal G8946: std_logic; attribute dont_touch of G8946: signal is true;
	signal G8947: std_logic; attribute dont_touch of G8947: signal is true;
	signal G8948: std_logic; attribute dont_touch of G8948: signal is true;
	signal G8949: std_logic; attribute dont_touch of G8949: signal is true;
	signal G8950: std_logic; attribute dont_touch of G8950: signal is true;
	signal G8951: std_logic; attribute dont_touch of G8951: signal is true;
	signal G8952: std_logic; attribute dont_touch of G8952: signal is true;
	signal G8953: std_logic; attribute dont_touch of G8953: signal is true;
	signal G8954: std_logic; attribute dont_touch of G8954: signal is true;
	signal G8955: std_logic; attribute dont_touch of G8955: signal is true;
	signal G8956: std_logic; attribute dont_touch of G8956: signal is true;
	signal G8957: std_logic; attribute dont_touch of G8957: signal is true;
	signal G8958: std_logic; attribute dont_touch of G8958: signal is true;
	signal G8959: std_logic; attribute dont_touch of G8959: signal is true;
	signal G8960: std_logic; attribute dont_touch of G8960: signal is true;
	signal G8961: std_logic; attribute dont_touch of G8961: signal is true;
	signal G8962: std_logic; attribute dont_touch of G8962: signal is true;
	signal G8963: std_logic; attribute dont_touch of G8963: signal is true;
	signal G8964: std_logic; attribute dont_touch of G8964: signal is true;
	signal G8965: std_logic; attribute dont_touch of G8965: signal is true;
	signal G8966: std_logic; attribute dont_touch of G8966: signal is true;
	signal G8967: std_logic; attribute dont_touch of G8967: signal is true;
	signal G8968: std_logic; attribute dont_touch of G8968: signal is true;
	signal G8969: std_logic; attribute dont_touch of G8969: signal is true;
	signal G8970: std_logic; attribute dont_touch of G8970: signal is true;
	signal G8971: std_logic; attribute dont_touch of G8971: signal is true;
	signal G8972: std_logic; attribute dont_touch of G8972: signal is true;
	signal G8973: std_logic; attribute dont_touch of G8973: signal is true;
	signal G8974: std_logic; attribute dont_touch of G8974: signal is true;
	signal G8975: std_logic; attribute dont_touch of G8975: signal is true;
	signal G8987: std_logic; attribute dont_touch of G8987: signal is true;
	signal G8988: std_logic; attribute dont_touch of G8988: signal is true;
	signal G8989: std_logic; attribute dont_touch of G8989: signal is true;
	signal G8990: std_logic; attribute dont_touch of G8990: signal is true;
	signal G8991: std_logic; attribute dont_touch of G8991: signal is true;
	signal G8992: std_logic; attribute dont_touch of G8992: signal is true;
	signal G8993: std_logic; attribute dont_touch of G8993: signal is true;
	signal G8994: std_logic; attribute dont_touch of G8994: signal is true;
	signal G8995: std_logic; attribute dont_touch of G8995: signal is true;
	signal G9009: std_logic; attribute dont_touch of G9009: signal is true;
	signal G9010: std_logic; attribute dont_touch of G9010: signal is true;
	signal G9024: std_logic; attribute dont_touch of G9024: signal is true;
	signal G9025: std_logic; attribute dont_touch of G9025: signal is true;
	signal G9026: std_logic; attribute dont_touch of G9026: signal is true;
	signal G9027: std_logic; attribute dont_touch of G9027: signal is true;
	signal G9028: std_logic; attribute dont_touch of G9028: signal is true;
	signal G9029: std_logic; attribute dont_touch of G9029: signal is true;
	signal G9030: std_logic; attribute dont_touch of G9030: signal is true;
	signal G9052: std_logic; attribute dont_touch of G9052: signal is true;
	signal G9076: std_logic; attribute dont_touch of G9076: signal is true;
	signal G9079: std_logic; attribute dont_touch of G9079: signal is true;
	signal G9082: std_logic; attribute dont_touch of G9082: signal is true;
	signal G9085: std_logic; attribute dont_touch of G9085: signal is true;
	signal G9088: std_logic; attribute dont_touch of G9088: signal is true;
	signal G9091: std_logic; attribute dont_touch of G9091: signal is true;
	signal G9094: std_logic; attribute dont_touch of G9094: signal is true;
	signal G9097: std_logic; attribute dont_touch of G9097: signal is true;
	signal G9100: std_logic; attribute dont_touch of G9100: signal is true;
	signal G9103: std_logic; attribute dont_touch of G9103: signal is true;
	signal G9106: std_logic; attribute dont_touch of G9106: signal is true;
	signal G9107: std_logic; attribute dont_touch of G9107: signal is true;
	signal G9108: std_logic; attribute dont_touch of G9108: signal is true;
	signal G9109: std_logic; attribute dont_touch of G9109: signal is true;
	signal G9110: std_logic; attribute dont_touch of G9110: signal is true;
	signal G9111: std_logic; attribute dont_touch of G9111: signal is true;
	signal G9124: std_logic; attribute dont_touch of G9124: signal is true;
	signal G9125: std_logic; attribute dont_touch of G9125: signal is true;
	signal G9150: std_logic; attribute dont_touch of G9150: signal is true;
	signal G9151: std_logic; attribute dont_touch of G9151: signal is true;
	signal G9173: std_logic; attribute dont_touch of G9173: signal is true;
	signal G9192: std_logic; attribute dont_touch of G9192: signal is true;
	signal G9204: std_logic; attribute dont_touch of G9204: signal is true;
	signal G9205: std_logic; attribute dont_touch of G9205: signal is true;
	signal G9223: std_logic; attribute dont_touch of G9223: signal is true;
	signal G9240: std_logic; attribute dont_touch of G9240: signal is true;
	signal G9256: std_logic; attribute dont_touch of G9256: signal is true;
	signal G9257: std_logic; attribute dont_touch of G9257: signal is true;
	signal G9258: std_logic; attribute dont_touch of G9258: signal is true;
	signal G9259: std_logic; attribute dont_touch of G9259: signal is true;
	signal G9260: std_logic; attribute dont_touch of G9260: signal is true;
	signal G9261: std_logic; attribute dont_touch of G9261: signal is true;
	signal G9262: std_logic; attribute dont_touch of G9262: signal is true;
	signal G9263: std_logic; attribute dont_touch of G9263: signal is true;
	signal G9264: std_logic; attribute dont_touch of G9264: signal is true;
	signal G9265: std_logic; attribute dont_touch of G9265: signal is true;
	signal G9266: std_logic; attribute dont_touch of G9266: signal is true;
	signal G9267: std_logic; attribute dont_touch of G9267: signal is true;
	signal G9268: std_logic; attribute dont_touch of G9268: signal is true;
	signal G9269: std_logic; attribute dont_touch of G9269: signal is true;
	signal G9270: std_logic; attribute dont_touch of G9270: signal is true;
	signal G9271: std_logic; attribute dont_touch of G9271: signal is true;
	signal G9272: std_logic; attribute dont_touch of G9272: signal is true;
	signal G9273: std_logic; attribute dont_touch of G9273: signal is true;
	signal G9274: std_logic; attribute dont_touch of G9274: signal is true;
	signal G9290: std_logic; attribute dont_touch of G9290: signal is true;
	signal G9291: std_logic; attribute dont_touch of G9291: signal is true;
	signal G9292: std_logic; attribute dont_touch of G9292: signal is true;
	signal G9308: std_logic; attribute dont_touch of G9308: signal is true;
	signal G9309: std_logic; attribute dont_touch of G9309: signal is true;
	signal G9310: std_logic; attribute dont_touch of G9310: signal is true;
	signal G9311: std_logic; attribute dont_touch of G9311: signal is true;
	signal G9312: std_logic; attribute dont_touch of G9312: signal is true;
	signal G9313: std_logic; attribute dont_touch of G9313: signal is true;
	signal G9316: std_logic; attribute dont_touch of G9316: signal is true;
	signal G9317: std_logic; attribute dont_touch of G9317: signal is true;
	signal G9324: std_logic; attribute dont_touch of G9324: signal is true;
	signal G9328: std_logic; attribute dont_touch of G9328: signal is true;
	signal G9331: std_logic; attribute dont_touch of G9331: signal is true;
	signal G9335: std_logic; attribute dont_touch of G9335: signal is true;
	signal G9338: std_logic; attribute dont_touch of G9338: signal is true;
	signal G9339: std_logic; attribute dont_touch of G9339: signal is true;
	signal G9340: std_logic; attribute dont_touch of G9340: signal is true;
	signal G9341: std_logic; attribute dont_touch of G9341: signal is true;
	signal G9342: std_logic; attribute dont_touch of G9342: signal is true;
	signal G9343: std_logic; attribute dont_touch of G9343: signal is true;
	signal G9344: std_logic; attribute dont_touch of G9344: signal is true;
	signal G9345: std_logic; attribute dont_touch of G9345: signal is true;
	signal G9346: std_logic; attribute dont_touch of G9346: signal is true;
	signal G9347: std_logic; attribute dont_touch of G9347: signal is true;
	signal G9348: std_logic; attribute dont_touch of G9348: signal is true;
	signal G9349: std_logic; attribute dont_touch of G9349: signal is true;
	signal G9350: std_logic; attribute dont_touch of G9350: signal is true;
	signal G9351: std_logic; attribute dont_touch of G9351: signal is true;
	signal G9352: std_logic; attribute dont_touch of G9352: signal is true;
	signal G9353: std_logic; attribute dont_touch of G9353: signal is true;
	signal G9354: std_logic; attribute dont_touch of G9354: signal is true;
	signal G9355: std_logic; attribute dont_touch of G9355: signal is true;
	signal G9356: std_logic; attribute dont_touch of G9356: signal is true;
	signal G9357: std_logic; attribute dont_touch of G9357: signal is true;
	signal G9358: std_logic; attribute dont_touch of G9358: signal is true;
	signal G9359: std_logic; attribute dont_touch of G9359: signal is true;
	signal G9360: std_logic; attribute dont_touch of G9360: signal is true;
	signal G9361: std_logic; attribute dont_touch of G9361: signal is true;
	signal G9362: std_logic; attribute dont_touch of G9362: signal is true;
	signal G9363: std_logic; attribute dont_touch of G9363: signal is true;
	signal G9364: std_logic; attribute dont_touch of G9364: signal is true;
	signal G9365: std_logic; attribute dont_touch of G9365: signal is true;
	signal G9366: std_logic; attribute dont_touch of G9366: signal is true;
	signal G9367: std_logic; attribute dont_touch of G9367: signal is true;
	signal G9384: std_logic; attribute dont_touch of G9384: signal is true;
	signal G9385: std_logic; attribute dont_touch of G9385: signal is true;
	signal G9386: std_logic; attribute dont_touch of G9386: signal is true;
	signal G9387: std_logic; attribute dont_touch of G9387: signal is true;
	signal G9388: std_logic; attribute dont_touch of G9388: signal is true;
	signal G9389: std_logic; attribute dont_touch of G9389: signal is true;
	signal G9390: std_logic; attribute dont_touch of G9390: signal is true;
	signal G9391: std_logic; attribute dont_touch of G9391: signal is true;
	signal G9392: std_logic; attribute dont_touch of G9392: signal is true;
	signal G9409: std_logic; attribute dont_touch of G9409: signal is true;
	signal G9410: std_logic; attribute dont_touch of G9410: signal is true;
	signal G9411: std_logic; attribute dont_touch of G9411: signal is true;
	signal G9412: std_logic; attribute dont_touch of G9412: signal is true;
	signal G9413: std_logic; attribute dont_touch of G9413: signal is true;
	signal G9414: std_logic; attribute dont_touch of G9414: signal is true;
	signal G9415: std_logic; attribute dont_touch of G9415: signal is true;
	signal G9416: std_logic; attribute dont_touch of G9416: signal is true;
	signal G9417: std_logic; attribute dont_touch of G9417: signal is true;
	signal G9418: std_logic; attribute dont_touch of G9418: signal is true;
	signal G9419: std_logic; attribute dont_touch of G9419: signal is true;
	signal G9420: std_logic; attribute dont_touch of G9420: signal is true;
	signal G9421: std_logic; attribute dont_touch of G9421: signal is true;
	signal G9422: std_logic; attribute dont_touch of G9422: signal is true;
	signal G9423: std_logic; attribute dont_touch of G9423: signal is true;
	signal G9424: std_logic; attribute dont_touch of G9424: signal is true;
	signal G9425: std_logic; attribute dont_touch of G9425: signal is true;
	signal G9426: std_logic; attribute dont_touch of G9426: signal is true;
	signal G9427: std_logic; attribute dont_touch of G9427: signal is true;
	signal G9428: std_logic; attribute dont_touch of G9428: signal is true;
	signal G9429: std_logic; attribute dont_touch of G9429: signal is true;
	signal G9430: std_logic; attribute dont_touch of G9430: signal is true;
	signal G9431: std_logic; attribute dont_touch of G9431: signal is true;
	signal G9432: std_logic; attribute dont_touch of G9432: signal is true;
	signal G9447: std_logic; attribute dont_touch of G9447: signal is true;
	signal G9448: std_logic; attribute dont_touch of G9448: signal is true;
	signal G9449: std_logic; attribute dont_touch of G9449: signal is true;
	signal G9450: std_logic; attribute dont_touch of G9450: signal is true;
	signal G9452: std_logic; attribute dont_touch of G9452: signal is true;
	signal G9453: std_logic; attribute dont_touch of G9453: signal is true;
	signal G9454: std_logic; attribute dont_touch of G9454: signal is true;
	signal G9473: std_logic; attribute dont_touch of G9473: signal is true;
	signal G9474: std_logic; attribute dont_touch of G9474: signal is true;
	signal G9489: std_logic; attribute dont_touch of G9489: signal is true;
	signal G9490: std_logic; attribute dont_touch of G9490: signal is true;
	signal G9505: std_logic; attribute dont_touch of G9505: signal is true;
	signal G9506: std_logic; attribute dont_touch of G9506: signal is true;
	signal G9507: std_logic; attribute dont_touch of G9507: signal is true;
	signal G9508: std_logic; attribute dont_touch of G9508: signal is true;
	signal G9509: std_logic; attribute dont_touch of G9509: signal is true;
	signal G9510: std_logic; attribute dont_touch of G9510: signal is true;
	signal G9511: std_logic; attribute dont_touch of G9511: signal is true;
	signal G9512: std_logic; attribute dont_touch of G9512: signal is true;
	signal G9515: std_logic; attribute dont_touch of G9515: signal is true;
	signal G9516: std_logic; attribute dont_touch of G9516: signal is true;
	signal G9519: std_logic; attribute dont_touch of G9519: signal is true;
	signal G9522: std_logic; attribute dont_touch of G9522: signal is true;
	signal G9525: std_logic; attribute dont_touch of G9525: signal is true;
	signal G9526: std_logic; attribute dont_touch of G9526: signal is true;
	signal G9527: std_logic; attribute dont_touch of G9527: signal is true;
	signal G9528: std_logic; attribute dont_touch of G9528: signal is true;
	signal G9529: std_logic; attribute dont_touch of G9529: signal is true;
	signal G9530: std_logic; attribute dont_touch of G9530: signal is true;
	signal G9531: std_logic; attribute dont_touch of G9531: signal is true;
	signal G9532: std_logic; attribute dont_touch of G9532: signal is true;
	signal G9533: std_logic; attribute dont_touch of G9533: signal is true;
	signal G9534: std_logic; attribute dont_touch of G9534: signal is true;
	signal G9535: std_logic; attribute dont_touch of G9535: signal is true;
	signal G9536: std_logic; attribute dont_touch of G9536: signal is true;
	signal G9553: std_logic; attribute dont_touch of G9553: signal is true;
	signal G9554: std_logic; attribute dont_touch of G9554: signal is true;
	signal G9555: std_logic; attribute dont_touch of G9555: signal is true;
	signal G9556: std_logic; attribute dont_touch of G9556: signal is true;
	signal G9557: std_logic; attribute dont_touch of G9557: signal is true;
	signal G9560: std_logic; attribute dont_touch of G9560: signal is true;
	signal G9563: std_logic; attribute dont_touch of G9563: signal is true;
	signal G9566: std_logic; attribute dont_touch of G9566: signal is true;
	signal G9569: std_logic; attribute dont_touch of G9569: signal is true;
	signal G9572: std_logic; attribute dont_touch of G9572: signal is true;
	signal G9573: std_logic; attribute dont_touch of G9573: signal is true;
	signal G9576: std_logic; attribute dont_touch of G9576: signal is true;
	signal G9579: std_logic; attribute dont_touch of G9579: signal is true;
	signal G9582: std_logic; attribute dont_touch of G9582: signal is true;
	signal G9583: std_logic; attribute dont_touch of G9583: signal is true;
	signal G9584: std_logic; attribute dont_touch of G9584: signal is true;
	signal G9585: std_logic; attribute dont_touch of G9585: signal is true;
	signal G9586: std_logic; attribute dont_touch of G9586: signal is true;
	signal G9587: std_logic; attribute dont_touch of G9587: signal is true;
	signal G9588: std_logic; attribute dont_touch of G9588: signal is true;
	signal G9589: std_logic; attribute dont_touch of G9589: signal is true;
	signal G9590: std_logic; attribute dont_touch of G9590: signal is true;
	signal G9591: std_logic; attribute dont_touch of G9591: signal is true;
	signal G9592: std_logic; attribute dont_touch of G9592: signal is true;
	signal G9593: std_logic; attribute dont_touch of G9593: signal is true;
	signal G9594: std_logic; attribute dont_touch of G9594: signal is true;
	signal G9595: std_logic; attribute dont_touch of G9595: signal is true;
	signal G9596: std_logic; attribute dont_touch of G9596: signal is true;
	signal G9597: std_logic; attribute dont_touch of G9597: signal is true;
	signal G9598: std_logic; attribute dont_touch of G9598: signal is true;
	signal G9599: std_logic; attribute dont_touch of G9599: signal is true;
	signal G9600: std_logic; attribute dont_touch of G9600: signal is true;
	signal G9601: std_logic; attribute dont_touch of G9601: signal is true;
	signal G9602: std_logic; attribute dont_touch of G9602: signal is true;
	signal G9603: std_logic; attribute dont_touch of G9603: signal is true;
	signal G9604: std_logic; attribute dont_touch of G9604: signal is true;
	signal G9605: std_logic; attribute dont_touch of G9605: signal is true;
	signal G9606: std_logic; attribute dont_touch of G9606: signal is true;
	signal G9607: std_logic; attribute dont_touch of G9607: signal is true;
	signal G9608: std_logic; attribute dont_touch of G9608: signal is true;
	signal G9609: std_logic; attribute dont_touch of G9609: signal is true;
	signal G9610: std_logic; attribute dont_touch of G9610: signal is true;
	signal G9611: std_logic; attribute dont_touch of G9611: signal is true;
	signal G9612: std_logic; attribute dont_touch of G9612: signal is true;
	signal G9613: std_logic; attribute dont_touch of G9613: signal is true;
	signal G9614: std_logic; attribute dont_touch of G9614: signal is true;
	signal G9615: std_logic; attribute dont_touch of G9615: signal is true;
	signal G9616: std_logic; attribute dont_touch of G9616: signal is true;
	signal G9617: std_logic; attribute dont_touch of G9617: signal is true;
	signal G9618: std_logic; attribute dont_touch of G9618: signal is true;
	signal G9619: std_logic; attribute dont_touch of G9619: signal is true;
	signal G9620: std_logic; attribute dont_touch of G9620: signal is true;
	signal G9621: std_logic; attribute dont_touch of G9621: signal is true;
	signal G9622: std_logic; attribute dont_touch of G9622: signal is true;
	signal G9623: std_logic; attribute dont_touch of G9623: signal is true;
	signal G9624: std_logic; attribute dont_touch of G9624: signal is true;
	signal G9641: std_logic; attribute dont_touch of G9641: signal is true;
	signal G9642: std_logic; attribute dont_touch of G9642: signal is true;
	signal G9643: std_logic; attribute dont_touch of G9643: signal is true;
	signal G9644: std_logic; attribute dont_touch of G9644: signal is true;
	signal G9645: std_logic; attribute dont_touch of G9645: signal is true;
	signal G9646: std_logic; attribute dont_touch of G9646: signal is true;
	signal G9647: std_logic; attribute dont_touch of G9647: signal is true;
	signal G9648: std_logic; attribute dont_touch of G9648: signal is true;
	signal G9649: std_logic; attribute dont_touch of G9649: signal is true;
	signal G9650: std_logic; attribute dont_touch of G9650: signal is true;
	signal G9651: std_logic; attribute dont_touch of G9651: signal is true;
	signal G9652: std_logic; attribute dont_touch of G9652: signal is true;
	signal G9653: std_logic; attribute dont_touch of G9653: signal is true;
	signal G9654: std_logic; attribute dont_touch of G9654: signal is true;
	signal G9655: std_logic; attribute dont_touch of G9655: signal is true;
	signal G9656: std_logic; attribute dont_touch of G9656: signal is true;
	signal G9657: std_logic; attribute dont_touch of G9657: signal is true;
	signal G9658: std_logic; attribute dont_touch of G9658: signal is true;
	signal G9659: std_logic; attribute dont_touch of G9659: signal is true;
	signal G9660: std_logic; attribute dont_touch of G9660: signal is true;
	signal G9661: std_logic; attribute dont_touch of G9661: signal is true;
	signal G9662: std_logic; attribute dont_touch of G9662: signal is true;
	signal G9663: std_logic; attribute dont_touch of G9663: signal is true;
	signal G9664: std_logic; attribute dont_touch of G9664: signal is true;
	signal G9665: std_logic; attribute dont_touch of G9665: signal is true;
	signal G9666: std_logic; attribute dont_touch of G9666: signal is true;
	signal G9667: std_logic; attribute dont_touch of G9667: signal is true;
	signal G9668: std_logic; attribute dont_touch of G9668: signal is true;
	signal G9669: std_logic; attribute dont_touch of G9669: signal is true;
	signal G9670: std_logic; attribute dont_touch of G9670: signal is true;
	signal G9671: std_logic; attribute dont_touch of G9671: signal is true;
	signal G9672: std_logic; attribute dont_touch of G9672: signal is true;
	signal G9673: std_logic; attribute dont_touch of G9673: signal is true;
	signal G9676: std_logic; attribute dont_touch of G9676: signal is true;
	signal G9679: std_logic; attribute dont_touch of G9679: signal is true;
	signal G9680: std_logic; attribute dont_touch of G9680: signal is true;
	signal G9683: std_logic; attribute dont_touch of G9683: signal is true;
	signal G9686: std_logic; attribute dont_touch of G9686: signal is true;
	signal G9689: std_logic; attribute dont_touch of G9689: signal is true;
	signal G9690: std_logic; attribute dont_touch of G9690: signal is true;
	signal G9691: std_logic; attribute dont_touch of G9691: signal is true;
	signal G9692: std_logic; attribute dont_touch of G9692: signal is true;
	signal G9693: std_logic; attribute dont_touch of G9693: signal is true;
	signal G9694: std_logic; attribute dont_touch of G9694: signal is true;
	signal G9695: std_logic; attribute dont_touch of G9695: signal is true;
	signal G9696: std_logic; attribute dont_touch of G9696: signal is true;
	signal G9697: std_logic; attribute dont_touch of G9697: signal is true;
	signal G9698: std_logic; attribute dont_touch of G9698: signal is true;
	signal G9699: std_logic; attribute dont_touch of G9699: signal is true;
	signal G9700: std_logic; attribute dont_touch of G9700: signal is true;
	signal G9701: std_logic; attribute dont_touch of G9701: signal is true;
	signal G9702: std_logic; attribute dont_touch of G9702: signal is true;
	signal G9703: std_logic; attribute dont_touch of G9703: signal is true;
	signal G9704: std_logic; attribute dont_touch of G9704: signal is true;
	signal G9705: std_logic; attribute dont_touch of G9705: signal is true;
	signal G9706: std_logic; attribute dont_touch of G9706: signal is true;
	signal G9707: std_logic; attribute dont_touch of G9707: signal is true;
	signal G9708: std_logic; attribute dont_touch of G9708: signal is true;
	signal G9709: std_logic; attribute dont_touch of G9709: signal is true;
	signal G9710: std_logic; attribute dont_touch of G9710: signal is true;
	signal G9711: std_logic; attribute dont_touch of G9711: signal is true;
	signal G9712: std_logic; attribute dont_touch of G9712: signal is true;
	signal G9713: std_logic; attribute dont_touch of G9713: signal is true;
	signal G9714: std_logic; attribute dont_touch of G9714: signal is true;
	signal G9715: std_logic; attribute dont_touch of G9715: signal is true;
	signal G9716: std_logic; attribute dont_touch of G9716: signal is true;
	signal G9717: std_logic; attribute dont_touch of G9717: signal is true;
	signal G9718: std_logic; attribute dont_touch of G9718: signal is true;
	signal G9719: std_logic; attribute dont_touch of G9719: signal is true;
	signal G9720: std_logic; attribute dont_touch of G9720: signal is true;
	signal G9721: std_logic; attribute dont_touch of G9721: signal is true;
	signal G9722: std_logic; attribute dont_touch of G9722: signal is true;
	signal G9723: std_logic; attribute dont_touch of G9723: signal is true;
	signal G9724: std_logic; attribute dont_touch of G9724: signal is true;
	signal G9725: std_logic; attribute dont_touch of G9725: signal is true;
	signal G9726: std_logic; attribute dont_touch of G9726: signal is true;
	signal G9727: std_logic; attribute dont_touch of G9727: signal is true;
	signal G9728: std_logic; attribute dont_touch of G9728: signal is true;
	signal G9729: std_logic; attribute dont_touch of G9729: signal is true;
	signal G9730: std_logic; attribute dont_touch of G9730: signal is true;
	signal G9731: std_logic; attribute dont_touch of G9731: signal is true;
	signal G9732: std_logic; attribute dont_touch of G9732: signal is true;
	signal G9733: std_logic; attribute dont_touch of G9733: signal is true;
	signal G9734: std_logic; attribute dont_touch of G9734: signal is true;
	signal G9735: std_logic; attribute dont_touch of G9735: signal is true;
	signal G9736: std_logic; attribute dont_touch of G9736: signal is true;
	signal G9737: std_logic; attribute dont_touch of G9737: signal is true;
	signal G9738: std_logic; attribute dont_touch of G9738: signal is true;
	signal G9739: std_logic; attribute dont_touch of G9739: signal is true;
	signal G9740: std_logic; attribute dont_touch of G9740: signal is true;
	signal G9741: std_logic; attribute dont_touch of G9741: signal is true;
	signal G9742: std_logic; attribute dont_touch of G9742: signal is true;
	signal G9745: std_logic; attribute dont_touch of G9745: signal is true;
	signal G9746: std_logic; attribute dont_touch of G9746: signal is true;
	signal G9747: std_logic; attribute dont_touch of G9747: signal is true;
	signal G9750: std_logic; attribute dont_touch of G9750: signal is true;
	signal G9751: std_logic; attribute dont_touch of G9751: signal is true;
	signal G9754: std_logic; attribute dont_touch of G9754: signal is true;
	signal G9757: std_logic; attribute dont_touch of G9757: signal is true;
	signal G9758: std_logic; attribute dont_touch of G9758: signal is true;
	signal G9759: std_logic; attribute dont_touch of G9759: signal is true;
	signal G9760: std_logic; attribute dont_touch of G9760: signal is true;
	signal G9761: std_logic; attribute dont_touch of G9761: signal is true;
	signal G9762: std_logic; attribute dont_touch of G9762: signal is true;
	signal G9763: std_logic; attribute dont_touch of G9763: signal is true;
	signal G9764: std_logic; attribute dont_touch of G9764: signal is true;
	signal G9765: std_logic; attribute dont_touch of G9765: signal is true;
	signal G9766: std_logic; attribute dont_touch of G9766: signal is true;
	signal G9767: std_logic; attribute dont_touch of G9767: signal is true;
	signal G9768: std_logic; attribute dont_touch of G9768: signal is true;
	signal G9769: std_logic; attribute dont_touch of G9769: signal is true;
	signal G9770: std_logic; attribute dont_touch of G9770: signal is true;
	signal G9771: std_logic; attribute dont_touch of G9771: signal is true;
	signal G9772: std_logic; attribute dont_touch of G9772: signal is true;
	signal G9773: std_logic; attribute dont_touch of G9773: signal is true;
	signal G9774: std_logic; attribute dont_touch of G9774: signal is true;
	signal G9775: std_logic; attribute dont_touch of G9775: signal is true;
	signal G9776: std_logic; attribute dont_touch of G9776: signal is true;
	signal G9777: std_logic; attribute dont_touch of G9777: signal is true;
	signal G9778: std_logic; attribute dont_touch of G9778: signal is true;
	signal G9779: std_logic; attribute dont_touch of G9779: signal is true;
	signal G9780: std_logic; attribute dont_touch of G9780: signal is true;
	signal G9781: std_logic; attribute dont_touch of G9781: signal is true;
	signal G9782: std_logic; attribute dont_touch of G9782: signal is true;
	signal G9785: std_logic; attribute dont_touch of G9785: signal is true;
	signal G9802: std_logic; attribute dont_touch of G9802: signal is true;
	signal G9803: std_logic; attribute dont_touch of G9803: signal is true;
	signal G9804: std_logic; attribute dont_touch of G9804: signal is true;
	signal G9807: std_logic; attribute dont_touch of G9807: signal is true;
	signal G9808: std_logic; attribute dont_touch of G9808: signal is true;
	signal G9809: std_logic; attribute dont_touch of G9809: signal is true;
	signal G9812: std_logic; attribute dont_touch of G9812: signal is true;
	signal G9813: std_logic; attribute dont_touch of G9813: signal is true;
	signal G9814: std_logic; attribute dont_touch of G9814: signal is true;
	signal G9815: std_logic; attribute dont_touch of G9815: signal is true;
	signal G9816: std_logic; attribute dont_touch of G9816: signal is true;
	signal G9817: std_logic; attribute dont_touch of G9817: signal is true;
	signal G9818: std_logic; attribute dont_touch of G9818: signal is true;
	signal G9819: std_logic; attribute dont_touch of G9819: signal is true;
	signal G9820: std_logic; attribute dont_touch of G9820: signal is true;
	signal G9821: std_logic; attribute dont_touch of G9821: signal is true;
	signal G9822: std_logic; attribute dont_touch of G9822: signal is true;
	signal G9823: std_logic; attribute dont_touch of G9823: signal is true;
	signal G9824: std_logic; attribute dont_touch of G9824: signal is true;
	signal G9825: std_logic; attribute dont_touch of G9825: signal is true;
	signal G9826: std_logic; attribute dont_touch of G9826: signal is true;
	signal G9827: std_logic; attribute dont_touch of G9827: signal is true;
	signal G9828: std_logic; attribute dont_touch of G9828: signal is true;
	signal G9829: std_logic; attribute dont_touch of G9829: signal is true;
	signal G9830: std_logic; attribute dont_touch of G9830: signal is true;
	signal G9831: std_logic; attribute dont_touch of G9831: signal is true;
	signal G9832: std_logic; attribute dont_touch of G9832: signal is true;
	signal G9833: std_logic; attribute dont_touch of G9833: signal is true;
	signal G9834: std_logic; attribute dont_touch of G9834: signal is true;
	signal G9835: std_logic; attribute dont_touch of G9835: signal is true;
	signal G9836: std_logic; attribute dont_touch of G9836: signal is true;
	signal G9837: std_logic; attribute dont_touch of G9837: signal is true;
	signal G9838: std_logic; attribute dont_touch of G9838: signal is true;
	signal G9839: std_logic; attribute dont_touch of G9839: signal is true;
	signal G9840: std_logic; attribute dont_touch of G9840: signal is true;
	signal G9841: std_logic; attribute dont_touch of G9841: signal is true;
	signal G9842: std_logic; attribute dont_touch of G9842: signal is true;
	signal G9843: std_logic; attribute dont_touch of G9843: signal is true;
	signal G9844: std_logic; attribute dont_touch of G9844: signal is true;
	signal G9845: std_logic; attribute dont_touch of G9845: signal is true;
	signal G9846: std_logic; attribute dont_touch of G9846: signal is true;
	signal G9847: std_logic; attribute dont_touch of G9847: signal is true;
	signal G9848: std_logic; attribute dont_touch of G9848: signal is true;
	signal G9849: std_logic; attribute dont_touch of G9849: signal is true;
	signal G9850: std_logic; attribute dont_touch of G9850: signal is true;
	signal G9851: std_logic; attribute dont_touch of G9851: signal is true;
	signal G9852: std_logic; attribute dont_touch of G9852: signal is true;
	signal G9853: std_logic; attribute dont_touch of G9853: signal is true;
	signal G9854: std_logic; attribute dont_touch of G9854: signal is true;
	signal G9855: std_logic; attribute dont_touch of G9855: signal is true;
	signal G9856: std_logic; attribute dont_touch of G9856: signal is true;
	signal G9857: std_logic; attribute dont_touch of G9857: signal is true;
	signal G9858: std_logic; attribute dont_touch of G9858: signal is true;
	signal G9859: std_logic; attribute dont_touch of G9859: signal is true;
	signal G9860: std_logic; attribute dont_touch of G9860: signal is true;
	signal G9861: std_logic; attribute dont_touch of G9861: signal is true;
	signal G9862: std_logic; attribute dont_touch of G9862: signal is true;
	signal G9863: std_logic; attribute dont_touch of G9863: signal is true;
	signal G9864: std_logic; attribute dont_touch of G9864: signal is true;
	signal G9865: std_logic; attribute dont_touch of G9865: signal is true;
	signal G9866: std_logic; attribute dont_touch of G9866: signal is true;
	signal G9867: std_logic; attribute dont_touch of G9867: signal is true;
	signal G9868: std_logic; attribute dont_touch of G9868: signal is true;
	signal G9869: std_logic; attribute dont_touch of G9869: signal is true;
	signal G9870: std_logic; attribute dont_touch of G9870: signal is true;
	signal G9871: std_logic; attribute dont_touch of G9871: signal is true;
	signal G9872: std_logic; attribute dont_touch of G9872: signal is true;
	signal G9873: std_logic; attribute dont_touch of G9873: signal is true;
	signal G9874: std_logic; attribute dont_touch of G9874: signal is true;
	signal G9875: std_logic; attribute dont_touch of G9875: signal is true;
	signal G9876: std_logic; attribute dont_touch of G9876: signal is true;
	signal G9877: std_logic; attribute dont_touch of G9877: signal is true;
	signal G9878: std_logic; attribute dont_touch of G9878: signal is true;
	signal G9879: std_logic; attribute dont_touch of G9879: signal is true;
	signal G9880: std_logic; attribute dont_touch of G9880: signal is true;
	signal G9881: std_logic; attribute dont_touch of G9881: signal is true;
	signal G9882: std_logic; attribute dont_touch of G9882: signal is true;
	signal G9883: std_logic; attribute dont_touch of G9883: signal is true;
	signal G9884: std_logic; attribute dont_touch of G9884: signal is true;
	signal G9885: std_logic; attribute dont_touch of G9885: signal is true;
	signal G9886: std_logic; attribute dont_touch of G9886: signal is true;
	signal G9887: std_logic; attribute dont_touch of G9887: signal is true;
	signal G9888: std_logic; attribute dont_touch of G9888: signal is true;
	signal G9889: std_logic; attribute dont_touch of G9889: signal is true;
	signal G9890: std_logic; attribute dont_touch of G9890: signal is true;
	signal G9891: std_logic; attribute dont_touch of G9891: signal is true;
	signal G9892: std_logic; attribute dont_touch of G9892: signal is true;
	signal G9893: std_logic; attribute dont_touch of G9893: signal is true;
	signal G9894: std_logic; attribute dont_touch of G9894: signal is true;
	signal G9895: std_logic; attribute dont_touch of G9895: signal is true;
	signal G9896: std_logic; attribute dont_touch of G9896: signal is true;
	signal G9897: std_logic; attribute dont_touch of G9897: signal is true;
	signal G9898: std_logic; attribute dont_touch of G9898: signal is true;
	signal G9899: std_logic; attribute dont_touch of G9899: signal is true;
	signal G9900: std_logic; attribute dont_touch of G9900: signal is true;
	signal G9901: std_logic; attribute dont_touch of G9901: signal is true;
	signal G9902: std_logic; attribute dont_touch of G9902: signal is true;
	signal G9903: std_logic; attribute dont_touch of G9903: signal is true;
	signal G9904: std_logic; attribute dont_touch of G9904: signal is true;
	signal G9905: std_logic; attribute dont_touch of G9905: signal is true;
	signal G9906: std_logic; attribute dont_touch of G9906: signal is true;
	signal G9907: std_logic; attribute dont_touch of G9907: signal is true;
	signal G9908: std_logic; attribute dont_touch of G9908: signal is true;
	signal G9909: std_logic; attribute dont_touch of G9909: signal is true;
	signal G9910: std_logic; attribute dont_touch of G9910: signal is true;
	signal G9911: std_logic; attribute dont_touch of G9911: signal is true;
	signal G9912: std_logic; attribute dont_touch of G9912: signal is true;
	signal G9913: std_logic; attribute dont_touch of G9913: signal is true;
	signal G9914: std_logic; attribute dont_touch of G9914: signal is true;
	signal G9915: std_logic; attribute dont_touch of G9915: signal is true;
	signal G9916: std_logic; attribute dont_touch of G9916: signal is true;
	signal G9917: std_logic; attribute dont_touch of G9917: signal is true;
	signal G9918: std_logic; attribute dont_touch of G9918: signal is true;
	signal G9919: std_logic; attribute dont_touch of G9919: signal is true;
	signal G9920: std_logic; attribute dont_touch of G9920: signal is true;
	signal G9921: std_logic; attribute dont_touch of G9921: signal is true;
	signal G9922: std_logic; attribute dont_touch of G9922: signal is true;
	signal G9923: std_logic; attribute dont_touch of G9923: signal is true;
	signal G9924: std_logic; attribute dont_touch of G9924: signal is true;
	signal G9925: std_logic; attribute dont_touch of G9925: signal is true;
	signal G9926: std_logic; attribute dont_touch of G9926: signal is true;
	signal G9927: std_logic; attribute dont_touch of G9927: signal is true;
	signal G9928: std_logic; attribute dont_touch of G9928: signal is true;
	signal G9929: std_logic; attribute dont_touch of G9929: signal is true;
	signal G9930: std_logic; attribute dont_touch of G9930: signal is true;
	signal G9931: std_logic; attribute dont_touch of G9931: signal is true;
	signal G9932: std_logic; attribute dont_touch of G9932: signal is true;
	signal G9933: std_logic; attribute dont_touch of G9933: signal is true;
	signal G9934: std_logic; attribute dont_touch of G9934: signal is true;
	signal G9935: std_logic; attribute dont_touch of G9935: signal is true;
	signal G9936: std_logic; attribute dont_touch of G9936: signal is true;
	signal G9937: std_logic; attribute dont_touch of G9937: signal is true;
	signal G9938: std_logic; attribute dont_touch of G9938: signal is true;
	signal G9939: std_logic; attribute dont_touch of G9939: signal is true;
	signal G9940: std_logic; attribute dont_touch of G9940: signal is true;
	signal G9941: std_logic; attribute dont_touch of G9941: signal is true;
	signal G9942: std_logic; attribute dont_touch of G9942: signal is true;
	signal G9943: std_logic; attribute dont_touch of G9943: signal is true;
	signal G9944: std_logic; attribute dont_touch of G9944: signal is true;
	signal G9945: std_logic; attribute dont_touch of G9945: signal is true;
	signal G9946: std_logic; attribute dont_touch of G9946: signal is true;
	signal G9947: std_logic; attribute dont_touch of G9947: signal is true;
	signal G9948: std_logic; attribute dont_touch of G9948: signal is true;
	signal G9949: std_logic; attribute dont_touch of G9949: signal is true;
	signal G9950: std_logic; attribute dont_touch of G9950: signal is true;
	signal G9951: std_logic; attribute dont_touch of G9951: signal is true;
	signal G9952: std_logic; attribute dont_touch of G9952: signal is true;
	signal G9953: std_logic; attribute dont_touch of G9953: signal is true;
	signal G9954: std_logic; attribute dont_touch of G9954: signal is true;
	signal G9955: std_logic; attribute dont_touch of G9955: signal is true;
	signal G9956: std_logic; attribute dont_touch of G9956: signal is true;
	signal G9957: std_logic; attribute dont_touch of G9957: signal is true;
	signal G9958: std_logic; attribute dont_touch of G9958: signal is true;
	signal G9959: std_logic; attribute dont_touch of G9959: signal is true;
	signal G9960: std_logic; attribute dont_touch of G9960: signal is true;
	signal G9962: std_logic; attribute dont_touch of G9962: signal is true;
	signal G9963: std_logic; attribute dont_touch of G9963: signal is true;
	signal G9964: std_logic; attribute dont_touch of G9964: signal is true;
	signal G9965: std_logic; attribute dont_touch of G9965: signal is true;
	signal G9966: std_logic; attribute dont_touch of G9966: signal is true;
	signal G9967: std_logic; attribute dont_touch of G9967: signal is true;
	signal G9968: std_logic; attribute dont_touch of G9968: signal is true;
	signal G9974: std_logic; attribute dont_touch of G9974: signal is true;
	signal G9980: std_logic; attribute dont_touch of G9980: signal is true;
	signal G9984: std_logic; attribute dont_touch of G9984: signal is true;
	signal G9987: std_logic; attribute dont_touch of G9987: signal is true;
	signal G9990: std_logic; attribute dont_touch of G9990: signal is true;
	signal G9993: std_logic; attribute dont_touch of G9993: signal is true;
	signal G9994: std_logic; attribute dont_touch of G9994: signal is true;
	signal G9995: std_logic; attribute dont_touch of G9995: signal is true;
	signal G10001: std_logic; attribute dont_touch of G10001: signal is true;
	signal G10007: std_logic; attribute dont_touch of G10007: signal is true;
	signal G10013: std_logic; attribute dont_touch of G10013: signal is true;
	signal G10019: std_logic; attribute dont_touch of G10019: signal is true;
	signal G10025: std_logic; attribute dont_touch of G10025: signal is true;
	signal G10031: std_logic; attribute dont_touch of G10031: signal is true;
	signal G10032: std_logic; attribute dont_touch of G10032: signal is true;
	signal G10033: std_logic; attribute dont_touch of G10033: signal is true;
	signal G10034: std_logic; attribute dont_touch of G10034: signal is true;
	signal G10035: std_logic; attribute dont_touch of G10035: signal is true;
	signal G10039: std_logic; attribute dont_touch of G10039: signal is true;
	signal G10040: std_logic; attribute dont_touch of G10040: signal is true;
	signal G10041: std_logic; attribute dont_touch of G10041: signal is true;
	signal G10042: std_logic; attribute dont_touch of G10042: signal is true;
	signal G10043: std_logic; attribute dont_touch of G10043: signal is true;
	signal G10044: std_logic; attribute dont_touch of G10044: signal is true;
	signal G10047: std_logic; attribute dont_touch of G10047: signal is true;
	signal G10050: std_logic; attribute dont_touch of G10050: signal is true;
	signal G10051: std_logic; attribute dont_touch of G10051: signal is true;
	signal G10056: std_logic; attribute dont_touch of G10056: signal is true;
	signal G10057: std_logic; attribute dont_touch of G10057: signal is true;
	signal G10058: std_logic; attribute dont_touch of G10058: signal is true;
	signal G10062: std_logic; attribute dont_touch of G10062: signal is true;
	signal G10063: std_logic; attribute dont_touch of G10063: signal is true;
	signal G10064: std_logic; attribute dont_touch of G10064: signal is true;
	signal G10065: std_logic; attribute dont_touch of G10065: signal is true;
	signal G10069: std_logic; attribute dont_touch of G10069: signal is true;
	signal G10074: std_logic; attribute dont_touch of G10074: signal is true;
	signal G10075: std_logic; attribute dont_touch of G10075: signal is true;
	signal G10079: std_logic; attribute dont_touch of G10079: signal is true;
	signal G10080: std_logic; attribute dont_touch of G10080: signal is true;
	signal G10083: std_logic; attribute dont_touch of G10083: signal is true;
	signal G10087: std_logic; attribute dont_touch of G10087: signal is true;
	signal G10088: std_logic; attribute dont_touch of G10088: signal is true;
	signal G10091: std_logic; attribute dont_touch of G10091: signal is true;
	signal G10092: std_logic; attribute dont_touch of G10092: signal is true;
	signal G10093: std_logic; attribute dont_touch of G10093: signal is true;
	signal G10094: std_logic; attribute dont_touch of G10094: signal is true;
	signal G10098: std_logic; attribute dont_touch of G10098: signal is true;
	signal G10101: std_logic; attribute dont_touch of G10101: signal is true;
	signal G10104: std_logic; attribute dont_touch of G10104: signal is true;
	signal G10107: std_logic; attribute dont_touch of G10107: signal is true;
	signal G10110: std_logic; attribute dont_touch of G10110: signal is true;
	signal G10111: std_logic; attribute dont_touch of G10111: signal is true;
	signal G10114: std_logic; attribute dont_touch of G10114: signal is true;
	signal G10115: std_logic; attribute dont_touch of G10115: signal is true;
	signal G10116: std_logic; attribute dont_touch of G10116: signal is true;
	signal G10117: std_logic; attribute dont_touch of G10117: signal is true;
	signal G10118: std_logic; attribute dont_touch of G10118: signal is true;
	signal G10119: std_logic; attribute dont_touch of G10119: signal is true;
	signal G10120: std_logic; attribute dont_touch of G10120: signal is true;
	signal G10121: std_logic; attribute dont_touch of G10121: signal is true;
	signal G10122: std_logic; attribute dont_touch of G10122: signal is true;
	signal G10125: std_logic; attribute dont_touch of G10125: signal is true;
	signal G10126: std_logic; attribute dont_touch of G10126: signal is true;
	signal G10127: std_logic; attribute dont_touch of G10127: signal is true;
	signal G10128: std_logic; attribute dont_touch of G10128: signal is true;
	signal G10129: std_logic; attribute dont_touch of G10129: signal is true;
	signal G10130: std_logic; attribute dont_touch of G10130: signal is true;
	signal G10131: std_logic; attribute dont_touch of G10131: signal is true;
	signal G10132: std_logic; attribute dont_touch of G10132: signal is true;
	signal G10133: std_logic; attribute dont_touch of G10133: signal is true;
	signal G10134: std_logic; attribute dont_touch of G10134: signal is true;
	signal G10135: std_logic; attribute dont_touch of G10135: signal is true;
	signal G10136: std_logic; attribute dont_touch of G10136: signal is true;
	signal G10137: std_logic; attribute dont_touch of G10137: signal is true;
	signal G10138: std_logic; attribute dont_touch of G10138: signal is true;
	signal G10139: std_logic; attribute dont_touch of G10139: signal is true;
	signal G10140: std_logic; attribute dont_touch of G10140: signal is true;
	signal G10141: std_logic; attribute dont_touch of G10141: signal is true;
	signal G10142: std_logic; attribute dont_touch of G10142: signal is true;
	signal G10143: std_logic; attribute dont_touch of G10143: signal is true;
	signal G10144: std_logic; attribute dont_touch of G10144: signal is true;
	signal G10145: std_logic; attribute dont_touch of G10145: signal is true;
	signal G10148: std_logic; attribute dont_touch of G10148: signal is true;
	signal G10149: std_logic; attribute dont_touch of G10149: signal is true;
	signal G10150: std_logic; attribute dont_touch of G10150: signal is true;
	signal G10153: std_logic; attribute dont_touch of G10153: signal is true;
	signal G10154: std_logic; attribute dont_touch of G10154: signal is true;
	signal G10155: std_logic; attribute dont_touch of G10155: signal is true;
	signal G10156: std_logic; attribute dont_touch of G10156: signal is true;
	signal G10157: std_logic; attribute dont_touch of G10157: signal is true;
	signal G10158: std_logic; attribute dont_touch of G10158: signal is true;
	signal G10159: std_logic; attribute dont_touch of G10159: signal is true;
	signal G10160: std_logic; attribute dont_touch of G10160: signal is true;
	signal G10161: std_logic; attribute dont_touch of G10161: signal is true;
	signal G10162: std_logic; attribute dont_touch of G10162: signal is true;
	signal G10163: std_logic; attribute dont_touch of G10163: signal is true;
	signal G10164: std_logic; attribute dont_touch of G10164: signal is true;
	signal G10165: std_logic; attribute dont_touch of G10165: signal is true;
	signal G10166: std_logic; attribute dont_touch of G10166: signal is true;
	signal G10167: std_logic; attribute dont_touch of G10167: signal is true;
	signal G10168: std_logic; attribute dont_touch of G10168: signal is true;
	signal G10169: std_logic; attribute dont_touch of G10169: signal is true;
	signal G10170: std_logic; attribute dont_touch of G10170: signal is true;
	signal G10171: std_logic; attribute dont_touch of G10171: signal is true;
	signal G10172: std_logic; attribute dont_touch of G10172: signal is true;
	signal G10173: std_logic; attribute dont_touch of G10173: signal is true;
	signal G10174: std_logic; attribute dont_touch of G10174: signal is true;
	signal G10175: std_logic; attribute dont_touch of G10175: signal is true;
	signal G10176: std_logic; attribute dont_touch of G10176: signal is true;
	signal G10177: std_logic; attribute dont_touch of G10177: signal is true;
	signal G10178: std_logic; attribute dont_touch of G10178: signal is true;
	signal G10179: std_logic; attribute dont_touch of G10179: signal is true;
	signal G10182: std_logic; attribute dont_touch of G10182: signal is true;
	signal G10183: std_logic; attribute dont_touch of G10183: signal is true;
	signal G10184: std_logic; attribute dont_touch of G10184: signal is true;
	signal G10185: std_logic; attribute dont_touch of G10185: signal is true;
	signal G10186: std_logic; attribute dont_touch of G10186: signal is true;
	signal G10187: std_logic; attribute dont_touch of G10187: signal is true;
	signal G10188: std_logic; attribute dont_touch of G10188: signal is true;
	signal G10189: std_logic; attribute dont_touch of G10189: signal is true;
	signal G10190: std_logic; attribute dont_touch of G10190: signal is true;
	signal G10191: std_logic; attribute dont_touch of G10191: signal is true;
	signal G10192: std_logic; attribute dont_touch of G10192: signal is true;
	signal G10193: std_logic; attribute dont_touch of G10193: signal is true;
	signal G10194: std_logic; attribute dont_touch of G10194: signal is true;
	signal G10195: std_logic; attribute dont_touch of G10195: signal is true;
	signal G10196: std_logic; attribute dont_touch of G10196: signal is true;
	signal G10197: std_logic; attribute dont_touch of G10197: signal is true;
	signal G10198: std_logic; attribute dont_touch of G10198: signal is true;
	signal G10199: std_logic; attribute dont_touch of G10199: signal is true;
	signal G10200: std_logic; attribute dont_touch of G10200: signal is true;
	signal G10201: std_logic; attribute dont_touch of G10201: signal is true;
	signal G10202: std_logic; attribute dont_touch of G10202: signal is true;
	signal G10203: std_logic; attribute dont_touch of G10203: signal is true;
	signal G10204: std_logic; attribute dont_touch of G10204: signal is true;
	signal G10205: std_logic; attribute dont_touch of G10205: signal is true;
	signal G10206: std_logic; attribute dont_touch of G10206: signal is true;
	signal G10207: std_logic; attribute dont_touch of G10207: signal is true;
	signal G10208: std_logic; attribute dont_touch of G10208: signal is true;
	signal G10211: std_logic; attribute dont_touch of G10211: signal is true;
	signal G10214: std_logic; attribute dont_touch of G10214: signal is true;
	signal G10217: std_logic; attribute dont_touch of G10217: signal is true;
	signal G10220: std_logic; attribute dont_touch of G10220: signal is true;
	signal G10223: std_logic; attribute dont_touch of G10223: signal is true;
	signal G10226: std_logic; attribute dont_touch of G10226: signal is true;
	signal G10227: std_logic; attribute dont_touch of G10227: signal is true;
	signal G10228: std_logic; attribute dont_touch of G10228: signal is true;
	signal G10229: std_logic; attribute dont_touch of G10229: signal is true;
	signal G10230: std_logic; attribute dont_touch of G10230: signal is true;
	signal G10231: std_logic; attribute dont_touch of G10231: signal is true;
	signal G10232: std_logic; attribute dont_touch of G10232: signal is true;
	signal G10233: std_logic; attribute dont_touch of G10233: signal is true;
	signal G10234: std_logic; attribute dont_touch of G10234: signal is true;
	signal G10235: std_logic; attribute dont_touch of G10235: signal is true;
	signal G10236: std_logic; attribute dont_touch of G10236: signal is true;
	signal G10237: std_logic; attribute dont_touch of G10237: signal is true;
	signal G10238: std_logic; attribute dont_touch of G10238: signal is true;
	signal G10239: std_logic; attribute dont_touch of G10239: signal is true;
	signal G10240: std_logic; attribute dont_touch of G10240: signal is true;
	signal G10241: std_logic; attribute dont_touch of G10241: signal is true;
	signal G10242: std_logic; attribute dont_touch of G10242: signal is true;
	signal G10243: std_logic; attribute dont_touch of G10243: signal is true;
	signal G10244: std_logic; attribute dont_touch of G10244: signal is true;
	signal G10247: std_logic; attribute dont_touch of G10247: signal is true;
	signal G10248: std_logic; attribute dont_touch of G10248: signal is true;
	signal G10249: std_logic; attribute dont_touch of G10249: signal is true;
	signal G10250: std_logic; attribute dont_touch of G10250: signal is true;
	signal G10251: std_logic; attribute dont_touch of G10251: signal is true;
	signal G10252: std_logic; attribute dont_touch of G10252: signal is true;
	signal G10253: std_logic; attribute dont_touch of G10253: signal is true;
	signal G10254: std_logic; attribute dont_touch of G10254: signal is true;
	signal G10255: std_logic; attribute dont_touch of G10255: signal is true;
	signal G10256: std_logic; attribute dont_touch of G10256: signal is true;
	signal G10257: std_logic; attribute dont_touch of G10257: signal is true;
	signal G10258: std_logic; attribute dont_touch of G10258: signal is true;
	signal G10259: std_logic; attribute dont_touch of G10259: signal is true;
	signal G10260: std_logic; attribute dont_touch of G10260: signal is true;
	signal G10261: std_logic; attribute dont_touch of G10261: signal is true;
	signal G10262: std_logic; attribute dont_touch of G10262: signal is true;
	signal G10263: std_logic; attribute dont_touch of G10263: signal is true;
	signal G10264: std_logic; attribute dont_touch of G10264: signal is true;
	signal G10265: std_logic; attribute dont_touch of G10265: signal is true;
	signal G10266: std_logic; attribute dont_touch of G10266: signal is true;
	signal G10267: std_logic; attribute dont_touch of G10267: signal is true;
	signal G10268: std_logic; attribute dont_touch of G10268: signal is true;
	signal G10269: std_logic; attribute dont_touch of G10269: signal is true;
	signal G10270: std_logic; attribute dont_touch of G10270: signal is true;
	signal G10271: std_logic; attribute dont_touch of G10271: signal is true;
	signal G10272: std_logic; attribute dont_touch of G10272: signal is true;
	signal G10275: std_logic; attribute dont_touch of G10275: signal is true;
	signal G10276: std_logic; attribute dont_touch of G10276: signal is true;
	signal G10277: std_logic; attribute dont_touch of G10277: signal is true;
	signal G10278: std_logic; attribute dont_touch of G10278: signal is true;
	signal G10279: std_logic; attribute dont_touch of G10279: signal is true;
	signal G10280: std_logic; attribute dont_touch of G10280: signal is true;
	signal G10281: std_logic; attribute dont_touch of G10281: signal is true;
	signal G10282: std_logic; attribute dont_touch of G10282: signal is true;
	signal G10283: std_logic; attribute dont_touch of G10283: signal is true;
	signal G10284: std_logic; attribute dont_touch of G10284: signal is true;
	signal G10285: std_logic; attribute dont_touch of G10285: signal is true;
	signal G10286: std_logic; attribute dont_touch of G10286: signal is true;
	signal G10287: std_logic; attribute dont_touch of G10287: signal is true;
	signal G10288: std_logic; attribute dont_touch of G10288: signal is true;
	signal G10289: std_logic; attribute dont_touch of G10289: signal is true;
	signal G10290: std_logic; attribute dont_touch of G10290: signal is true;
	signal G10291: std_logic; attribute dont_touch of G10291: signal is true;
	signal G10292: std_logic; attribute dont_touch of G10292: signal is true;
	signal G10293: std_logic; attribute dont_touch of G10293: signal is true;
	signal G10294: std_logic; attribute dont_touch of G10294: signal is true;
	signal G10295: std_logic; attribute dont_touch of G10295: signal is true;
	signal G10296: std_logic; attribute dont_touch of G10296: signal is true;
	signal G10297: std_logic; attribute dont_touch of G10297: signal is true;
	signal G10298: std_logic; attribute dont_touch of G10298: signal is true;
	signal G10299: std_logic; attribute dont_touch of G10299: signal is true;
	signal G10300: std_logic; attribute dont_touch of G10300: signal is true;
	signal G10301: std_logic; attribute dont_touch of G10301: signal is true;
	signal G10302: std_logic; attribute dont_touch of G10302: signal is true;
	signal G10303: std_logic; attribute dont_touch of G10303: signal is true;
	signal G10304: std_logic; attribute dont_touch of G10304: signal is true;
	signal G10305: std_logic; attribute dont_touch of G10305: signal is true;
	signal G10306: std_logic; attribute dont_touch of G10306: signal is true;
	signal G10307: std_logic; attribute dont_touch of G10307: signal is true;
	signal G10308: std_logic; attribute dont_touch of G10308: signal is true;
	signal G10309: std_logic; attribute dont_touch of G10309: signal is true;
	signal G10310: std_logic; attribute dont_touch of G10310: signal is true;
	signal G10311: std_logic; attribute dont_touch of G10311: signal is true;
	signal G10312: std_logic; attribute dont_touch of G10312: signal is true;
	signal G10313: std_logic; attribute dont_touch of G10313: signal is true;
	signal G10314: std_logic; attribute dont_touch of G10314: signal is true;
	signal G10315: std_logic; attribute dont_touch of G10315: signal is true;
	signal G10316: std_logic; attribute dont_touch of G10316: signal is true;
	signal G10317: std_logic; attribute dont_touch of G10317: signal is true;
	signal G10318: std_logic; attribute dont_touch of G10318: signal is true;
	signal G10319: std_logic; attribute dont_touch of G10319: signal is true;
	signal G10320: std_logic; attribute dont_touch of G10320: signal is true;
	signal G10321: std_logic; attribute dont_touch of G10321: signal is true;
	signal G10322: std_logic; attribute dont_touch of G10322: signal is true;
	signal G10323: std_logic; attribute dont_touch of G10323: signal is true;
	signal G10324: std_logic; attribute dont_touch of G10324: signal is true;
	signal G10325: std_logic; attribute dont_touch of G10325: signal is true;
	signal G10326: std_logic; attribute dont_touch of G10326: signal is true;
	signal G10327: std_logic; attribute dont_touch of G10327: signal is true;
	signal G10328: std_logic; attribute dont_touch of G10328: signal is true;
	signal G10329: std_logic; attribute dont_touch of G10329: signal is true;
	signal G10330: std_logic; attribute dont_touch of G10330: signal is true;
	signal G10331: std_logic; attribute dont_touch of G10331: signal is true;
	signal G10332: std_logic; attribute dont_touch of G10332: signal is true;
	signal G10333: std_logic; attribute dont_touch of G10333: signal is true;
	signal G10334: std_logic; attribute dont_touch of G10334: signal is true;
	signal G10335: std_logic; attribute dont_touch of G10335: signal is true;
	signal G10336: std_logic; attribute dont_touch of G10336: signal is true;
	signal G10339: std_logic; attribute dont_touch of G10339: signal is true;
	signal G10342: std_logic; attribute dont_touch of G10342: signal is true;
	signal G10343: std_logic; attribute dont_touch of G10343: signal is true;
	signal G10344: std_logic; attribute dont_touch of G10344: signal is true;
	signal G10345: std_logic; attribute dont_touch of G10345: signal is true;
	signal G10346: std_logic; attribute dont_touch of G10346: signal is true;
	signal G10347: std_logic; attribute dont_touch of G10347: signal is true;
	signal G10348: std_logic; attribute dont_touch of G10348: signal is true;
	signal G10349: std_logic; attribute dont_touch of G10349: signal is true;
	signal G10350: std_logic; attribute dont_touch of G10350: signal is true;
	signal G10351: std_logic; attribute dont_touch of G10351: signal is true;
	signal G10352: std_logic; attribute dont_touch of G10352: signal is true;
	signal G10353: std_logic; attribute dont_touch of G10353: signal is true;
	signal G10354: std_logic; attribute dont_touch of G10354: signal is true;
	signal G10355: std_logic; attribute dont_touch of G10355: signal is true;
	signal G10356: std_logic; attribute dont_touch of G10356: signal is true;
	signal G10357: std_logic; attribute dont_touch of G10357: signal is true;
	signal G10358: std_logic; attribute dont_touch of G10358: signal is true;
	signal G10359: std_logic; attribute dont_touch of G10359: signal is true;
	signal G10360: std_logic; attribute dont_touch of G10360: signal is true;
	signal G10361: std_logic; attribute dont_touch of G10361: signal is true;
	signal G10362: std_logic; attribute dont_touch of G10362: signal is true;
	signal G10363: std_logic; attribute dont_touch of G10363: signal is true;
	signal G10364: std_logic; attribute dont_touch of G10364: signal is true;
	signal G10365: std_logic; attribute dont_touch of G10365: signal is true;
	signal G10366: std_logic; attribute dont_touch of G10366: signal is true;
	signal G10367: std_logic; attribute dont_touch of G10367: signal is true;
	signal G10368: std_logic; attribute dont_touch of G10368: signal is true;
	signal G10369: std_logic; attribute dont_touch of G10369: signal is true;
	signal G10370: std_logic; attribute dont_touch of G10370: signal is true;
	signal G10371: std_logic; attribute dont_touch of G10371: signal is true;
	signal G10372: std_logic; attribute dont_touch of G10372: signal is true;
	signal G10373: std_logic; attribute dont_touch of G10373: signal is true;
	signal G10374: std_logic; attribute dont_touch of G10374: signal is true;
	signal G10375: std_logic; attribute dont_touch of G10375: signal is true;
	signal G10376: std_logic; attribute dont_touch of G10376: signal is true;
	signal G10378: std_logic; attribute dont_touch of G10378: signal is true;
	signal G10380: std_logic; attribute dont_touch of G10380: signal is true;
	signal G10381: std_logic; attribute dont_touch of G10381: signal is true;
	signal G10382: std_logic; attribute dont_touch of G10382: signal is true;
	signal G10383: std_logic; attribute dont_touch of G10383: signal is true;
	signal G10384: std_logic; attribute dont_touch of G10384: signal is true;
	signal G10385: std_logic; attribute dont_touch of G10385: signal is true;
	signal G10386: std_logic; attribute dont_touch of G10386: signal is true;
	signal G10387: std_logic; attribute dont_touch of G10387: signal is true;
	signal G10388: std_logic; attribute dont_touch of G10388: signal is true;
	signal G10389: std_logic; attribute dont_touch of G10389: signal is true;
	signal G10390: std_logic; attribute dont_touch of G10390: signal is true;
	signal G10391: std_logic; attribute dont_touch of G10391: signal is true;
	signal G10392: std_logic; attribute dont_touch of G10392: signal is true;
	signal G10393: std_logic; attribute dont_touch of G10393: signal is true;
	signal G10394: std_logic; attribute dont_touch of G10394: signal is true;
	signal G10395: std_logic; attribute dont_touch of G10395: signal is true;
	signal G10396: std_logic; attribute dont_touch of G10396: signal is true;
	signal G10400: std_logic; attribute dont_touch of G10400: signal is true;
	signal G10401: std_logic; attribute dont_touch of G10401: signal is true;
	signal G10402: std_logic; attribute dont_touch of G10402: signal is true;
	signal G10405: std_logic; attribute dont_touch of G10405: signal is true;
	signal G10408: std_logic; attribute dont_touch of G10408: signal is true;
	signal G10411: std_logic; attribute dont_touch of G10411: signal is true;
	signal G10414: std_logic; attribute dont_touch of G10414: signal is true;
	signal G10417: std_logic; attribute dont_touch of G10417: signal is true;
	signal G10420: std_logic; attribute dont_touch of G10420: signal is true;
	signal G10421: std_logic; attribute dont_touch of G10421: signal is true;
	signal G10422: std_logic; attribute dont_touch of G10422: signal is true;
	signal G10423: std_logic; attribute dont_touch of G10423: signal is true;
	signal G10424: std_logic; attribute dont_touch of G10424: signal is true;
	signal G10425: std_logic; attribute dont_touch of G10425: signal is true;
	signal G10426: std_logic; attribute dont_touch of G10426: signal is true;
	signal G10427: std_logic; attribute dont_touch of G10427: signal is true;
	signal G10428: std_logic; attribute dont_touch of G10428: signal is true;
	signal G10429: std_logic; attribute dont_touch of G10429: signal is true;
	signal G10430: std_logic; attribute dont_touch of G10430: signal is true;
	signal G10431: std_logic; attribute dont_touch of G10431: signal is true;
	signal G10432: std_logic; attribute dont_touch of G10432: signal is true;
	signal G10433: std_logic; attribute dont_touch of G10433: signal is true;
	signal G10434: std_logic; attribute dont_touch of G10434: signal is true;
	signal G10435: std_logic; attribute dont_touch of G10435: signal is true;
	signal G10436: std_logic; attribute dont_touch of G10436: signal is true;
	signal G10437: std_logic; attribute dont_touch of G10437: signal is true;
	signal G10438: std_logic; attribute dont_touch of G10438: signal is true;
	signal G10439: std_logic; attribute dont_touch of G10439: signal is true;
	signal G10440: std_logic; attribute dont_touch of G10440: signal is true;
	signal G10441: std_logic; attribute dont_touch of G10441: signal is true;
	signal G10442: std_logic; attribute dont_touch of G10442: signal is true;
	signal G10443: std_logic; attribute dont_touch of G10443: signal is true;
	signal G10444: std_logic; attribute dont_touch of G10444: signal is true;
	signal G10445: std_logic; attribute dont_touch of G10445: signal is true;
	signal G10446: std_logic; attribute dont_touch of G10446: signal is true;
	signal G10447: std_logic; attribute dont_touch of G10447: signal is true;
	signal G10448: std_logic; attribute dont_touch of G10448: signal is true;
	signal G10449: std_logic; attribute dont_touch of G10449: signal is true;
	signal G10450: std_logic; attribute dont_touch of G10450: signal is true;
	signal G10451: std_logic; attribute dont_touch of G10451: signal is true;
	signal G10452: std_logic; attribute dont_touch of G10452: signal is true;
	signal G10453: std_logic; attribute dont_touch of G10453: signal is true;
	signal G10454: std_logic; attribute dont_touch of G10454: signal is true;
	signal G10456: std_logic; attribute dont_touch of G10456: signal is true;
	signal G10458: std_logic; attribute dont_touch of G10458: signal is true;
	signal G10460: std_logic; attribute dont_touch of G10460: signal is true;
	signal G10462: std_logic; attribute dont_touch of G10462: signal is true;
	signal G10464: std_logic; attribute dont_touch of G10464: signal is true;
	signal G10466: std_logic; attribute dont_touch of G10466: signal is true;
	signal G10467: std_logic; attribute dont_touch of G10467: signal is true;
	signal G10468: std_logic; attribute dont_touch of G10468: signal is true;
	signal G10469: std_logic; attribute dont_touch of G10469: signal is true;
	signal G10470: std_logic; attribute dont_touch of G10470: signal is true;
	signal G10471: std_logic; attribute dont_touch of G10471: signal is true;
	signal G10472: std_logic; attribute dont_touch of G10472: signal is true;
	signal G10473: std_logic; attribute dont_touch of G10473: signal is true;
	signal G10474: std_logic; attribute dont_touch of G10474: signal is true;
	signal G10475: std_logic; attribute dont_touch of G10475: signal is true;
	signal G10476: std_logic; attribute dont_touch of G10476: signal is true;
	signal G10477: std_logic; attribute dont_touch of G10477: signal is true;
	signal G10478: std_logic; attribute dont_touch of G10478: signal is true;
	signal G10479: std_logic; attribute dont_touch of G10479: signal is true;
	signal G10480: std_logic; attribute dont_touch of G10480: signal is true;
	signal G10481: std_logic; attribute dont_touch of G10481: signal is true;
	signal G10482: std_logic; attribute dont_touch of G10482: signal is true;
	signal G10483: std_logic; attribute dont_touch of G10483: signal is true;
	signal G10484: std_logic; attribute dont_touch of G10484: signal is true;
	signal G10485: std_logic; attribute dont_touch of G10485: signal is true;
	signal G10486: std_logic; attribute dont_touch of G10486: signal is true;
	signal G10487: std_logic; attribute dont_touch of G10487: signal is true;
	signal G10488: std_logic; attribute dont_touch of G10488: signal is true;
	signal G10489: std_logic; attribute dont_touch of G10489: signal is true;
	signal G10490: std_logic; attribute dont_touch of G10490: signal is true;
	signal G10491: std_logic; attribute dont_touch of G10491: signal is true;
	signal G10492: std_logic; attribute dont_touch of G10492: signal is true;
	signal G10493: std_logic; attribute dont_touch of G10493: signal is true;
	signal G10494: std_logic; attribute dont_touch of G10494: signal is true;
	signal G10495: std_logic; attribute dont_touch of G10495: signal is true;
	signal G10496: std_logic; attribute dont_touch of G10496: signal is true;
	signal G10497: std_logic; attribute dont_touch of G10497: signal is true;
	signal G10498: std_logic; attribute dont_touch of G10498: signal is true;
	signal G10499: std_logic; attribute dont_touch of G10499: signal is true;
	signal G10500: std_logic; attribute dont_touch of G10500: signal is true;
	signal G10501: std_logic; attribute dont_touch of G10501: signal is true;
	signal G10502: std_logic; attribute dont_touch of G10502: signal is true;
	signal G10503: std_logic; attribute dont_touch of G10503: signal is true;
	signal G10504: std_logic; attribute dont_touch of G10504: signal is true;
	signal G10505: std_logic; attribute dont_touch of G10505: signal is true;
	signal G10506: std_logic; attribute dont_touch of G10506: signal is true;
	signal G10507: std_logic; attribute dont_touch of G10507: signal is true;
	signal G10508: std_logic; attribute dont_touch of G10508: signal is true;
	signal G10509: std_logic; attribute dont_touch of G10509: signal is true;
	signal G10510: std_logic; attribute dont_touch of G10510: signal is true;
	signal G10511: std_logic; attribute dont_touch of G10511: signal is true;
	signal G10512: std_logic; attribute dont_touch of G10512: signal is true;
	signal G10513: std_logic; attribute dont_touch of G10513: signal is true;
	signal G10514: std_logic; attribute dont_touch of G10514: signal is true;
	signal G10515: std_logic; attribute dont_touch of G10515: signal is true;
	signal G10518: std_logic; attribute dont_touch of G10518: signal is true;
	signal G10521: std_logic; attribute dont_touch of G10521: signal is true;
	signal G10522: std_logic; attribute dont_touch of G10522: signal is true;
	signal G10523: std_logic; attribute dont_touch of G10523: signal is true;
	signal G10524: std_logic; attribute dont_touch of G10524: signal is true;
	signal G10525: std_logic; attribute dont_touch of G10525: signal is true;
	signal G10526: std_logic; attribute dont_touch of G10526: signal is true;
	signal G10527: std_logic; attribute dont_touch of G10527: signal is true;
	signal G10528: std_logic; attribute dont_touch of G10528: signal is true;
	signal G10529: std_logic; attribute dont_touch of G10529: signal is true;
	signal G10530: std_logic; attribute dont_touch of G10530: signal is true;
	signal G10531: std_logic; attribute dont_touch of G10531: signal is true;
	signal G10532: std_logic; attribute dont_touch of G10532: signal is true;
	signal G10533: std_logic; attribute dont_touch of G10533: signal is true;
	signal G10534: std_logic; attribute dont_touch of G10534: signal is true;
	signal G10535: std_logic; attribute dont_touch of G10535: signal is true;
	signal G10536: std_logic; attribute dont_touch of G10536: signal is true;
	signal G10537: std_logic; attribute dont_touch of G10537: signal is true;
	signal G10538: std_logic; attribute dont_touch of G10538: signal is true;
	signal G10539: std_logic; attribute dont_touch of G10539: signal is true;
	signal G10540: std_logic; attribute dont_touch of G10540: signal is true;
	signal G10541: std_logic; attribute dont_touch of G10541: signal is true;
	signal G10542: std_logic; attribute dont_touch of G10542: signal is true;
	signal G10543: std_logic; attribute dont_touch of G10543: signal is true;
	signal G10544: std_logic; attribute dont_touch of G10544: signal is true;
	signal G10545: std_logic; attribute dont_touch of G10545: signal is true;
	signal G10546: std_logic; attribute dont_touch of G10546: signal is true;
	signal G10547: std_logic; attribute dont_touch of G10547: signal is true;
	signal G10548: std_logic; attribute dont_touch of G10548: signal is true;
	signal G10549: std_logic; attribute dont_touch of G10549: signal is true;
	signal G10550: std_logic; attribute dont_touch of G10550: signal is true;
	signal G10551: std_logic; attribute dont_touch of G10551: signal is true;
	signal G10552: std_logic; attribute dont_touch of G10552: signal is true;
	signal G10553: std_logic; attribute dont_touch of G10553: signal is true;
	signal G10554: std_logic; attribute dont_touch of G10554: signal is true;
	signal G10555: std_logic; attribute dont_touch of G10555: signal is true;
	signal G10556: std_logic; attribute dont_touch of G10556: signal is true;
	signal G10557: std_logic; attribute dont_touch of G10557: signal is true;
	signal G10558: std_logic; attribute dont_touch of G10558: signal is true;
	signal G10559: std_logic; attribute dont_touch of G10559: signal is true;
	signal G10560: std_logic; attribute dont_touch of G10560: signal is true;
	signal G10561: std_logic; attribute dont_touch of G10561: signal is true;
	signal G10562: std_logic; attribute dont_touch of G10562: signal is true;
	signal G10563: std_logic; attribute dont_touch of G10563: signal is true;
	signal G10564: std_logic; attribute dont_touch of G10564: signal is true;
	signal G10567: std_logic; attribute dont_touch of G10567: signal is true;
	signal G10570: std_logic; attribute dont_touch of G10570: signal is true;
	signal G10571: std_logic; attribute dont_touch of G10571: signal is true;
	signal G10574: std_logic; attribute dont_touch of G10574: signal is true;
	signal G10575: std_logic; attribute dont_touch of G10575: signal is true;
	signal G10576: std_logic; attribute dont_touch of G10576: signal is true;
	signal G10577: std_logic; attribute dont_touch of G10577: signal is true;
	signal G10578: std_logic; attribute dont_touch of G10578: signal is true;
	signal G10579: std_logic; attribute dont_touch of G10579: signal is true;
	signal G10580: std_logic; attribute dont_touch of G10580: signal is true;
	signal G10581: std_logic; attribute dont_touch of G10581: signal is true;
	signal G10582: std_logic; attribute dont_touch of G10582: signal is true;
	signal G10583: std_logic; attribute dont_touch of G10583: signal is true;
	signal G10584: std_logic; attribute dont_touch of G10584: signal is true;
	signal G10589: std_logic; attribute dont_touch of G10589: signal is true;
	signal G10590: std_logic; attribute dont_touch of G10590: signal is true;
	signal G10591: std_logic; attribute dont_touch of G10591: signal is true;
	signal G10592: std_logic; attribute dont_touch of G10592: signal is true;
	signal G10593: std_logic; attribute dont_touch of G10593: signal is true;
	signal G10594: std_logic; attribute dont_touch of G10594: signal is true;
	signal G10595: std_logic; attribute dont_touch of G10595: signal is true;
	signal G10596: std_logic; attribute dont_touch of G10596: signal is true;
	signal G10597: std_logic; attribute dont_touch of G10597: signal is true;
	signal G10598: std_logic; attribute dont_touch of G10598: signal is true;
	signal G10599: std_logic; attribute dont_touch of G10599: signal is true;
	signal G10600: std_logic; attribute dont_touch of G10600: signal is true;
	signal G10604: std_logic; attribute dont_touch of G10604: signal is true;
	signal G10608: std_logic; attribute dont_touch of G10608: signal is true;
	signal G10612: std_logic; attribute dont_touch of G10612: signal is true;
	signal G10616: std_logic; attribute dont_touch of G10616: signal is true;
	signal G10619: std_logic; attribute dont_touch of G10619: signal is true;
	signal G10620: std_logic; attribute dont_touch of G10620: signal is true;
	signal G10621: std_logic; attribute dont_touch of G10621: signal is true;
	signal G10622: std_logic; attribute dont_touch of G10622: signal is true;
	signal G10623: std_logic; attribute dont_touch of G10623: signal is true;
	signal G10624: std_logic; attribute dont_touch of G10624: signal is true;
	signal G10625: std_logic; attribute dont_touch of G10625: signal is true;
	signal G10626: std_logic; attribute dont_touch of G10626: signal is true;
	signal G10627: std_logic; attribute dont_touch of G10627: signal is true;
	signal G10629: std_logic; attribute dont_touch of G10629: signal is true;
	signal G10630: std_logic; attribute dont_touch of G10630: signal is true;
	signal G10633: std_logic; attribute dont_touch of G10633: signal is true;
	signal G10634: std_logic; attribute dont_touch of G10634: signal is true;
	signal G10635: std_logic; attribute dont_touch of G10635: signal is true;
	signal G10638: std_logic; attribute dont_touch of G10638: signal is true;
	signal G10639: std_logic; attribute dont_touch of G10639: signal is true;
	signal G10642: std_logic; attribute dont_touch of G10642: signal is true;
	signal G10643: std_logic; attribute dont_touch of G10643: signal is true;
	signal G10646: std_logic; attribute dont_touch of G10646: signal is true;
	signal G10649: std_logic; attribute dont_touch of G10649: signal is true;
	signal G10652: std_logic; attribute dont_touch of G10652: signal is true;
	signal G10655: std_logic; attribute dont_touch of G10655: signal is true;
	signal G10658: std_logic; attribute dont_touch of G10658: signal is true;
	signal G10661: std_logic; attribute dont_touch of G10661: signal is true;
	signal G10662: std_logic; attribute dont_touch of G10662: signal is true;
	signal G10663: std_logic; attribute dont_touch of G10663: signal is true;
	signal G10664: std_logic; attribute dont_touch of G10664: signal is true;
	signal G10665: std_logic; attribute dont_touch of G10665: signal is true;
	signal G10666: std_logic; attribute dont_touch of G10666: signal is true;
	signal G10667: std_logic; attribute dont_touch of G10667: signal is true;
	signal G10668: std_logic; attribute dont_touch of G10668: signal is true;
	signal G10669: std_logic; attribute dont_touch of G10669: signal is true;
	signal G10670: std_logic; attribute dont_touch of G10670: signal is true;
	signal G10671: std_logic; attribute dont_touch of G10671: signal is true;
	signal G10672: std_logic; attribute dont_touch of G10672: signal is true;
	signal G10673: std_logic; attribute dont_touch of G10673: signal is true;
	signal G10674: std_logic; attribute dont_touch of G10674: signal is true;
	signal G10675: std_logic; attribute dont_touch of G10675: signal is true;
	signal G10676: std_logic; attribute dont_touch of G10676: signal is true;
	signal G10679: std_logic; attribute dont_touch of G10679: signal is true;
	signal G10680: std_logic; attribute dont_touch of G10680: signal is true;
	signal G10681: std_logic; attribute dont_touch of G10681: signal is true;
	signal G10682: std_logic; attribute dont_touch of G10682: signal is true;
	signal G10683: std_logic; attribute dont_touch of G10683: signal is true;
	signal G10684: std_logic; attribute dont_touch of G10684: signal is true;
	signal G10685: std_logic; attribute dont_touch of G10685: signal is true;
	signal G10686: std_logic; attribute dont_touch of G10686: signal is true;
	signal G10687: std_logic; attribute dont_touch of G10687: signal is true;
	signal G10690: std_logic; attribute dont_touch of G10690: signal is true;
	signal G10691: std_logic; attribute dont_touch of G10691: signal is true;
	signal G10692: std_logic; attribute dont_touch of G10692: signal is true;
	signal G10695: std_logic; attribute dont_touch of G10695: signal is true;
	signal G10696: std_logic; attribute dont_touch of G10696: signal is true;
	signal G10697: std_logic; attribute dont_touch of G10697: signal is true;
	signal G10698: std_logic; attribute dont_touch of G10698: signal is true;
	signal G10699: std_logic; attribute dont_touch of G10699: signal is true;
	signal G10700: std_logic; attribute dont_touch of G10700: signal is true;
	signal G10701: std_logic; attribute dont_touch of G10701: signal is true;
	signal G10702: std_logic; attribute dont_touch of G10702: signal is true;
	signal G10705: std_logic; attribute dont_touch of G10705: signal is true;
	signal G10706: std_logic; attribute dont_touch of G10706: signal is true;
	signal G10707: std_logic; attribute dont_touch of G10707: signal is true;
	signal G10708: std_logic; attribute dont_touch of G10708: signal is true;
	signal G10711: std_logic; attribute dont_touch of G10711: signal is true;
	signal G10712: std_logic; attribute dont_touch of G10712: signal is true;
	signal G10715: std_logic; attribute dont_touch of G10715: signal is true;
	signal G10716: std_logic; attribute dont_touch of G10716: signal is true;
	signal G10717: std_logic; attribute dont_touch of G10717: signal is true;
	signal G10718: std_logic; attribute dont_touch of G10718: signal is true;
	signal G10719: std_logic; attribute dont_touch of G10719: signal is true;
	signal G10720: std_logic; attribute dont_touch of G10720: signal is true;
	signal G10721: std_logic; attribute dont_touch of G10721: signal is true;
	signal G10722: std_logic; attribute dont_touch of G10722: signal is true;
	signal G10723: std_logic; attribute dont_touch of G10723: signal is true;
	signal G10724: std_logic; attribute dont_touch of G10724: signal is true;
	signal G10725: std_logic; attribute dont_touch of G10725: signal is true;
	signal G10726: std_logic; attribute dont_touch of G10726: signal is true;
	signal G10727: std_logic; attribute dont_touch of G10727: signal is true;
	signal G10728: std_logic; attribute dont_touch of G10728: signal is true;
	signal G10729: std_logic; attribute dont_touch of G10729: signal is true;
	signal G10730: std_logic; attribute dont_touch of G10730: signal is true;
	signal G10731: std_logic; attribute dont_touch of G10731: signal is true;
	signal G10732: std_logic; attribute dont_touch of G10732: signal is true;
	signal G10733: std_logic; attribute dont_touch of G10733: signal is true;
	signal G10734: std_logic; attribute dont_touch of G10734: signal is true;
	signal G10735: std_logic; attribute dont_touch of G10735: signal is true;
	signal G10736: std_logic; attribute dont_touch of G10736: signal is true;
	signal G10737: std_logic; attribute dont_touch of G10737: signal is true;
	signal G10738: std_logic; attribute dont_touch of G10738: signal is true;
	signal G10739: std_logic; attribute dont_touch of G10739: signal is true;
	signal G10740: std_logic; attribute dont_touch of G10740: signal is true;
	signal G10741: std_logic; attribute dont_touch of G10741: signal is true;
	signal G10742: std_logic; attribute dont_touch of G10742: signal is true;
	signal G10743: std_logic; attribute dont_touch of G10743: signal is true;
	signal G10744: std_logic; attribute dont_touch of G10744: signal is true;
	signal G10745: std_logic; attribute dont_touch of G10745: signal is true;
	signal G10746: std_logic; attribute dont_touch of G10746: signal is true;
	signal G10747: std_logic; attribute dont_touch of G10747: signal is true;
	signal G10750: std_logic; attribute dont_touch of G10750: signal is true;
	signal G10751: std_logic; attribute dont_touch of G10751: signal is true;
	signal G10752: std_logic; attribute dont_touch of G10752: signal is true;
	signal G10753: std_logic; attribute dont_touch of G10753: signal is true;
	signal G10754: std_logic; attribute dont_touch of G10754: signal is true;
	signal G10758: std_logic; attribute dont_touch of G10758: signal is true;
	signal G10759: std_logic; attribute dont_touch of G10759: signal is true;
	signal G10760: std_logic; attribute dont_touch of G10760: signal is true;
	signal G10761: std_logic; attribute dont_touch of G10761: signal is true;
	signal G10762: std_logic; attribute dont_touch of G10762: signal is true;
	signal G10763: std_logic; attribute dont_touch of G10763: signal is true;
	signal G10764: std_logic; attribute dont_touch of G10764: signal is true;
	signal G10765: std_logic; attribute dont_touch of G10765: signal is true;
	signal G10766: std_logic; attribute dont_touch of G10766: signal is true;
	signal G10767: std_logic; attribute dont_touch of G10767: signal is true;
	signal G10768: std_logic; attribute dont_touch of G10768: signal is true;
	signal G10769: std_logic; attribute dont_touch of G10769: signal is true;
	signal G10770: std_logic; attribute dont_touch of G10770: signal is true;
	signal G10771: std_logic; attribute dont_touch of G10771: signal is true;
	signal G10772: std_logic; attribute dont_touch of G10772: signal is true;
	signal G10773: std_logic; attribute dont_touch of G10773: signal is true;
	signal G10774: std_logic; attribute dont_touch of G10774: signal is true;
	signal G10775: std_logic; attribute dont_touch of G10775: signal is true;
	signal G10776: std_logic; attribute dont_touch of G10776: signal is true;
	signal G10777: std_logic; attribute dont_touch of G10777: signal is true;
	signal G10778: std_logic; attribute dont_touch of G10778: signal is true;
	signal G10779: std_logic; attribute dont_touch of G10779: signal is true;
	signal G10780: std_logic; attribute dont_touch of G10780: signal is true;
	signal G10781: std_logic; attribute dont_touch of G10781: signal is true;
	signal G10782: std_logic; attribute dont_touch of G10782: signal is true;
	signal G10783: std_logic; attribute dont_touch of G10783: signal is true;
	signal G10784: std_logic; attribute dont_touch of G10784: signal is true;
	signal G10785: std_logic; attribute dont_touch of G10785: signal is true;
	signal G10786: std_logic; attribute dont_touch of G10786: signal is true;
	signal G10787: std_logic; attribute dont_touch of G10787: signal is true;
	signal G10788: std_logic; attribute dont_touch of G10788: signal is true;
	signal G10791: std_logic; attribute dont_touch of G10791: signal is true;
	signal G10792: std_logic; attribute dont_touch of G10792: signal is true;
	signal G10793: std_logic; attribute dont_touch of G10793: signal is true;
	signal G10794: std_logic; attribute dont_touch of G10794: signal is true;
	signal G10795: std_logic; attribute dont_touch of G10795: signal is true;
	signal G10796: std_logic; attribute dont_touch of G10796: signal is true;
	signal G10797: std_logic; attribute dont_touch of G10797: signal is true;
	signal G10798: std_logic; attribute dont_touch of G10798: signal is true;
	signal G10799: std_logic; attribute dont_touch of G10799: signal is true;
	signal G10800: std_logic; attribute dont_touch of G10800: signal is true;
	signal G10802: std_logic; attribute dont_touch of G10802: signal is true;
	signal G10803: std_logic; attribute dont_touch of G10803: signal is true;
	signal G10804: std_logic; attribute dont_touch of G10804: signal is true;
	signal G10805: std_logic; attribute dont_touch of G10805: signal is true;
	signal G10806: std_logic; attribute dont_touch of G10806: signal is true;
	signal G10807: std_logic; attribute dont_touch of G10807: signal is true;
	signal G10808: std_logic; attribute dont_touch of G10808: signal is true;
	signal G10809: std_logic; attribute dont_touch of G10809: signal is true;
	signal G10818: std_logic; attribute dont_touch of G10818: signal is true;
	signal G10819: std_logic; attribute dont_touch of G10819: signal is true;
	signal G10820: std_logic; attribute dont_touch of G10820: signal is true;
	signal G10821: std_logic; attribute dont_touch of G10821: signal is true;
	signal G10822: std_logic; attribute dont_touch of G10822: signal is true;
	signal G10825: std_logic; attribute dont_touch of G10825: signal is true;
	signal G10826: std_logic; attribute dont_touch of G10826: signal is true;
	signal G10827: std_logic; attribute dont_touch of G10827: signal is true;
	signal G10848: std_logic; attribute dont_touch of G10848: signal is true;
	signal G10849: std_logic; attribute dont_touch of G10849: signal is true;
	signal G10850: std_logic; attribute dont_touch of G10850: signal is true;
	signal G10851: std_logic; attribute dont_touch of G10851: signal is true;
	signal G10852: std_logic; attribute dont_touch of G10852: signal is true;
	signal G10853: std_logic; attribute dont_touch of G10853: signal is true;
	signal G10854: std_logic; attribute dont_touch of G10854: signal is true;
	signal G10855: std_logic; attribute dont_touch of G10855: signal is true;
	signal G10856: std_logic; attribute dont_touch of G10856: signal is true;
	signal G10857: std_logic; attribute dont_touch of G10857: signal is true;
	signal G10858: std_logic; attribute dont_touch of G10858: signal is true;
	signal G10859: std_logic; attribute dont_touch of G10859: signal is true;
	signal G10860: std_logic; attribute dont_touch of G10860: signal is true;
	signal G10861: std_logic; attribute dont_touch of G10861: signal is true;
	signal G10862: std_logic; attribute dont_touch of G10862: signal is true;
	signal G10863: std_logic; attribute dont_touch of G10863: signal is true;
	signal G10864: std_logic; attribute dont_touch of G10864: signal is true;
	signal G10865: std_logic; attribute dont_touch of G10865: signal is true;
	signal G10866: std_logic; attribute dont_touch of G10866: signal is true;
	signal G10867: std_logic; attribute dont_touch of G10867: signal is true;
	signal G10868: std_logic; attribute dont_touch of G10868: signal is true;
	signal G10869: std_logic; attribute dont_touch of G10869: signal is true;
	signal G10870: std_logic; attribute dont_touch of G10870: signal is true;
	signal G10871: std_logic; attribute dont_touch of G10871: signal is true;
	signal G10872: std_logic; attribute dont_touch of G10872: signal is true;
	signal G10873: std_logic; attribute dont_touch of G10873: signal is true;
	signal G10874: std_logic; attribute dont_touch of G10874: signal is true;
	signal G10875: std_logic; attribute dont_touch of G10875: signal is true;
	signal G10876: std_logic; attribute dont_touch of G10876: signal is true;
	signal G10877: std_logic; attribute dont_touch of G10877: signal is true;
	signal G10878: std_logic; attribute dont_touch of G10878: signal is true;
	signal G10879: std_logic; attribute dont_touch of G10879: signal is true;
	signal G10880: std_logic; attribute dont_touch of G10880: signal is true;
	signal G10881: std_logic; attribute dont_touch of G10881: signal is true;
	signal G10882: std_logic; attribute dont_touch of G10882: signal is true;
	signal G10883: std_logic; attribute dont_touch of G10883: signal is true;
	signal G10884: std_logic; attribute dont_touch of G10884: signal is true;
	signal G10885: std_logic; attribute dont_touch of G10885: signal is true;
	signal G10886: std_logic; attribute dont_touch of G10886: signal is true;
	signal G10887: std_logic; attribute dont_touch of G10887: signal is true;
	signal G10888: std_logic; attribute dont_touch of G10888: signal is true;
	signal G10889: std_logic; attribute dont_touch of G10889: signal is true;
	signal G10890: std_logic; attribute dont_touch of G10890: signal is true;
	signal G10891: std_logic; attribute dont_touch of G10891: signal is true;
	signal G10892: std_logic; attribute dont_touch of G10892: signal is true;
	signal G10893: std_logic; attribute dont_touch of G10893: signal is true;
	signal G10894: std_logic; attribute dont_touch of G10894: signal is true;
	signal G10895: std_logic; attribute dont_touch of G10895: signal is true;
	signal G10896: std_logic; attribute dont_touch of G10896: signal is true;
	signal G10897: std_logic; attribute dont_touch of G10897: signal is true;
	signal G10898: std_logic; attribute dont_touch of G10898: signal is true;
	signal G10899: std_logic; attribute dont_touch of G10899: signal is true;
	signal G10900: std_logic; attribute dont_touch of G10900: signal is true;
	signal G10901: std_logic; attribute dont_touch of G10901: signal is true;
	signal G10902: std_logic; attribute dont_touch of G10902: signal is true;
	signal G10903: std_logic; attribute dont_touch of G10903: signal is true;
	signal G10904: std_logic; attribute dont_touch of G10904: signal is true;
	signal G10905: std_logic; attribute dont_touch of G10905: signal is true;
	signal G10906: std_logic; attribute dont_touch of G10906: signal is true;
	signal G10907: std_logic; attribute dont_touch of G10907: signal is true;
	signal G10908: std_logic; attribute dont_touch of G10908: signal is true;
	signal G10909: std_logic; attribute dont_touch of G10909: signal is true;
	signal G10910: std_logic; attribute dont_touch of G10910: signal is true;
	signal G10911: std_logic; attribute dont_touch of G10911: signal is true;
	signal G10912: std_logic; attribute dont_touch of G10912: signal is true;
	signal G10913: std_logic; attribute dont_touch of G10913: signal is true;
	signal G10923: std_logic; attribute dont_touch of G10923: signal is true;
	signal G10926: std_logic; attribute dont_touch of G10926: signal is true;
	signal G10927: std_logic; attribute dont_touch of G10927: signal is true;
	signal G10928: std_logic; attribute dont_touch of G10928: signal is true;
	signal G10929: std_logic; attribute dont_touch of G10929: signal is true;
	signal G10930: std_logic; attribute dont_touch of G10930: signal is true;
	signal G10931: std_logic; attribute dont_touch of G10931: signal is true;
	signal G10932: std_logic; attribute dont_touch of G10932: signal is true;
	signal G10933: std_logic; attribute dont_touch of G10933: signal is true;
	signal G10934: std_logic; attribute dont_touch of G10934: signal is true;
	signal G10935: std_logic; attribute dont_touch of G10935: signal is true;
	signal G10936: std_logic; attribute dont_touch of G10936: signal is true;
	signal G10937: std_logic; attribute dont_touch of G10937: signal is true;
	signal G10946: std_logic; attribute dont_touch of G10946: signal is true;
	signal G10947: std_logic; attribute dont_touch of G10947: signal is true;
	signal G10948: std_logic; attribute dont_touch of G10948: signal is true;
	signal G10949: std_logic; attribute dont_touch of G10949: signal is true;
	signal G10950: std_logic; attribute dont_touch of G10950: signal is true;
	signal G10969: std_logic; attribute dont_touch of G10969: signal is true;
	signal G10970: std_logic; attribute dont_touch of G10970: signal is true;
	signal G10971: std_logic; attribute dont_touch of G10971: signal is true;
	signal G10972: std_logic; attribute dont_touch of G10972: signal is true;
	signal G10973: std_logic; attribute dont_touch of G10973: signal is true;
	signal G10974: std_logic; attribute dont_touch of G10974: signal is true;
	signal G11005: std_logic; attribute dont_touch of G11005: signal is true;
	signal G11006: std_logic; attribute dont_touch of G11006: signal is true;
	signal G11007: std_logic; attribute dont_touch of G11007: signal is true;
	signal G11008: std_logic; attribute dont_touch of G11008: signal is true;
	signal G11009: std_logic; attribute dont_touch of G11009: signal is true;
	signal G11010: std_logic; attribute dont_touch of G11010: signal is true;
	signal G11011: std_logic; attribute dont_touch of G11011: signal is true;
	signal G11012: std_logic; attribute dont_touch of G11012: signal is true;
	signal G11013: std_logic; attribute dont_touch of G11013: signal is true;
	signal G11014: std_logic; attribute dont_touch of G11014: signal is true;
	signal G11015: std_logic; attribute dont_touch of G11015: signal is true;
	signal G11016: std_logic; attribute dont_touch of G11016: signal is true;
	signal G11017: std_logic; attribute dont_touch of G11017: signal is true;
	signal G11018: std_logic; attribute dont_touch of G11018: signal is true;
	signal G11019: std_logic; attribute dont_touch of G11019: signal is true;
	signal G11020: std_logic; attribute dont_touch of G11020: signal is true;
	signal G11021: std_logic; attribute dont_touch of G11021: signal is true;
	signal G11022: std_logic; attribute dont_touch of G11022: signal is true;
	signal G11023: std_logic; attribute dont_touch of G11023: signal is true;
	signal G11024: std_logic; attribute dont_touch of G11024: signal is true;
	signal G11025: std_logic; attribute dont_touch of G11025: signal is true;
	signal G11026: std_logic; attribute dont_touch of G11026: signal is true;
	signal G11027: std_logic; attribute dont_touch of G11027: signal is true;
	signal G11028: std_logic; attribute dont_touch of G11028: signal is true;
	signal G11029: std_logic; attribute dont_touch of G11029: signal is true;
	signal G11030: std_logic; attribute dont_touch of G11030: signal is true;
	signal G11031: std_logic; attribute dont_touch of G11031: signal is true;
	signal G11032: std_logic; attribute dont_touch of G11032: signal is true;
	signal G11033: std_logic; attribute dont_touch of G11033: signal is true;
	signal G11034: std_logic; attribute dont_touch of G11034: signal is true;
	signal G11035: std_logic; attribute dont_touch of G11035: signal is true;
	signal G11036: std_logic; attribute dont_touch of G11036: signal is true;
	signal G11037: std_logic; attribute dont_touch of G11037: signal is true;
	signal G11038: std_logic; attribute dont_touch of G11038: signal is true;
	signal G11039: std_logic; attribute dont_touch of G11039: signal is true;
	signal G11040: std_logic; attribute dont_touch of G11040: signal is true;
	signal G11041: std_logic; attribute dont_touch of G11041: signal is true;
	signal G11042: std_logic; attribute dont_touch of G11042: signal is true;
	signal G11043: std_logic; attribute dont_touch of G11043: signal is true;
	signal G11044: std_logic; attribute dont_touch of G11044: signal is true;
	signal G11045: std_logic; attribute dont_touch of G11045: signal is true;
	signal G11046: std_logic; attribute dont_touch of G11046: signal is true;
	signal G11047: std_logic; attribute dont_touch of G11047: signal is true;
	signal G11048: std_logic; attribute dont_touch of G11048: signal is true;
	signal G11049: std_logic; attribute dont_touch of G11049: signal is true;
	signal G11050: std_logic; attribute dont_touch of G11050: signal is true;
	signal G11051: std_logic; attribute dont_touch of G11051: signal is true;
	signal G11052: std_logic; attribute dont_touch of G11052: signal is true;
	signal G11053: std_logic; attribute dont_touch of G11053: signal is true;
	signal G11054: std_logic; attribute dont_touch of G11054: signal is true;
	signal G11055: std_logic; attribute dont_touch of G11055: signal is true;
	signal G11056: std_logic; attribute dont_touch of G11056: signal is true;
	signal G11057: std_logic; attribute dont_touch of G11057: signal is true;
	signal G11058: std_logic; attribute dont_touch of G11058: signal is true;
	signal G11059: std_logic; attribute dont_touch of G11059: signal is true;
	signal G11060: std_logic; attribute dont_touch of G11060: signal is true;
	signal G11061: std_logic; attribute dont_touch of G11061: signal is true;
	signal G11062: std_logic; attribute dont_touch of G11062: signal is true;
	signal G11063: std_logic; attribute dont_touch of G11063: signal is true;
	signal G11064: std_logic; attribute dont_touch of G11064: signal is true;
	signal G11065: std_logic; attribute dont_touch of G11065: signal is true;
	signal G11066: std_logic; attribute dont_touch of G11066: signal is true;
	signal G11067: std_logic; attribute dont_touch of G11067: signal is true;
	signal G11068: std_logic; attribute dont_touch of G11068: signal is true;
	signal G11069: std_logic; attribute dont_touch of G11069: signal is true;
	signal G11070: std_logic; attribute dont_touch of G11070: signal is true;
	signal G11071: std_logic; attribute dont_touch of G11071: signal is true;
	signal G11072: std_logic; attribute dont_touch of G11072: signal is true;
	signal G11073: std_logic; attribute dont_touch of G11073: signal is true;
	signal G11074: std_logic; attribute dont_touch of G11074: signal is true;
	signal G11075: std_logic; attribute dont_touch of G11075: signal is true;
	signal G11076: std_logic; attribute dont_touch of G11076: signal is true;
	signal G11077: std_logic; attribute dont_touch of G11077: signal is true;
	signal G11078: std_logic; attribute dont_touch of G11078: signal is true;
	signal G11079: std_logic; attribute dont_touch of G11079: signal is true;
	signal G11080: std_logic; attribute dont_touch of G11080: signal is true;
	signal G11081: std_logic; attribute dont_touch of G11081: signal is true;
	signal G11082: std_logic; attribute dont_touch of G11082: signal is true;
	signal G11083: std_logic; attribute dont_touch of G11083: signal is true;
	signal G11084: std_logic; attribute dont_touch of G11084: signal is true;
	signal G11085: std_logic; attribute dont_touch of G11085: signal is true;
	signal G11086: std_logic; attribute dont_touch of G11086: signal is true;
	signal G11087: std_logic; attribute dont_touch of G11087: signal is true;
	signal G11088: std_logic; attribute dont_touch of G11088: signal is true;
	signal G11091: std_logic; attribute dont_touch of G11091: signal is true;
	signal G11092: std_logic; attribute dont_touch of G11092: signal is true;
	signal G11093: std_logic; attribute dont_touch of G11093: signal is true;
	signal G11094: std_logic; attribute dont_touch of G11094: signal is true;
	signal G11095: std_logic; attribute dont_touch of G11095: signal is true;
	signal G11096: std_logic; attribute dont_touch of G11096: signal is true;
	signal G11097: std_logic; attribute dont_touch of G11097: signal is true;
	signal G11098: std_logic; attribute dont_touch of G11098: signal is true;
	signal G11099: std_logic; attribute dont_touch of G11099: signal is true;
	signal G11100: std_logic; attribute dont_touch of G11100: signal is true;
	signal G11101: std_logic; attribute dont_touch of G11101: signal is true;
	signal G11102: std_logic; attribute dont_touch of G11102: signal is true;
	signal G11103: std_logic; attribute dont_touch of G11103: signal is true;
	signal G11104: std_logic; attribute dont_touch of G11104: signal is true;
	signal G11105: std_logic; attribute dont_touch of G11105: signal is true;
	signal G11106: std_logic; attribute dont_touch of G11106: signal is true;
	signal G11107: std_logic; attribute dont_touch of G11107: signal is true;
	signal G11108: std_logic; attribute dont_touch of G11108: signal is true;
	signal G11109: std_logic; attribute dont_touch of G11109: signal is true;
	signal G11110: std_logic; attribute dont_touch of G11110: signal is true;
	signal G11111: std_logic; attribute dont_touch of G11111: signal is true;
	signal G11112: std_logic; attribute dont_touch of G11112: signal is true;
	signal G11143: std_logic; attribute dont_touch of G11143: signal is true;
	signal G11144: std_logic; attribute dont_touch of G11144: signal is true;
	signal G11145: std_logic; attribute dont_touch of G11145: signal is true;
	signal G11146: std_logic; attribute dont_touch of G11146: signal is true;
	signal G11147: std_logic; attribute dont_touch of G11147: signal is true;
	signal G11148: std_logic; attribute dont_touch of G11148: signal is true;
	signal G11149: std_logic; attribute dont_touch of G11149: signal is true;
	signal G11150: std_logic; attribute dont_touch of G11150: signal is true;
	signal G11151: std_logic; attribute dont_touch of G11151: signal is true;
	signal G11152: std_logic; attribute dont_touch of G11152: signal is true;
	signal G11153: std_logic; attribute dont_touch of G11153: signal is true;
	signal G11154: std_logic; attribute dont_touch of G11154: signal is true;
	signal G11155: std_logic; attribute dont_touch of G11155: signal is true;
	signal G11156: std_logic; attribute dont_touch of G11156: signal is true;
	signal G11157: std_logic; attribute dont_touch of G11157: signal is true;
	signal G11158: std_logic; attribute dont_touch of G11158: signal is true;
	signal G11159: std_logic; attribute dont_touch of G11159: signal is true;
	signal G11160: std_logic; attribute dont_touch of G11160: signal is true;
	signal G11161: std_logic; attribute dont_touch of G11161: signal is true;
	signal G11162: std_logic; attribute dont_touch of G11162: signal is true;
	signal G11164: std_logic; attribute dont_touch of G11164: signal is true;
	signal G11165: std_logic; attribute dont_touch of G11165: signal is true;
	signal G11166: std_logic; attribute dont_touch of G11166: signal is true;
	signal G11167: std_logic; attribute dont_touch of G11167: signal is true;
	signal G11168: std_logic; attribute dont_touch of G11168: signal is true;
	signal G11169: std_logic; attribute dont_touch of G11169: signal is true;
	signal G11170: std_logic; attribute dont_touch of G11170: signal is true;
	signal G11171: std_logic; attribute dont_touch of G11171: signal is true;
	signal G11172: std_logic; attribute dont_touch of G11172: signal is true;
	signal G11173: std_logic; attribute dont_touch of G11173: signal is true;
	signal G11174: std_logic; attribute dont_touch of G11174: signal is true;
	signal G11175: std_logic; attribute dont_touch of G11175: signal is true;
	signal G11176: std_logic; attribute dont_touch of G11176: signal is true;
	signal G11177: std_logic; attribute dont_touch of G11177: signal is true;
	signal G11178: std_logic; attribute dont_touch of G11178: signal is true;
	signal G11179: std_logic; attribute dont_touch of G11179: signal is true;
	signal G11180: std_logic; attribute dont_touch of G11180: signal is true;
	signal G11181: std_logic; attribute dont_touch of G11181: signal is true;
	signal G11182: std_logic; attribute dont_touch of G11182: signal is true;
	signal G11183: std_logic; attribute dont_touch of G11183: signal is true;
	signal G11184: std_logic; attribute dont_touch of G11184: signal is true;
	signal G11185: std_logic; attribute dont_touch of G11185: signal is true;
	signal G11186: std_logic; attribute dont_touch of G11186: signal is true;
	signal G11187: std_logic; attribute dont_touch of G11187: signal is true;
	signal G11188: std_logic; attribute dont_touch of G11188: signal is true;
	signal G11189: std_logic; attribute dont_touch of G11189: signal is true;
	signal G11190: std_logic; attribute dont_touch of G11190: signal is true;
	signal G11191: std_logic; attribute dont_touch of G11191: signal is true;
	signal G11192: std_logic; attribute dont_touch of G11192: signal is true;
	signal G11193: std_logic; attribute dont_touch of G11193: signal is true;
	signal G11194: std_logic; attribute dont_touch of G11194: signal is true;
	signal G11195: std_logic; attribute dont_touch of G11195: signal is true;
	signal G11196: std_logic; attribute dont_touch of G11196: signal is true;
	signal G11197: std_logic; attribute dont_touch of G11197: signal is true;
	signal G11198: std_logic; attribute dont_touch of G11198: signal is true;
	signal G11199: std_logic; attribute dont_touch of G11199: signal is true;
	signal G11200: std_logic; attribute dont_touch of G11200: signal is true;
	signal G11201: std_logic; attribute dont_touch of G11201: signal is true;
	signal G11202: std_logic; attribute dont_touch of G11202: signal is true;
	signal G11203: std_logic; attribute dont_touch of G11203: signal is true;
	signal G11204: std_logic; attribute dont_touch of G11204: signal is true;
	signal G11205: std_logic; attribute dont_touch of G11205: signal is true;
	signal G11207: std_logic; attribute dont_touch of G11207: signal is true;
	signal G11208: std_logic; attribute dont_touch of G11208: signal is true;
	signal G11209: std_logic; attribute dont_touch of G11209: signal is true;
	signal G11210: std_logic; attribute dont_touch of G11210: signal is true;
	signal G11211: std_logic; attribute dont_touch of G11211: signal is true;
	signal G11212: std_logic; attribute dont_touch of G11212: signal is true;
	signal G11213: std_logic; attribute dont_touch of G11213: signal is true;
	signal G11214: std_logic; attribute dont_touch of G11214: signal is true;
	signal G11215: std_logic; attribute dont_touch of G11215: signal is true;
	signal G11216: std_logic; attribute dont_touch of G11216: signal is true;
	signal G11217: std_logic; attribute dont_touch of G11217: signal is true;
	signal G11218: std_logic; attribute dont_touch of G11218: signal is true;
	signal G11219: std_logic; attribute dont_touch of G11219: signal is true;
	signal G11220: std_logic; attribute dont_touch of G11220: signal is true;
	signal G11221: std_logic; attribute dont_touch of G11221: signal is true;
	signal G11222: std_logic; attribute dont_touch of G11222: signal is true;
	signal G11223: std_logic; attribute dont_touch of G11223: signal is true;
	signal G11224: std_logic; attribute dont_touch of G11224: signal is true;
	signal G11225: std_logic; attribute dont_touch of G11225: signal is true;
	signal G11226: std_logic; attribute dont_touch of G11226: signal is true;
	signal G11227: std_logic; attribute dont_touch of G11227: signal is true;
	signal G11228: std_logic; attribute dont_touch of G11228: signal is true;
	signal G11229: std_logic; attribute dont_touch of G11229: signal is true;
	signal G11230: std_logic; attribute dont_touch of G11230: signal is true;
	signal G11231: std_logic; attribute dont_touch of G11231: signal is true;
	signal G11232: std_logic; attribute dont_touch of G11232: signal is true;
	signal G11233: std_logic; attribute dont_touch of G11233: signal is true;
	signal G11234: std_logic; attribute dont_touch of G11234: signal is true;
	signal G11235: std_logic; attribute dont_touch of G11235: signal is true;
	signal G11236: std_logic; attribute dont_touch of G11236: signal is true;
	signal G11237: std_logic; attribute dont_touch of G11237: signal is true;
	signal G11238: std_logic; attribute dont_touch of G11238: signal is true;
	signal G11239: std_logic; attribute dont_touch of G11239: signal is true;
	signal G11240: std_logic; attribute dont_touch of G11240: signal is true;
	signal G11241: std_logic; attribute dont_touch of G11241: signal is true;
	signal G11242: std_logic; attribute dont_touch of G11242: signal is true;
	signal G11243: std_logic; attribute dont_touch of G11243: signal is true;
	signal G11244: std_logic; attribute dont_touch of G11244: signal is true;
	signal G11245: std_logic; attribute dont_touch of G11245: signal is true;
	signal G11246: std_logic; attribute dont_touch of G11246: signal is true;
	signal G11247: std_logic; attribute dont_touch of G11247: signal is true;
	signal G11248: std_logic; attribute dont_touch of G11248: signal is true;
	signal G11249: std_logic; attribute dont_touch of G11249: signal is true;
	signal G11252: std_logic; attribute dont_touch of G11252: signal is true;
	signal G11253: std_logic; attribute dont_touch of G11253: signal is true;
	signal G11254: std_logic; attribute dont_touch of G11254: signal is true;
	signal G11255: std_logic; attribute dont_touch of G11255: signal is true;
	signal G11256: std_logic; attribute dont_touch of G11256: signal is true;
	signal G11257: std_logic; attribute dont_touch of G11257: signal is true;
	signal G11258: std_logic; attribute dont_touch of G11258: signal is true;
	signal G11259: std_logic; attribute dont_touch of G11259: signal is true;
	signal G11260: std_logic; attribute dont_touch of G11260: signal is true;
	signal G11261: std_logic; attribute dont_touch of G11261: signal is true;
	signal G11262: std_logic; attribute dont_touch of G11262: signal is true;
	signal G11263: std_logic; attribute dont_touch of G11263: signal is true;
	signal G11264: std_logic; attribute dont_touch of G11264: signal is true;
	signal G11265: std_logic; attribute dont_touch of G11265: signal is true;
	signal G11266: std_logic; attribute dont_touch of G11266: signal is true;
	signal G11267: std_logic; attribute dont_touch of G11267: signal is true;
	signal G11268: std_logic; attribute dont_touch of G11268: signal is true;
	signal G11269: std_logic; attribute dont_touch of G11269: signal is true;
	signal G11270: std_logic; attribute dont_touch of G11270: signal is true;
	signal G11271: std_logic; attribute dont_touch of G11271: signal is true;
	signal G11272: std_logic; attribute dont_touch of G11272: signal is true;
	signal G11273: std_logic; attribute dont_touch of G11273: signal is true;
	signal G11274: std_logic; attribute dont_touch of G11274: signal is true;
	signal G11275: std_logic; attribute dont_touch of G11275: signal is true;
	signal G11276: std_logic; attribute dont_touch of G11276: signal is true;
	signal G11277: std_logic; attribute dont_touch of G11277: signal is true;
	signal G11278: std_logic; attribute dont_touch of G11278: signal is true;
	signal G11279: std_logic; attribute dont_touch of G11279: signal is true;
	signal G11280: std_logic; attribute dont_touch of G11280: signal is true;
	signal G11281: std_logic; attribute dont_touch of G11281: signal is true;
	signal G11282: std_logic; attribute dont_touch of G11282: signal is true;
	signal G11283: std_logic; attribute dont_touch of G11283: signal is true;
	signal G11284: std_logic; attribute dont_touch of G11284: signal is true;
	signal G11285: std_logic; attribute dont_touch of G11285: signal is true;
	signal G11286: std_logic; attribute dont_touch of G11286: signal is true;
	signal G11287: std_logic; attribute dont_touch of G11287: signal is true;
	signal G11288: std_logic; attribute dont_touch of G11288: signal is true;
	signal G11289: std_logic; attribute dont_touch of G11289: signal is true;
	signal G11290: std_logic; attribute dont_touch of G11290: signal is true;
	signal G11291: std_logic; attribute dont_touch of G11291: signal is true;
	signal G11292: std_logic; attribute dont_touch of G11292: signal is true;
	signal G11293: std_logic; attribute dont_touch of G11293: signal is true;
	signal G11294: std_logic; attribute dont_touch of G11294: signal is true;
	signal G11295: std_logic; attribute dont_touch of G11295: signal is true;
	signal G11296: std_logic; attribute dont_touch of G11296: signal is true;
	signal G11297: std_logic; attribute dont_touch of G11297: signal is true;
	signal G11298: std_logic; attribute dont_touch of G11298: signal is true;
	signal G11299: std_logic; attribute dont_touch of G11299: signal is true;
	signal G11300: std_logic; attribute dont_touch of G11300: signal is true;
	signal G11301: std_logic; attribute dont_touch of G11301: signal is true;
	signal G11302: std_logic; attribute dont_touch of G11302: signal is true;
	signal G11303: std_logic; attribute dont_touch of G11303: signal is true;
	signal G11304: std_logic; attribute dont_touch of G11304: signal is true;
	signal G11305: std_logic; attribute dont_touch of G11305: signal is true;
	signal G11306: std_logic; attribute dont_touch of G11306: signal is true;
	signal G11307: std_logic; attribute dont_touch of G11307: signal is true;
	signal G11308: std_logic; attribute dont_touch of G11308: signal is true;
	signal G11309: std_logic; attribute dont_touch of G11309: signal is true;
	signal G11310: std_logic; attribute dont_touch of G11310: signal is true;
	signal G11311: std_logic; attribute dont_touch of G11311: signal is true;
	signal G11312: std_logic; attribute dont_touch of G11312: signal is true;
	signal G11313: std_logic; attribute dont_touch of G11313: signal is true;
	signal G11314: std_logic; attribute dont_touch of G11314: signal is true;
	signal G11315: std_logic; attribute dont_touch of G11315: signal is true;
	signal G11316: std_logic; attribute dont_touch of G11316: signal is true;
	signal G11317: std_logic; attribute dont_touch of G11317: signal is true;
	signal G11318: std_logic; attribute dont_touch of G11318: signal is true;
	signal G11319: std_logic; attribute dont_touch of G11319: signal is true;
	signal G11320: std_logic; attribute dont_touch of G11320: signal is true;
	signal G11321: std_logic; attribute dont_touch of G11321: signal is true;
	signal G11322: std_logic; attribute dont_touch of G11322: signal is true;
	signal G11323: std_logic; attribute dont_touch of G11323: signal is true;
	signal G11324: std_logic; attribute dont_touch of G11324: signal is true;
	signal G11325: std_logic; attribute dont_touch of G11325: signal is true;
	signal G11326: std_logic; attribute dont_touch of G11326: signal is true;
	signal G11327: std_logic; attribute dont_touch of G11327: signal is true;
	signal G11328: std_logic; attribute dont_touch of G11328: signal is true;
	signal G11329: std_logic; attribute dont_touch of G11329: signal is true;
	signal G11330: std_logic; attribute dont_touch of G11330: signal is true;
	signal G11331: std_logic; attribute dont_touch of G11331: signal is true;
	signal G11332: std_logic; attribute dont_touch of G11332: signal is true;
	signal G11333: std_logic; attribute dont_touch of G11333: signal is true;
	signal G11334: std_logic; attribute dont_touch of G11334: signal is true;
	signal G11335: std_logic; attribute dont_touch of G11335: signal is true;
	signal G11336: std_logic; attribute dont_touch of G11336: signal is true;
	signal G11337: std_logic; attribute dont_touch of G11337: signal is true;
	signal G11338: std_logic; attribute dont_touch of G11338: signal is true;
	signal G11339: std_logic; attribute dont_touch of G11339: signal is true;
	signal G11340: std_logic; attribute dont_touch of G11340: signal is true;
	signal G11341: std_logic; attribute dont_touch of G11341: signal is true;
	signal G11342: std_logic; attribute dont_touch of G11342: signal is true;
	signal G11343: std_logic; attribute dont_touch of G11343: signal is true;
	signal G11344: std_logic; attribute dont_touch of G11344: signal is true;
	signal G11345: std_logic; attribute dont_touch of G11345: signal is true;
	signal G11346: std_logic; attribute dont_touch of G11346: signal is true;
	signal G11347: std_logic; attribute dont_touch of G11347: signal is true;
	signal G11348: std_logic; attribute dont_touch of G11348: signal is true;
	signal G11349: std_logic; attribute dont_touch of G11349: signal is true;
	signal G11350: std_logic; attribute dont_touch of G11350: signal is true;
	signal G11351: std_logic; attribute dont_touch of G11351: signal is true;
	signal G11352: std_logic; attribute dont_touch of G11352: signal is true;
	signal G11353: std_logic; attribute dont_touch of G11353: signal is true;
	signal G11354: std_logic; attribute dont_touch of G11354: signal is true;
	signal G11357: std_logic; attribute dont_touch of G11357: signal is true;
	signal G11360: std_logic; attribute dont_touch of G11360: signal is true;
	signal G11363: std_logic; attribute dont_touch of G11363: signal is true;
	signal G11366: std_logic; attribute dont_touch of G11366: signal is true;
	signal G11369: std_logic; attribute dont_touch of G11369: signal is true;
	signal G11372: std_logic; attribute dont_touch of G11372: signal is true;
	signal G11373: std_logic; attribute dont_touch of G11373: signal is true;
	signal G11376: std_logic; attribute dont_touch of G11376: signal is true;
	signal G11377: std_logic; attribute dont_touch of G11377: signal is true;
	signal G11380: std_logic; attribute dont_touch of G11380: signal is true;
	signal G11381: std_logic; attribute dont_touch of G11381: signal is true;
	signal G11384: std_logic; attribute dont_touch of G11384: signal is true;
	signal G11387: std_logic; attribute dont_touch of G11387: signal is true;
	signal G11388: std_logic; attribute dont_touch of G11388: signal is true;
	signal G11389: std_logic; attribute dont_touch of G11389: signal is true;
	signal G11390: std_logic; attribute dont_touch of G11390: signal is true;
	signal G11391: std_logic; attribute dont_touch of G11391: signal is true;
	signal G11392: std_logic; attribute dont_touch of G11392: signal is true;
	signal G11393: std_logic; attribute dont_touch of G11393: signal is true;
	signal G11394: std_logic; attribute dont_touch of G11394: signal is true;
	signal G11395: std_logic; attribute dont_touch of G11395: signal is true;
	signal G11396: std_logic; attribute dont_touch of G11396: signal is true;
	signal G11397: std_logic; attribute dont_touch of G11397: signal is true;
	signal G11398: std_logic; attribute dont_touch of G11398: signal is true;
	signal G11399: std_logic; attribute dont_touch of G11399: signal is true;
	signal G11400: std_logic; attribute dont_touch of G11400: signal is true;
	signal G11401: std_logic; attribute dont_touch of G11401: signal is true;
	signal G11402: std_logic; attribute dont_touch of G11402: signal is true;
	signal G11403: std_logic; attribute dont_touch of G11403: signal is true;
	signal G11404: std_logic; attribute dont_touch of G11404: signal is true;
	signal G11405: std_logic; attribute dont_touch of G11405: signal is true;
	signal G11406: std_logic; attribute dont_touch of G11406: signal is true;
	signal G11407: std_logic; attribute dont_touch of G11407: signal is true;
	signal G11408: std_logic; attribute dont_touch of G11408: signal is true;
	signal G11409: std_logic; attribute dont_touch of G11409: signal is true;
	signal G11410: std_logic; attribute dont_touch of G11410: signal is true;
	signal G11411: std_logic; attribute dont_touch of G11411: signal is true;
	signal G11412: std_logic; attribute dont_touch of G11412: signal is true;
	signal G11413: std_logic; attribute dont_touch of G11413: signal is true;
	signal G11414: std_logic; attribute dont_touch of G11414: signal is true;
	signal G11415: std_logic; attribute dont_touch of G11415: signal is true;
	signal G11416: std_logic; attribute dont_touch of G11416: signal is true;
	signal G11417: std_logic; attribute dont_touch of G11417: signal is true;
	signal G11418: std_logic; attribute dont_touch of G11418: signal is true;
	signal G11419: std_logic; attribute dont_touch of G11419: signal is true;
	signal G11420: std_logic; attribute dont_touch of G11420: signal is true;
	signal G11421: std_logic; attribute dont_touch of G11421: signal is true;
	signal G11422: std_logic; attribute dont_touch of G11422: signal is true;
	signal G11423: std_logic; attribute dont_touch of G11423: signal is true;
	signal G11424: std_logic; attribute dont_touch of G11424: signal is true;
	signal G11425: std_logic; attribute dont_touch of G11425: signal is true;
	signal G11426: std_logic; attribute dont_touch of G11426: signal is true;
	signal G11427: std_logic; attribute dont_touch of G11427: signal is true;
	signal G11428: std_logic; attribute dont_touch of G11428: signal is true;
	signal G11429: std_logic; attribute dont_touch of G11429: signal is true;
	signal G11430: std_logic; attribute dont_touch of G11430: signal is true;
	signal G11431: std_logic; attribute dont_touch of G11431: signal is true;
	signal G11432: std_logic; attribute dont_touch of G11432: signal is true;
	signal G11433: std_logic; attribute dont_touch of G11433: signal is true;
	signal G11434: std_logic; attribute dont_touch of G11434: signal is true;
	signal G11435: std_logic; attribute dont_touch of G11435: signal is true;
	signal G11436: std_logic; attribute dont_touch of G11436: signal is true;
	signal G11437: std_logic; attribute dont_touch of G11437: signal is true;
	signal G11438: std_logic; attribute dont_touch of G11438: signal is true;
	signal G11439: std_logic; attribute dont_touch of G11439: signal is true;
	signal G11440: std_logic; attribute dont_touch of G11440: signal is true;
	signal G11441: std_logic; attribute dont_touch of G11441: signal is true;
	signal G11442: std_logic; attribute dont_touch of G11442: signal is true;
	signal G11443: std_logic; attribute dont_touch of G11443: signal is true;
	signal G11444: std_logic; attribute dont_touch of G11444: signal is true;
	signal G11445: std_logic; attribute dont_touch of G11445: signal is true;
	signal G11446: std_logic; attribute dont_touch of G11446: signal is true;
	signal G11447: std_logic; attribute dont_touch of G11447: signal is true;
	signal G11448: std_logic; attribute dont_touch of G11448: signal is true;
	signal G11449: std_logic; attribute dont_touch of G11449: signal is true;
	signal G11450: std_logic; attribute dont_touch of G11450: signal is true;
	signal G11451: std_logic; attribute dont_touch of G11451: signal is true;
	signal G11452: std_logic; attribute dont_touch of G11452: signal is true;
	signal G11453: std_logic; attribute dont_touch of G11453: signal is true;
	signal G11454: std_logic; attribute dont_touch of G11454: signal is true;
	signal G11455: std_logic; attribute dont_touch of G11455: signal is true;
	signal G11456: std_logic; attribute dont_touch of G11456: signal is true;
	signal G11457: std_logic; attribute dont_touch of G11457: signal is true;
	signal G11458: std_logic; attribute dont_touch of G11458: signal is true;
	signal G11459: std_logic; attribute dont_touch of G11459: signal is true;
	signal G11460: std_logic; attribute dont_touch of G11460: signal is true;
	signal G11461: std_logic; attribute dont_touch of G11461: signal is true;
	signal G11462: std_logic; attribute dont_touch of G11462: signal is true;
	signal G11463: std_logic; attribute dont_touch of G11463: signal is true;
	signal G11464: std_logic; attribute dont_touch of G11464: signal is true;
	signal G11465: std_logic; attribute dont_touch of G11465: signal is true;
	signal G11466: std_logic; attribute dont_touch of G11466: signal is true;
	signal G11467: std_logic; attribute dont_touch of G11467: signal is true;
	signal G11468: std_logic; attribute dont_touch of G11468: signal is true;
	signal G11469: std_logic; attribute dont_touch of G11469: signal is true;
	signal G11470: std_logic; attribute dont_touch of G11470: signal is true;
	signal G11471: std_logic; attribute dont_touch of G11471: signal is true;
	signal G11472: std_logic; attribute dont_touch of G11472: signal is true;
	signal G11473: std_logic; attribute dont_touch of G11473: signal is true;
	signal G11474: std_logic; attribute dont_touch of G11474: signal is true;
	signal G11475: std_logic; attribute dont_touch of G11475: signal is true;
	signal G11478: std_logic; attribute dont_touch of G11478: signal is true;
	signal G11479: std_logic; attribute dont_touch of G11479: signal is true;
	signal G11480: std_logic; attribute dont_touch of G11480: signal is true;
	signal G11481: std_logic; attribute dont_touch of G11481: signal is true;
	signal G11482: std_logic; attribute dont_touch of G11482: signal is true;
	signal G11483: std_logic; attribute dont_touch of G11483: signal is true;
	signal G11484: std_logic; attribute dont_touch of G11484: signal is true;
	signal G11485: std_logic; attribute dont_touch of G11485: signal is true;
	signal G11486: std_logic; attribute dont_touch of G11486: signal is true;
	signal G11487: std_logic; attribute dont_touch of G11487: signal is true;
	signal G11488: std_logic; attribute dont_touch of G11488: signal is true;
	signal G11490: std_logic; attribute dont_touch of G11490: signal is true;
	signal G11491: std_logic; attribute dont_touch of G11491: signal is true;
	signal G11492: std_logic; attribute dont_touch of G11492: signal is true;
	signal G11495: std_logic; attribute dont_touch of G11495: signal is true;
	signal G11496: std_logic; attribute dont_touch of G11496: signal is true;
	signal G11497: std_logic; attribute dont_touch of G11497: signal is true;
	signal G11498: std_logic; attribute dont_touch of G11498: signal is true;
	signal G11499: std_logic; attribute dont_touch of G11499: signal is true;
	signal G11500: std_logic; attribute dont_touch of G11500: signal is true;
	signal G11501: std_logic; attribute dont_touch of G11501: signal is true;
	signal G11502: std_logic; attribute dont_touch of G11502: signal is true;
	signal G11503: std_logic; attribute dont_touch of G11503: signal is true;
	signal G11504: std_logic; attribute dont_touch of G11504: signal is true;
	signal G11505: std_logic; attribute dont_touch of G11505: signal is true;
	signal G11506: std_logic; attribute dont_touch of G11506: signal is true;
	signal G11507: std_logic; attribute dont_touch of G11507: signal is true;
	signal G11508: std_logic; attribute dont_touch of G11508: signal is true;
	signal G11509: std_logic; attribute dont_touch of G11509: signal is true;
	signal G11510: std_logic; attribute dont_touch of G11510: signal is true;
	signal G11511: std_logic; attribute dont_touch of G11511: signal is true;
	signal G11512: std_logic; attribute dont_touch of G11512: signal is true;
	signal G11513: std_logic; attribute dont_touch of G11513: signal is true;
	signal G11514: std_logic; attribute dont_touch of G11514: signal is true;
	signal G11515: std_logic; attribute dont_touch of G11515: signal is true;
	signal G11518: std_logic; attribute dont_touch of G11518: signal is true;
	signal G11519: std_logic; attribute dont_touch of G11519: signal is true;
	signal G11538: std_logic; attribute dont_touch of G11538: signal is true;
	signal G11539: std_logic; attribute dont_touch of G11539: signal is true;
	signal G11540: std_logic; attribute dont_touch of G11540: signal is true;
	signal G11541: std_logic; attribute dont_touch of G11541: signal is true;
	signal G11542: std_logic; attribute dont_touch of G11542: signal is true;
	signal G11543: std_logic; attribute dont_touch of G11543: signal is true;
	signal G11544: std_logic; attribute dont_touch of G11544: signal is true;
	signal G11545: std_logic; attribute dont_touch of G11545: signal is true;
	signal G11546: std_logic; attribute dont_touch of G11546: signal is true;
	signal G11547: std_logic; attribute dont_touch of G11547: signal is true;
	signal G11548: std_logic; attribute dont_touch of G11548: signal is true;
	signal G11549: std_logic; attribute dont_touch of G11549: signal is true;
	signal G11550: std_logic; attribute dont_touch of G11550: signal is true;
	signal G11551: std_logic; attribute dont_touch of G11551: signal is true;
	signal G11552: std_logic; attribute dont_touch of G11552: signal is true;
	signal G11553: std_logic; attribute dont_touch of G11553: signal is true;
	signal G11554: std_logic; attribute dont_touch of G11554: signal is true;
	signal G11555: std_logic; attribute dont_touch of G11555: signal is true;
	signal G11556: std_logic; attribute dont_touch of G11556: signal is true;
	signal G11557: std_logic; attribute dont_touch of G11557: signal is true;
	signal G11558: std_logic; attribute dont_touch of G11558: signal is true;
	signal G11559: std_logic; attribute dont_touch of G11559: signal is true;
	signal G11560: std_logic; attribute dont_touch of G11560: signal is true;
	signal G11561: std_logic; attribute dont_touch of G11561: signal is true;
	signal G11571: std_logic; attribute dont_touch of G11571: signal is true;
	signal G11572: std_logic; attribute dont_touch of G11572: signal is true;
	signal G11573: std_logic; attribute dont_touch of G11573: signal is true;
	signal G11574: std_logic; attribute dont_touch of G11574: signal is true;
	signal G11575: std_logic; attribute dont_touch of G11575: signal is true;
	signal G11576: std_logic; attribute dont_touch of G11576: signal is true;
	signal G11577: std_logic; attribute dont_touch of G11577: signal is true;
	signal G11578: std_logic; attribute dont_touch of G11578: signal is true;
	signal G11579: std_logic; attribute dont_touch of G11579: signal is true;
	signal G11580: std_logic; attribute dont_touch of G11580: signal is true;
	signal G11581: std_logic; attribute dont_touch of G11581: signal is true;
	signal G11582: std_logic; attribute dont_touch of G11582: signal is true;
	signal G11583: std_logic; attribute dont_touch of G11583: signal is true;
	signal G11584: std_logic; attribute dont_touch of G11584: signal is true;
	signal G11585: std_logic; attribute dont_touch of G11585: signal is true;
	signal G11586: std_logic; attribute dont_touch of G11586: signal is true;
	signal G11587: std_logic; attribute dont_touch of G11587: signal is true;
	signal G11588: std_logic; attribute dont_touch of G11588: signal is true;
	signal G11589: std_logic; attribute dont_touch of G11589: signal is true;
	signal G11590: std_logic; attribute dont_touch of G11590: signal is true;
	signal G11591: std_logic; attribute dont_touch of G11591: signal is true;
	signal G11592: std_logic; attribute dont_touch of G11592: signal is true;
	signal G11593: std_logic; attribute dont_touch of G11593: signal is true;
	signal G11594: std_logic; attribute dont_touch of G11594: signal is true;
	signal G11595: std_logic; attribute dont_touch of G11595: signal is true;
	signal G11596: std_logic; attribute dont_touch of G11596: signal is true;
	signal G11597: std_logic; attribute dont_touch of G11597: signal is true;
	signal G11598: std_logic; attribute dont_touch of G11598: signal is true;
	signal G11599: std_logic; attribute dont_touch of G11599: signal is true;
	signal G11600: std_logic; attribute dont_touch of G11600: signal is true;
	signal G11601: std_logic; attribute dont_touch of G11601: signal is true;
	signal G11602: std_logic; attribute dont_touch of G11602: signal is true;
	signal G11603: std_logic; attribute dont_touch of G11603: signal is true;
	signal G11604: std_logic; attribute dont_touch of G11604: signal is true;
	signal G11605: std_logic; attribute dont_touch of G11605: signal is true;
	signal G11606: std_logic; attribute dont_touch of G11606: signal is true;
	signal G11607: std_logic; attribute dont_touch of G11607: signal is true;
	signal G11608: std_logic; attribute dont_touch of G11608: signal is true;
	signal G11609: std_logic; attribute dont_touch of G11609: signal is true;
	signal G11610: std_logic; attribute dont_touch of G11610: signal is true;
	signal G11611: std_logic; attribute dont_touch of G11611: signal is true;
	signal G11612: std_logic; attribute dont_touch of G11612: signal is true;
	signal G11613: std_logic; attribute dont_touch of G11613: signal is true;
	signal G11614: std_logic; attribute dont_touch of G11614: signal is true;
	signal G11615: std_logic; attribute dont_touch of G11615: signal is true;
	signal G11616: std_logic; attribute dont_touch of G11616: signal is true;
	signal G11617: std_logic; attribute dont_touch of G11617: signal is true;
	signal G11618: std_logic; attribute dont_touch of G11618: signal is true;
	signal G11619: std_logic; attribute dont_touch of G11619: signal is true;
	signal G11620: std_logic; attribute dont_touch of G11620: signal is true;
	signal G11621: std_logic; attribute dont_touch of G11621: signal is true;
	signal G11622: std_logic; attribute dont_touch of G11622: signal is true;
	signal G11623: std_logic; attribute dont_touch of G11623: signal is true;
	signal G11624: std_logic; attribute dont_touch of G11624: signal is true;
	signal G11625: std_logic; attribute dont_touch of G11625: signal is true;
	signal G11626: std_logic; attribute dont_touch of G11626: signal is true;
	signal G11627: std_logic; attribute dont_touch of G11627: signal is true;
	signal G11628: std_logic; attribute dont_touch of G11628: signal is true;
	signal G11629: std_logic; attribute dont_touch of G11629: signal is true;
	signal G11630: std_logic; attribute dont_touch of G11630: signal is true;
	signal G11631: std_logic; attribute dont_touch of G11631: signal is true;
	signal G11632: std_logic; attribute dont_touch of G11632: signal is true;
	signal G11633: std_logic; attribute dont_touch of G11633: signal is true;
	signal G11634: std_logic; attribute dont_touch of G11634: signal is true;
	signal G11635: std_logic; attribute dont_touch of G11635: signal is true;
	signal G11636: std_logic; attribute dont_touch of G11636: signal is true;
	signal G11637: std_logic; attribute dont_touch of G11637: signal is true;
	signal G11638: std_logic; attribute dont_touch of G11638: signal is true;
	signal G11639: std_logic; attribute dont_touch of G11639: signal is true;
	signal G11640: std_logic; attribute dont_touch of G11640: signal is true;
	signal G11641: std_logic; attribute dont_touch of G11641: signal is true;
	signal G11642: std_logic; attribute dont_touch of G11642: signal is true;
	signal G11643: std_logic; attribute dont_touch of G11643: signal is true;
	signal G11644: std_logic; attribute dont_touch of G11644: signal is true;
	signal G11645: std_logic; attribute dont_touch of G11645: signal is true;
	signal G11646: std_logic; attribute dont_touch of G11646: signal is true;
	signal G11647: std_logic; attribute dont_touch of G11647: signal is true;
	signal G11648: std_logic; attribute dont_touch of G11648: signal is true;
	signal G11649: std_logic; attribute dont_touch of G11649: signal is true;
	signal G11650: std_logic; attribute dont_touch of G11650: signal is true;
	signal G11651: std_logic; attribute dont_touch of G11651: signal is true;
	signal G11652: std_logic; attribute dont_touch of G11652: signal is true;
	signal G11653: std_logic; attribute dont_touch of G11653: signal is true;
	signal G11654: std_logic; attribute dont_touch of G11654: signal is true;
	signal G11655: std_logic; attribute dont_touch of G11655: signal is true;
	signal G11656: std_logic; attribute dont_touch of G11656: signal is true;
	signal G11657: std_logic; attribute dont_touch of G11657: signal is true;
	signal I4777: std_logic; attribute dont_touch of I4777: signal is true;
	signal I4780: std_logic; attribute dont_touch of I4780: signal is true;
	signal I4783: std_logic; attribute dont_touch of I4783: signal is true;
	signal I4786: std_logic; attribute dont_touch of I4786: signal is true;
	signal I4820: std_logic; attribute dont_touch of I4820: signal is true;
	signal I4850: std_logic; attribute dont_touch of I4850: signal is true;
	signal I4859: std_logic; attribute dont_touch of I4859: signal is true;
	signal I4866: std_logic; attribute dont_touch of I4866: signal is true;
	signal I4869: std_logic; attribute dont_touch of I4869: signal is true;
	signal I4873: std_logic; attribute dont_touch of I4873: signal is true;
	signal I4876: std_logic; attribute dont_touch of I4876: signal is true;
	signal I4879: std_logic; attribute dont_touch of I4879: signal is true;
	signal I4883: std_logic; attribute dont_touch of I4883: signal is true;
	signal I4886: std_logic; attribute dont_touch of I4886: signal is true;
	signal I4891: std_logic; attribute dont_touch of I4891: signal is true;
	signal I4894: std_logic; attribute dont_touch of I4894: signal is true;
	signal I4900: std_logic; attribute dont_touch of I4900: signal is true;
	signal I4903: std_logic; attribute dont_touch of I4903: signal is true;
	signal I4906: std_logic; attribute dont_touch of I4906: signal is true;
	signal I4910: std_logic; attribute dont_touch of I4910: signal is true;
	signal I4911: std_logic; attribute dont_touch of I4911: signal is true;
	signal I4912: std_logic; attribute dont_touch of I4912: signal is true;
	signal I4917: std_logic; attribute dont_touch of I4917: signal is true;
	signal I4920: std_logic; attribute dont_touch of I4920: signal is true;
	signal I4924: std_logic; attribute dont_touch of I4924: signal is true;
	signal I4928: std_logic; attribute dont_touch of I4928: signal is true;
	signal I4929: std_logic; attribute dont_touch of I4929: signal is true;
	signal I4930: std_logic; attribute dont_touch of I4930: signal is true;
	signal I4935: std_logic; attribute dont_touch of I4935: signal is true;
	signal I4938: std_logic; attribute dont_touch of I4938: signal is true;
	signal I4941: std_logic; attribute dont_touch of I4941: signal is true;
	signal I4942: std_logic; attribute dont_touch of I4942: signal is true;
	signal I4943: std_logic; attribute dont_touch of I4943: signal is true;
	signal I4948: std_logic; attribute dont_touch of I4948: signal is true;
	signal I4951: std_logic; attribute dont_touch of I4951: signal is true;
	signal I4954: std_logic; attribute dont_touch of I4954: signal is true;
	signal I4955: std_logic; attribute dont_touch of I4955: signal is true;
	signal I4956: std_logic; attribute dont_touch of I4956: signal is true;
	signal I4961: std_logic; attribute dont_touch of I4961: signal is true;
	signal I4964: std_logic; attribute dont_touch of I4964: signal is true;
	signal I4965: std_logic; attribute dont_touch of I4965: signal is true;
	signal I4966: std_logic; attribute dont_touch of I4966: signal is true;
	signal I4971: std_logic; attribute dont_touch of I4971: signal is true;
	signal I4972: std_logic; attribute dont_touch of I4972: signal is true;
	signal I4973: std_logic; attribute dont_touch of I4973: signal is true;
	signal I4978: std_logic; attribute dont_touch of I4978: signal is true;
	signal I4979: std_logic; attribute dont_touch of I4979: signal is true;
	signal I4980: std_logic; attribute dont_touch of I4980: signal is true;
	signal I4985: std_logic; attribute dont_touch of I4985: signal is true;
	signal I4986: std_logic; attribute dont_touch of I4986: signal is true;
	signal I4987: std_logic; attribute dont_touch of I4987: signal is true;
	signal I4992: std_logic; attribute dont_touch of I4992: signal is true;
	signal I4995: std_logic; attribute dont_touch of I4995: signal is true;
	signal I4996: std_logic; attribute dont_touch of I4996: signal is true;
	signal I4997: std_logic; attribute dont_touch of I4997: signal is true;
	signal I5002: std_logic; attribute dont_touch of I5002: signal is true;
	signal I5005: std_logic; attribute dont_touch of I5005: signal is true;
	signal I5006: std_logic; attribute dont_touch of I5006: signal is true;
	signal I5007: std_logic; attribute dont_touch of I5007: signal is true;
	signal I5013: std_logic; attribute dont_touch of I5013: signal is true;
	signal I5014: std_logic; attribute dont_touch of I5014: signal is true;
	signal I5015: std_logic; attribute dont_touch of I5015: signal is true;
	signal I5020: std_logic; attribute dont_touch of I5020: signal is true;
	signal I5023: std_logic; attribute dont_touch of I5023: signal is true;
	signal I5024: std_logic; attribute dont_touch of I5024: signal is true;
	signal I5025: std_logic; attribute dont_touch of I5025: signal is true;
	signal I5031: std_logic; attribute dont_touch of I5031: signal is true;
	signal I5034: std_logic; attribute dont_touch of I5034: signal is true;
	signal I5035: std_logic; attribute dont_touch of I5035: signal is true;
	signal I5036: std_logic; attribute dont_touch of I5036: signal is true;
	signal I5041: std_logic; attribute dont_touch of I5041: signal is true;
	signal I5044: std_logic; attribute dont_touch of I5044: signal is true;
	signal I5047: std_logic; attribute dont_touch of I5047: signal is true;
	signal I5050: std_logic; attribute dont_touch of I5050: signal is true;
	signal I5053: std_logic; attribute dont_touch of I5053: signal is true;
	signal I5057: std_logic; attribute dont_touch of I5057: signal is true;
	signal I5060: std_logic; attribute dont_touch of I5060: signal is true;
	signal I5064: std_logic; attribute dont_touch of I5064: signal is true;
	signal I5067: std_logic; attribute dont_touch of I5067: signal is true;
	signal I5070: std_logic; attribute dont_touch of I5070: signal is true;
	signal I5073: std_logic; attribute dont_touch of I5073: signal is true;
	signal I5077: std_logic; attribute dont_touch of I5077: signal is true;
	signal I5080: std_logic; attribute dont_touch of I5080: signal is true;
	signal I5084: std_logic; attribute dont_touch of I5084: signal is true;
	signal I5085: std_logic; attribute dont_touch of I5085: signal is true;
	signal I5089: std_logic; attribute dont_touch of I5089: signal is true;
	signal I5092: std_logic; attribute dont_touch of I5092: signal is true;
	signal I5095: std_logic; attribute dont_touch of I5095: signal is true;
	signal I5098: std_logic; attribute dont_touch of I5098: signal is true;
	signal I5101: std_logic; attribute dont_touch of I5101: signal is true;
	signal I5104: std_logic; attribute dont_touch of I5104: signal is true;
	signal I5105: std_logic; attribute dont_touch of I5105: signal is true;
	signal I5106: std_logic; attribute dont_touch of I5106: signal is true;
	signal I5111: std_logic; attribute dont_touch of I5111: signal is true;
	signal I5116: std_logic; attribute dont_touch of I5116: signal is true;
	signal I5120: std_logic; attribute dont_touch of I5120: signal is true;
	signal I5126: std_logic; attribute dont_touch of I5126: signal is true;
	signal I5127: std_logic; attribute dont_touch of I5127: signal is true;
	signal I5128: std_logic; attribute dont_touch of I5128: signal is true;
	signal I5135: std_logic; attribute dont_touch of I5135: signal is true;
	signal I5136: std_logic; attribute dont_touch of I5136: signal is true;
	signal I5137: std_logic; attribute dont_touch of I5137: signal is true;
	signal I5142: std_logic; attribute dont_touch of I5142: signal is true;
	signal I5149: std_logic; attribute dont_touch of I5149: signal is true;
	signal I5164: std_logic; attribute dont_touch of I5164: signal is true;
	signal I5165: std_logic; attribute dont_touch of I5165: signal is true;
	signal I5166: std_logic; attribute dont_touch of I5166: signal is true;
	signal I5171: std_logic; attribute dont_touch of I5171: signal is true;
	signal I5174: std_logic; attribute dont_touch of I5174: signal is true;
	signal I5184: std_logic; attribute dont_touch of I5184: signal is true;
	signal I5185: std_logic; attribute dont_touch of I5185: signal is true;
	signal I5186: std_logic; attribute dont_touch of I5186: signal is true;
	signal I5192: std_logic; attribute dont_touch of I5192: signal is true;
	signal I5198: std_logic; attribute dont_touch of I5198: signal is true;
	signal I5202: std_logic; attribute dont_touch of I5202: signal is true;
	signal I5203: std_logic; attribute dont_touch of I5203: signal is true;
	signal I5204: std_logic; attribute dont_touch of I5204: signal is true;
	signal I5210: std_logic; attribute dont_touch of I5210: signal is true;
	signal I5218: std_logic; attribute dont_touch of I5218: signal is true;
	signal I5221: std_logic; attribute dont_touch of I5221: signal is true;
	signal I5224: std_logic; attribute dont_touch of I5224: signal is true;
	signal I5229: std_logic; attribute dont_touch of I5229: signal is true;
	signal I5230: std_logic; attribute dont_touch of I5230: signal is true;
	signal I5231: std_logic; attribute dont_touch of I5231: signal is true;
	signal I5237: std_logic; attribute dont_touch of I5237: signal is true;
	signal I5240: std_logic; attribute dont_touch of I5240: signal is true;
	signal I5245: std_logic; attribute dont_touch of I5245: signal is true;
	signal I5248: std_logic; attribute dont_touch of I5248: signal is true;
	signal I5251: std_logic; attribute dont_touch of I5251: signal is true;
	signal I5254: std_logic; attribute dont_touch of I5254: signal is true;
	signal I5258: std_logic; attribute dont_touch of I5258: signal is true;
	signal I5263: std_logic; attribute dont_touch of I5263: signal is true;
	signal I5264: std_logic; attribute dont_touch of I5264: signal is true;
	signal I5265: std_logic; attribute dont_touch of I5265: signal is true;
	signal I5271: std_logic; attribute dont_touch of I5271: signal is true;
	signal I5276: std_logic; attribute dont_touch of I5276: signal is true;
	signal I5279: std_logic; attribute dont_touch of I5279: signal is true;
	signal I5282: std_logic; attribute dont_touch of I5282: signal is true;
	signal I5283: std_logic; attribute dont_touch of I5283: signal is true;
	signal I5284: std_logic; attribute dont_touch of I5284: signal is true;
	signal I5289: std_logic; attribute dont_touch of I5289: signal is true;
	signal I5292: std_logic; attribute dont_touch of I5292: signal is true;
	signal I5295: std_logic; attribute dont_touch of I5295: signal is true;
	signal I5296: std_logic; attribute dont_touch of I5296: signal is true;
	signal I5297: std_logic; attribute dont_touch of I5297: signal is true;
	signal I5304: std_logic; attribute dont_touch of I5304: signal is true;
	signal I5308: std_logic; attribute dont_touch of I5308: signal is true;
	signal I5311: std_logic; attribute dont_touch of I5311: signal is true;
	signal I5315: std_logic; attribute dont_touch of I5315: signal is true;
	signal I5316: std_logic; attribute dont_touch of I5316: signal is true;
	signal I5317: std_logic; attribute dont_touch of I5317: signal is true;
	signal I5323: std_logic; attribute dont_touch of I5323: signal is true;
	signal I5324: std_logic; attribute dont_touch of I5324: signal is true;
	signal I5325: std_logic; attribute dont_touch of I5325: signal is true;
	signal I5332: std_logic; attribute dont_touch of I5332: signal is true;
	signal I5336: std_logic; attribute dont_touch of I5336: signal is true;
	signal I5341: std_logic; attribute dont_touch of I5341: signal is true;
	signal I5342: std_logic; attribute dont_touch of I5342: signal is true;
	signal I5343: std_logic; attribute dont_touch of I5343: signal is true;
	signal I5348: std_logic; attribute dont_touch of I5348: signal is true;
	signal I5351: std_logic; attribute dont_touch of I5351: signal is true;
	signal I5352: std_logic; attribute dont_touch of I5352: signal is true;
	signal I5357: std_logic; attribute dont_touch of I5357: signal is true;
	signal I5358: std_logic; attribute dont_touch of I5358: signal is true;
	signal I5363: std_logic; attribute dont_touch of I5363: signal is true;
	signal I5366: std_logic; attribute dont_touch of I5366: signal is true;
	signal I5371: std_logic; attribute dont_touch of I5371: signal is true;
	signal I5372: std_logic; attribute dont_touch of I5372: signal is true;
	signal I5373: std_logic; attribute dont_touch of I5373: signal is true;
	signal I5378: std_logic; attribute dont_touch of I5378: signal is true;
	signal I5383: std_logic; attribute dont_touch of I5383: signal is true;
	signal I5388: std_logic; attribute dont_touch of I5388: signal is true;
	signal I5391: std_logic; attribute dont_touch of I5391: signal is true;
	signal I5395: std_logic; attribute dont_touch of I5395: signal is true;
	signal I5399: std_logic; attribute dont_touch of I5399: signal is true;
	signal I5403: std_logic; attribute dont_touch of I5403: signal is true;
	signal I5406: std_logic; attribute dont_touch of I5406: signal is true;
	signal I5410: std_logic; attribute dont_touch of I5410: signal is true;
	signal I5414: std_logic; attribute dont_touch of I5414: signal is true;
	signal I5418: std_logic; attribute dont_touch of I5418: signal is true;
	signal I5421: std_logic; attribute dont_touch of I5421: signal is true;
	signal I5424: std_logic; attribute dont_touch of I5424: signal is true;
	signal I5427: std_logic; attribute dont_touch of I5427: signal is true;
	signal I5430: std_logic; attribute dont_touch of I5430: signal is true;
	signal I5435: std_logic; attribute dont_touch of I5435: signal is true;
	signal I5438: std_logic; attribute dont_touch of I5438: signal is true;
	signal I5441: std_logic; attribute dont_touch of I5441: signal is true;
	signal I5445: std_logic; attribute dont_touch of I5445: signal is true;
	signal I5449: std_logic; attribute dont_touch of I5449: signal is true;
	signal I5450: std_logic; attribute dont_touch of I5450: signal is true;
	signal I5451: std_logic; attribute dont_touch of I5451: signal is true;
	signal I5459: std_logic; attribute dont_touch of I5459: signal is true;
	signal I5460: std_logic; attribute dont_touch of I5460: signal is true;
	signal I5461: std_logic; attribute dont_touch of I5461: signal is true;
	signal I5468: std_logic; attribute dont_touch of I5468: signal is true;
	signal I5469: std_logic; attribute dont_touch of I5469: signal is true;
	signal I5470: std_logic; attribute dont_touch of I5470: signal is true;
	signal I5475: std_logic; attribute dont_touch of I5475: signal is true;
	signal I5478: std_logic; attribute dont_touch of I5478: signal is true;
	signal I5484: std_logic; attribute dont_touch of I5484: signal is true;
	signal I5485: std_logic; attribute dont_touch of I5485: signal is true;
	signal I5486: std_logic; attribute dont_touch of I5486: signal is true;
	signal I5494: std_logic; attribute dont_touch of I5494: signal is true;
	signal I5497: std_logic; attribute dont_touch of I5497: signal is true;
	signal I5500: std_logic; attribute dont_touch of I5500: signal is true;
	signal I5501: std_logic; attribute dont_touch of I5501: signal is true;
	signal I5502: std_logic; attribute dont_touch of I5502: signal is true;
	signal I5510: std_logic; attribute dont_touch of I5510: signal is true;
	signal I5513: std_logic; attribute dont_touch of I5513: signal is true;
	signal I5516: std_logic; attribute dont_touch of I5516: signal is true;
	signal I5517: std_logic; attribute dont_touch of I5517: signal is true;
	signal I5518: std_logic; attribute dont_touch of I5518: signal is true;
	signal I5525: std_logic; attribute dont_touch of I5525: signal is true;
	signal I5528: std_logic; attribute dont_touch of I5528: signal is true;
	signal I5529: std_logic; attribute dont_touch of I5529: signal is true;
	signal I5530: std_logic; attribute dont_touch of I5530: signal is true;
	signal I5538: std_logic; attribute dont_touch of I5538: signal is true;
	signal I5539: std_logic; attribute dont_touch of I5539: signal is true;
	signal I5540: std_logic; attribute dont_touch of I5540: signal is true;
	signal I5549: std_logic; attribute dont_touch of I5549: signal is true;
	signal I5555: std_logic; attribute dont_touch of I5555: signal is true;
	signal I5561: std_logic; attribute dont_touch of I5561: signal is true;
	signal I5565: std_logic; attribute dont_touch of I5565: signal is true;
	signal I5570: std_logic; attribute dont_touch of I5570: signal is true;
	signal I5571: std_logic; attribute dont_touch of I5571: signal is true;
	signal I5576: std_logic; attribute dont_touch of I5576: signal is true;
	signal I5579: std_logic; attribute dont_touch of I5579: signal is true;
	signal I5584: std_logic; attribute dont_touch of I5584: signal is true;
	signal I5588: std_logic; attribute dont_touch of I5588: signal is true;
	signal I5591: std_logic; attribute dont_touch of I5591: signal is true;
	signal I5592: std_logic; attribute dont_touch of I5592: signal is true;
	signal I5593: std_logic; attribute dont_touch of I5593: signal is true;
	signal I5599: std_logic; attribute dont_touch of I5599: signal is true;
	signal I5600: std_logic; attribute dont_touch of I5600: signal is true;
	signal I5604: std_logic; attribute dont_touch of I5604: signal is true;
	signal I5605: std_logic; attribute dont_touch of I5605: signal is true;
	signal I5606: std_logic; attribute dont_touch of I5606: signal is true;
	signal I5611: std_logic; attribute dont_touch of I5611: signal is true;
	signal I5612: std_logic; attribute dont_touch of I5612: signal is true;
	signal I5613: std_logic; attribute dont_touch of I5613: signal is true;
	signal I5618: std_logic; attribute dont_touch of I5618: signal is true;
	signal I5619: std_logic; attribute dont_touch of I5619: signal is true;
	signal I5620: std_logic; attribute dont_touch of I5620: signal is true;
	signal I5626: std_logic; attribute dont_touch of I5626: signal is true;
	signal I5629: std_logic; attribute dont_touch of I5629: signal is true;
	signal I5632: std_logic; attribute dont_touch of I5632: signal is true;
	signal I5638: std_logic; attribute dont_touch of I5638: signal is true;
	signal I5641: std_logic; attribute dont_touch of I5641: signal is true;
	signal I5646: std_logic; attribute dont_touch of I5646: signal is true;
	signal I5649: std_logic; attribute dont_touch of I5649: signal is true;
	signal I5652: std_logic; attribute dont_touch of I5652: signal is true;
	signal I5655: std_logic; attribute dont_touch of I5655: signal is true;
	signal I5658: std_logic; attribute dont_touch of I5658: signal is true;
	signal I5662: std_logic; attribute dont_touch of I5662: signal is true;
	signal I5667: std_logic; attribute dont_touch of I5667: signal is true;
	signal I5672: std_logic; attribute dont_touch of I5672: signal is true;
	signal I5675: std_logic; attribute dont_touch of I5675: signal is true;
	signal I5676: std_logic; attribute dont_touch of I5676: signal is true;
	signal I5677: std_logic; attribute dont_touch of I5677: signal is true;
	signal I5684: std_logic; attribute dont_touch of I5684: signal is true;
	signal I5689: std_logic; attribute dont_touch of I5689: signal is true;
	signal I5690: std_logic; attribute dont_touch of I5690: signal is true;
	signal I5695: std_logic; attribute dont_touch of I5695: signal is true;
	signal I5704: std_logic; attribute dont_touch of I5704: signal is true;
	signal I5707: std_logic; attribute dont_touch of I5707: signal is true;
	signal I5710: std_logic; attribute dont_touch of I5710: signal is true;
	signal I5713: std_logic; attribute dont_touch of I5713: signal is true;
	signal I5716: std_logic; attribute dont_touch of I5716: signal is true;
	signal I5719: std_logic; attribute dont_touch of I5719: signal is true;
	signal I5722: std_logic; attribute dont_touch of I5722: signal is true;
	signal I5725: std_logic; attribute dont_touch of I5725: signal is true;
	signal I5728: std_logic; attribute dont_touch of I5728: signal is true;
	signal I5731: std_logic; attribute dont_touch of I5731: signal is true;
	signal I5734: std_logic; attribute dont_touch of I5734: signal is true;
	signal I5737: std_logic; attribute dont_touch of I5737: signal is true;
	signal I5740: std_logic; attribute dont_touch of I5740: signal is true;
	signal I5751: std_logic; attribute dont_touch of I5751: signal is true;
	signal I5754: std_logic; attribute dont_touch of I5754: signal is true;
	signal I5765: std_logic; attribute dont_touch of I5765: signal is true;
	signal I5789: std_logic; attribute dont_touch of I5789: signal is true;
	signal I5792: std_logic; attribute dont_touch of I5792: signal is true;
	signal I5795: std_logic; attribute dont_touch of I5795: signal is true;
	signal I5798: std_logic; attribute dont_touch of I5798: signal is true;
	signal I5801: std_logic; attribute dont_touch of I5801: signal is true;
	signal I5804: std_logic; attribute dont_touch of I5804: signal is true;
	signal I5805: std_logic; attribute dont_touch of I5805: signal is true;
	signal I5809: std_logic; attribute dont_touch of I5809: signal is true;
	signal I5812: std_logic; attribute dont_touch of I5812: signal is true;
	signal I5815: std_logic; attribute dont_touch of I5815: signal is true;
	signal I5818: std_logic; attribute dont_touch of I5818: signal is true;
	signal I5821: std_logic; attribute dont_touch of I5821: signal is true;
	signal I5824: std_logic; attribute dont_touch of I5824: signal is true;
	signal I5827: std_logic; attribute dont_touch of I5827: signal is true;
	signal I5830: std_logic; attribute dont_touch of I5830: signal is true;
	signal I5833: std_logic; attribute dont_touch of I5833: signal is true;
	signal I5837: std_logic; attribute dont_touch of I5837: signal is true;
	signal I5840: std_logic; attribute dont_touch of I5840: signal is true;
	signal I5843: std_logic; attribute dont_touch of I5843: signal is true;
	signal I5847: std_logic; attribute dont_touch of I5847: signal is true;
	signal I5850: std_logic; attribute dont_touch of I5850: signal is true;
	signal I5854: std_logic; attribute dont_touch of I5854: signal is true;
	signal I5858: std_logic; attribute dont_touch of I5858: signal is true;
	signal I5862: std_logic; attribute dont_touch of I5862: signal is true;
	signal I5865: std_logic; attribute dont_touch of I5865: signal is true;
	signal I5866: std_logic; attribute dont_touch of I5866: signal is true;
	signal I5867: std_logic; attribute dont_touch of I5867: signal is true;
	signal I5878: std_logic; attribute dont_touch of I5878: signal is true;
	signal I5879: std_logic; attribute dont_touch of I5879: signal is true;
	signal I5880: std_logic; attribute dont_touch of I5880: signal is true;
	signal I5886: std_logic; attribute dont_touch of I5886: signal is true;
	signal I5887: std_logic; attribute dont_touch of I5887: signal is true;
	signal I5891: std_logic; attribute dont_touch of I5891: signal is true;
	signal I5892: std_logic; attribute dont_touch of I5892: signal is true;
	signal I5893: std_logic; attribute dont_touch of I5893: signal is true;
	signal I5909: std_logic; attribute dont_touch of I5909: signal is true;
	signal I5913: std_logic; attribute dont_touch of I5913: signal is true;
	signal I5916: std_logic; attribute dont_touch of I5916: signal is true;
	signal I5919: std_logic; attribute dont_touch of I5919: signal is true;
	signal I5922: std_logic; attribute dont_touch of I5922: signal is true;
	signal I5926: std_logic; attribute dont_touch of I5926: signal is true;
	signal I5929: std_logic; attribute dont_touch of I5929: signal is true;
	signal I5932: std_logic; attribute dont_touch of I5932: signal is true;
	signal I5935: std_logic; attribute dont_touch of I5935: signal is true;
	signal I5940: std_logic; attribute dont_touch of I5940: signal is true;
	signal I5943: std_logic; attribute dont_touch of I5943: signal is true;
	signal I5946: std_logic; attribute dont_touch of I5946: signal is true;
	signal I5949: std_logic; attribute dont_touch of I5949: signal is true;
	signal I5952: std_logic; attribute dont_touch of I5952: signal is true;
	signal I5957: std_logic; attribute dont_touch of I5957: signal is true;
	signal I5960: std_logic; attribute dont_touch of I5960: signal is true;
	signal I5963: std_logic; attribute dont_touch of I5963: signal is true;
	signal I5966: std_logic; attribute dont_touch of I5966: signal is true;
	signal I5970: std_logic; attribute dont_touch of I5970: signal is true;
	signal I5973: std_logic; attribute dont_touch of I5973: signal is true;
	signal I5976: std_logic; attribute dont_touch of I5976: signal is true;
	signal I5979: std_logic; attribute dont_touch of I5979: signal is true;
	signal I5982: std_logic; attribute dont_touch of I5982: signal is true;
	signal I5986: std_logic; attribute dont_touch of I5986: signal is true;
	signal I5989: std_logic; attribute dont_touch of I5989: signal is true;
	signal I5992: std_logic; attribute dont_touch of I5992: signal is true;
	signal I5995: std_logic; attribute dont_touch of I5995: signal is true;
	signal I5998: std_logic; attribute dont_touch of I5998: signal is true;
	signal I6001: std_logic; attribute dont_touch of I6001: signal is true;
	signal I6007: std_logic; attribute dont_touch of I6007: signal is true;
	signal I6010: std_logic; attribute dont_touch of I6010: signal is true;
	signal I6013: std_logic; attribute dont_touch of I6013: signal is true;
	signal I6016: std_logic; attribute dont_touch of I6016: signal is true;
	signal I6019: std_logic; attribute dont_touch of I6019: signal is true;
	signal I6022: std_logic; attribute dont_touch of I6022: signal is true;
	signal I6025: std_logic; attribute dont_touch of I6025: signal is true;
	signal I6028: std_logic; attribute dont_touch of I6028: signal is true;
	signal I6031: std_logic; attribute dont_touch of I6031: signal is true;
	signal I6034: std_logic; attribute dont_touch of I6034: signal is true;
	signal I6037: std_logic; attribute dont_touch of I6037: signal is true;
	signal I6040: std_logic; attribute dont_touch of I6040: signal is true;
	signal I6043: std_logic; attribute dont_touch of I6043: signal is true;
	signal I6046: std_logic; attribute dont_touch of I6046: signal is true;
	signal I6049: std_logic; attribute dont_touch of I6049: signal is true;
	signal I6052: std_logic; attribute dont_touch of I6052: signal is true;
	signal I6055: std_logic; attribute dont_touch of I6055: signal is true;
	signal I6061: std_logic; attribute dont_touch of I6061: signal is true;
	signal I6065: std_logic; attribute dont_touch of I6065: signal is true;
	signal I6068: std_logic; attribute dont_touch of I6068: signal is true;
	signal I6071: std_logic; attribute dont_touch of I6071: signal is true;
	signal I6074: std_logic; attribute dont_touch of I6074: signal is true;
	signal I6077: std_logic; attribute dont_touch of I6077: signal is true;
	signal I6080: std_logic; attribute dont_touch of I6080: signal is true;
	signal I6085: std_logic; attribute dont_touch of I6085: signal is true;
	signal I6088: std_logic; attribute dont_touch of I6088: signal is true;
	signal I6091: std_logic; attribute dont_touch of I6091: signal is true;
	signal I6094: std_logic; attribute dont_touch of I6094: signal is true;
	signal I6097: std_logic; attribute dont_touch of I6097: signal is true;
	signal I6102: std_logic; attribute dont_touch of I6102: signal is true;
	signal I6106: std_logic; attribute dont_touch of I6106: signal is true;
	signal I6109: std_logic; attribute dont_touch of I6109: signal is true;
	signal I6110: std_logic; attribute dont_touch of I6110: signal is true;
	signal I6111: std_logic; attribute dont_touch of I6111: signal is true;
	signal I6118: std_logic; attribute dont_touch of I6118: signal is true;
	signal I6121: std_logic; attribute dont_touch of I6121: signal is true;
	signal I6124: std_logic; attribute dont_touch of I6124: signal is true;
	signal I6125: std_logic; attribute dont_touch of I6125: signal is true;
	signal I6126: std_logic; attribute dont_touch of I6126: signal is true;
	signal I6133: std_logic; attribute dont_touch of I6133: signal is true;
	signal I6136: std_logic; attribute dont_touch of I6136: signal is true;
	signal I6137: std_logic; attribute dont_touch of I6137: signal is true;
	signal I6138: std_logic; attribute dont_touch of I6138: signal is true;
	signal I6143: std_logic; attribute dont_touch of I6143: signal is true;
	signal I6144: std_logic; attribute dont_touch of I6144: signal is true;
	signal I6145: std_logic; attribute dont_touch of I6145: signal is true;
	signal I6150: std_logic; attribute dont_touch of I6150: signal is true;
	signal I6156: std_logic; attribute dont_touch of I6156: signal is true;
	signal I6159: std_logic; attribute dont_touch of I6159: signal is true;
	signal I6163: std_logic; attribute dont_touch of I6163: signal is true;
	signal I6166: std_logic; attribute dont_touch of I6166: signal is true;
	signal I6167: std_logic; attribute dont_touch of I6167: signal is true;
	signal I6168: std_logic; attribute dont_touch of I6168: signal is true;
	signal I6173: std_logic; attribute dont_touch of I6173: signal is true;
	signal I6176: std_logic; attribute dont_touch of I6176: signal is true;
	signal I6177: std_logic; attribute dont_touch of I6177: signal is true;
	signal I6178: std_logic; attribute dont_touch of I6178: signal is true;
	signal I6183: std_logic; attribute dont_touch of I6183: signal is true;
	signal I6186: std_logic; attribute dont_touch of I6186: signal is true;
	signal I6187: std_logic; attribute dont_touch of I6187: signal is true;
	signal I6188: std_logic; attribute dont_touch of I6188: signal is true;
	signal I6193: std_logic; attribute dont_touch of I6193: signal is true;
	signal I6196: std_logic; attribute dont_touch of I6196: signal is true;
	signal I6199: std_logic; attribute dont_touch of I6199: signal is true;
	signal I6200: std_logic; attribute dont_touch of I6200: signal is true;
	signal I6201: std_logic; attribute dont_touch of I6201: signal is true;
	signal I6207: std_logic; attribute dont_touch of I6207: signal is true;
	signal I6208: std_logic; attribute dont_touch of I6208: signal is true;
	signal I6209: std_logic; attribute dont_touch of I6209: signal is true;
	signal I6217: std_logic; attribute dont_touch of I6217: signal is true;
	signal I6220: std_logic; attribute dont_touch of I6220: signal is true;
	signal I6224: std_logic; attribute dont_touch of I6224: signal is true;
	signal I6225: std_logic; attribute dont_touch of I6225: signal is true;
	signal I6226: std_logic; attribute dont_touch of I6226: signal is true;
	signal I6233: std_logic; attribute dont_touch of I6233: signal is true;
	signal I6240: std_logic; attribute dont_touch of I6240: signal is true;
	signal I6247: std_logic; attribute dont_touch of I6247: signal is true;
	signal I6256: std_logic; attribute dont_touch of I6256: signal is true;
	signal I6260: std_logic; attribute dont_touch of I6260: signal is true;
	signal I6264: std_logic; attribute dont_touch of I6264: signal is true;
	signal I6273: std_logic; attribute dont_touch of I6273: signal is true;
	signal I6277: std_logic; attribute dont_touch of I6277: signal is true;
	signal I6282: std_logic; attribute dont_touch of I6282: signal is true;
	signal I6287: std_logic; attribute dont_touch of I6287: signal is true;
	signal I6288: std_logic; attribute dont_touch of I6288: signal is true;
	signal I6289: std_logic; attribute dont_touch of I6289: signal is true;
	signal I6294: std_logic; attribute dont_touch of I6294: signal is true;
	signal I6299: std_logic; attribute dont_touch of I6299: signal is true;
	signal I6302: std_logic; attribute dont_touch of I6302: signal is true;
	signal I6309: std_logic; attribute dont_touch of I6309: signal is true;
	signal I6310: std_logic; attribute dont_touch of I6310: signal is true;
	signal I6316: std_logic; attribute dont_touch of I6316: signal is true;
	signal I6317: std_logic; attribute dont_touch of I6317: signal is true;
	signal I6322: std_logic; attribute dont_touch of I6322: signal is true;
	signal I6323: std_logic; attribute dont_touch of I6323: signal is true;
	signal I6324: std_logic; attribute dont_touch of I6324: signal is true;
	signal I6330: std_logic; attribute dont_touch of I6330: signal is true;
	signal I6331: std_logic; attribute dont_touch of I6331: signal is true;
	signal I6337: std_logic; attribute dont_touch of I6337: signal is true;
	signal I6338: std_logic; attribute dont_touch of I6338: signal is true;
	signal I6343: std_logic; attribute dont_touch of I6343: signal is true;
	signal I6347: std_logic; attribute dont_touch of I6347: signal is true;
	signal I6350: std_logic; attribute dont_touch of I6350: signal is true;
	signal I6351: std_logic; attribute dont_touch of I6351: signal is true;
	signal I6356: std_logic; attribute dont_touch of I6356: signal is true;
	signal I6360: std_logic; attribute dont_touch of I6360: signal is true;
	signal I6363: std_logic; attribute dont_touch of I6363: signal is true;
	signal I6367: std_logic; attribute dont_touch of I6367: signal is true;
	signal I6370: std_logic; attribute dont_touch of I6370: signal is true;
	signal I6373: std_logic; attribute dont_touch of I6373: signal is true;
	signal I6381: std_logic; attribute dont_touch of I6381: signal is true;
	signal I6385: std_logic; attribute dont_touch of I6385: signal is true;
	signal I6388: std_logic; attribute dont_touch of I6388: signal is true;
	signal I6391: std_logic; attribute dont_touch of I6391: signal is true;
	signal I6395: std_logic; attribute dont_touch of I6395: signal is true;
	signal I6398: std_logic; attribute dont_touch of I6398: signal is true;
	signal I6403: std_logic; attribute dont_touch of I6403: signal is true;
	signal I6406: std_logic; attribute dont_touch of I6406: signal is true;
	signal I6409: std_logic; attribute dont_touch of I6409: signal is true;
	signal I6414: std_logic; attribute dont_touch of I6414: signal is true;
	signal I6417: std_logic; attribute dont_touch of I6417: signal is true;
	signal I6421: std_logic; attribute dont_touch of I6421: signal is true;
	signal I6424: std_logic; attribute dont_touch of I6424: signal is true;
	signal I6428: std_logic; attribute dont_touch of I6428: signal is true;
	signal I6432: std_logic; attribute dont_touch of I6432: signal is true;
	signal I6436: std_logic; attribute dont_touch of I6436: signal is true;
	signal I6439: std_logic; attribute dont_touch of I6439: signal is true;
	signal I6443: std_logic; attribute dont_touch of I6443: signal is true;
	signal I6447: std_logic; attribute dont_touch of I6447: signal is true;
	signal I6448: std_logic; attribute dont_touch of I6448: signal is true;
	signal I6449: std_logic; attribute dont_touch of I6449: signal is true;
	signal I6454: std_logic; attribute dont_touch of I6454: signal is true;
	signal I6461: std_logic; attribute dont_touch of I6461: signal is true;
	signal I6467: std_logic; attribute dont_touch of I6467: signal is true;
	signal I6468: std_logic; attribute dont_touch of I6468: signal is true;
	signal I6469: std_logic; attribute dont_touch of I6469: signal is true;
	signal I6474: std_logic; attribute dont_touch of I6474: signal is true;
	signal I6477: std_logic; attribute dont_touch of I6477: signal is true;
	signal I6480: std_logic; attribute dont_touch of I6480: signal is true;
	signal I6484: std_logic; attribute dont_touch of I6484: signal is true;
	signal I6487: std_logic; attribute dont_touch of I6487: signal is true;
	signal I6488: std_logic; attribute dont_touch of I6488: signal is true;
	signal I6489: std_logic; attribute dont_touch of I6489: signal is true;
	signal I6495: std_logic; attribute dont_touch of I6495: signal is true;
	signal I6498: std_logic; attribute dont_touch of I6498: signal is true;
	signal I6501: std_logic; attribute dont_touch of I6501: signal is true;
	signal I6504: std_logic; attribute dont_touch of I6504: signal is true;
	signal I6507: std_logic; attribute dont_touch of I6507: signal is true;
	signal I6510: std_logic; attribute dont_touch of I6510: signal is true;
	signal I6513: std_logic; attribute dont_touch of I6513: signal is true;
	signal I6517: std_logic; attribute dont_touch of I6517: signal is true;
	signal I6520: std_logic; attribute dont_touch of I6520: signal is true;
	signal I6523: std_logic; attribute dont_touch of I6523: signal is true;
	signal I6528: std_logic; attribute dont_touch of I6528: signal is true;
	signal I6531: std_logic; attribute dont_touch of I6531: signal is true;
	signal I6535: std_logic; attribute dont_touch of I6535: signal is true;
	signal I6538: std_logic; attribute dont_touch of I6538: signal is true;
	signal I6543: std_logic; attribute dont_touch of I6543: signal is true;
	signal I6546: std_logic; attribute dont_touch of I6546: signal is true;
	signal I6549: std_logic; attribute dont_touch of I6549: signal is true;
	signal I6553: std_logic; attribute dont_touch of I6553: signal is true;
	signal I6557: std_logic; attribute dont_touch of I6557: signal is true;
	signal I6560: std_logic; attribute dont_touch of I6560: signal is true;
	signal I6565: std_logic; attribute dont_touch of I6565: signal is true;
	signal I6569: std_logic; attribute dont_touch of I6569: signal is true;
	signal I6572: std_logic; attribute dont_touch of I6572: signal is true;
	signal I6576: std_logic; attribute dont_touch of I6576: signal is true;
	signal I6580: std_logic; attribute dont_touch of I6580: signal is true;
	signal I6587: std_logic; attribute dont_touch of I6587: signal is true;
	signal I6590: std_logic; attribute dont_touch of I6590: signal is true;
	signal I6598: std_logic; attribute dont_touch of I6598: signal is true;
	signal I6601: std_logic; attribute dont_touch of I6601: signal is true;
	signal I6611: std_logic; attribute dont_touch of I6611: signal is true;
	signal I6616: std_logic; attribute dont_touch of I6616: signal is true;
	signal I6624: std_logic; attribute dont_touch of I6624: signal is true;
	signal I6630: std_logic; attribute dont_touch of I6630: signal is true;
	signal I6631: std_logic; attribute dont_touch of I6631: signal is true;
	signal I6639: std_logic; attribute dont_touch of I6639: signal is true;
	signal I6643: std_logic; attribute dont_touch of I6643: signal is true;
	signal I6648: std_logic; attribute dont_touch of I6648: signal is true;
	signal I6654: std_logic; attribute dont_touch of I6654: signal is true;
	signal I6661: std_logic; attribute dont_touch of I6661: signal is true;
	signal I6664: std_logic; attribute dont_touch of I6664: signal is true;
	signal I6665: std_logic; attribute dont_touch of I6665: signal is true;
	signal I6666: std_logic; attribute dont_touch of I6666: signal is true;
	signal I6671: std_logic; attribute dont_touch of I6671: signal is true;
	signal I6676: std_logic; attribute dont_touch of I6676: signal is true;
	signal I6679: std_logic; attribute dont_touch of I6679: signal is true;
	signal I6686: std_logic; attribute dont_touch of I6686: signal is true;
	signal I6690: std_logic; attribute dont_touch of I6690: signal is true;
	signal I6694: std_logic; attribute dont_touch of I6694: signal is true;
	signal I6702: std_logic; attribute dont_touch of I6702: signal is true;
	signal I6714: std_logic; attribute dont_touch of I6714: signal is true;
	signal I6715: std_logic; attribute dont_touch of I6715: signal is true;
	signal I6716: std_logic; attribute dont_touch of I6716: signal is true;
	signal I6726: std_logic; attribute dont_touch of I6726: signal is true;
	signal I6733: std_logic; attribute dont_touch of I6733: signal is true;
	signal I6738: std_logic; attribute dont_touch of I6738: signal is true;
	signal I6742: std_logic; attribute dont_touch of I6742: signal is true;
	signal I6746: std_logic; attribute dont_touch of I6746: signal is true;
	signal I6747: std_logic; attribute dont_touch of I6747: signal is true;
	signal I6748: std_logic; attribute dont_touch of I6748: signal is true;
	signal I6754: std_logic; attribute dont_touch of I6754: signal is true;
	signal I6757: std_logic; attribute dont_touch of I6757: signal is true;
	signal I6760: std_logic; attribute dont_touch of I6760: signal is true;
	signal I6761: std_logic; attribute dont_touch of I6761: signal is true;
	signal I6762: std_logic; attribute dont_touch of I6762: signal is true;
	signal I6767: std_logic; attribute dont_touch of I6767: signal is true;
	signal I6770: std_logic; attribute dont_touch of I6770: signal is true;
	signal I6771: std_logic; attribute dont_touch of I6771: signal is true;
	signal I6772: std_logic; attribute dont_touch of I6772: signal is true;
	signal I6777: std_logic; attribute dont_touch of I6777: signal is true;
	signal I6778: std_logic; attribute dont_touch of I6778: signal is true;
	signal I6779: std_logic; attribute dont_touch of I6779: signal is true;
	signal I6784: std_logic; attribute dont_touch of I6784: signal is true;
	signal I6789: std_logic; attribute dont_touch of I6789: signal is true;
	signal I6792: std_logic; attribute dont_touch of I6792: signal is true;
	signal I6793: std_logic; attribute dont_touch of I6793: signal is true;
	signal I6794: std_logic; attribute dont_touch of I6794: signal is true;
	signal I6799: std_logic; attribute dont_touch of I6799: signal is true;
	signal I6802: std_logic; attribute dont_touch of I6802: signal is true;
	signal I6805: std_logic; attribute dont_touch of I6805: signal is true;
	signal I6806: std_logic; attribute dont_touch of I6806: signal is true;
	signal I6807: std_logic; attribute dont_touch of I6807: signal is true;
	signal I6812: std_logic; attribute dont_touch of I6812: signal is true;
	signal I6815: std_logic; attribute dont_touch of I6815: signal is true;
	signal I6818: std_logic; attribute dont_touch of I6818: signal is true;
	signal I6821: std_logic; attribute dont_touch of I6821: signal is true;
	signal I6825: std_logic; attribute dont_touch of I6825: signal is true;
	signal I6826: std_logic; attribute dont_touch of I6826: signal is true;
	signal I6827: std_logic; attribute dont_touch of I6827: signal is true;
	signal I6832: std_logic; attribute dont_touch of I6832: signal is true;
	signal I6836: std_logic; attribute dont_touch of I6836: signal is true;
	signal I6837: std_logic; attribute dont_touch of I6837: signal is true;
	signal I6838: std_logic; attribute dont_touch of I6838: signal is true;
	signal I6844: std_logic; attribute dont_touch of I6844: signal is true;
	signal I6851: std_logic; attribute dont_touch of I6851: signal is true;
	signal I6856: std_logic; attribute dont_touch of I6856: signal is true;
	signal I6861: std_logic; attribute dont_touch of I6861: signal is true;
	signal I6867: std_logic; attribute dont_touch of I6867: signal is true;
	signal I6870: std_logic; attribute dont_touch of I6870: signal is true;
	signal I6876: std_logic; attribute dont_touch of I6876: signal is true;
	signal I6879: std_logic; attribute dont_touch of I6879: signal is true;
	signal I6880: std_logic; attribute dont_touch of I6880: signal is true;
	signal I6881: std_logic; attribute dont_touch of I6881: signal is true;
	signal I6888: std_logic; attribute dont_touch of I6888: signal is true;
	signal I6891: std_logic; attribute dont_touch of I6891: signal is true;
	signal I6894: std_logic; attribute dont_touch of I6894: signal is true;
	signal I6898: std_logic; attribute dont_touch of I6898: signal is true;
	signal I6901: std_logic; attribute dont_touch of I6901: signal is true;
	signal I6904: std_logic; attribute dont_touch of I6904: signal is true;
	signal I6907: std_logic; attribute dont_touch of I6907: signal is true;
	signal I6911: std_logic; attribute dont_touch of I6911: signal is true;
	signal I6914: std_logic; attribute dont_touch of I6914: signal is true;
	signal I6917: std_logic; attribute dont_touch of I6917: signal is true;
	signal I6921: std_logic; attribute dont_touch of I6921: signal is true;
	signal I6924: std_logic; attribute dont_touch of I6924: signal is true;
	signal I6929: std_logic; attribute dont_touch of I6929: signal is true;
	signal I6932: std_logic; attribute dont_touch of I6932: signal is true;
	signal I6938: std_logic; attribute dont_touch of I6938: signal is true;
	signal I6941: std_logic; attribute dont_touch of I6941: signal is true;
	signal I6944: std_logic; attribute dont_touch of I6944: signal is true;
	signal I6947: std_logic; attribute dont_touch of I6947: signal is true;
	signal I6952: std_logic; attribute dont_touch of I6952: signal is true;
	signal I6955: std_logic; attribute dont_touch of I6955: signal is true;
	signal I6958: std_logic; attribute dont_touch of I6958: signal is true;
	signal I6962: std_logic; attribute dont_touch of I6962: signal is true;
	signal I6965: std_logic; attribute dont_touch of I6965: signal is true;
	signal I6968: std_logic; attribute dont_touch of I6968: signal is true;
	signal I6971: std_logic; attribute dont_touch of I6971: signal is true;
	signal I6976: std_logic; attribute dont_touch of I6976: signal is true;
	signal I6979: std_logic; attribute dont_touch of I6979: signal is true;
	signal I6982: std_logic; attribute dont_touch of I6982: signal is true;
	signal I6985: std_logic; attribute dont_touch of I6985: signal is true;
	signal I6988: std_logic; attribute dont_touch of I6988: signal is true;
	signal I6989: std_logic; attribute dont_touch of I6989: signal is true;
	signal I6990: std_logic; attribute dont_touch of I6990: signal is true;
	signal I6996: std_logic; attribute dont_touch of I6996: signal is true;
	signal I6999: std_logic; attribute dont_touch of I6999: signal is true;
	signal I7002: std_logic; attribute dont_touch of I7002: signal is true;
	signal I7006: std_logic; attribute dont_touch of I7006: signal is true;
	signal I7009: std_logic; attribute dont_touch of I7009: signal is true;
	signal I7014: std_logic; attribute dont_touch of I7014: signal is true;
	signal I7017: std_logic; attribute dont_touch of I7017: signal is true;
	signal I7022: std_logic; attribute dont_touch of I7022: signal is true;
	signal I7029: std_logic; attribute dont_touch of I7029: signal is true;
	signal I7033: std_logic; attribute dont_touch of I7033: signal is true;
	signal I7034: std_logic; attribute dont_touch of I7034: signal is true;
	signal I7035: std_logic; attribute dont_touch of I7035: signal is true;
	signal I7043: std_logic; attribute dont_touch of I7043: signal is true;
	signal I7048: std_logic; attribute dont_touch of I7048: signal is true;
	signal I7054: std_logic; attribute dont_touch of I7054: signal is true;
	signal I7061: std_logic; attribute dont_touch of I7061: signal is true;
	signal I7064: std_logic; attribute dont_touch of I7064: signal is true;
	signal I7070: std_logic; attribute dont_touch of I7070: signal is true;
	signal I7076: std_logic; attribute dont_touch of I7076: signal is true;
	signal I7086: std_logic; attribute dont_touch of I7086: signal is true;
	signal I7096: std_logic; attribute dont_touch of I7096: signal is true;
	signal I7099: std_logic; attribute dont_touch of I7099: signal is true;
	signal I7104: std_logic; attribute dont_touch of I7104: signal is true;
	signal I7109: std_logic; attribute dont_touch of I7109: signal is true;
	signal I7112: std_logic; attribute dont_touch of I7112: signal is true;
	signal I7118: std_logic; attribute dont_touch of I7118: signal is true;
	signal I7131: std_logic; attribute dont_touch of I7131: signal is true;
	signal I7140: std_logic; attribute dont_touch of I7140: signal is true;
	signal I7143: std_logic; attribute dont_touch of I7143: signal is true;
	signal I7151: std_logic; attribute dont_touch of I7151: signal is true;
	signal I7154: std_logic; attribute dont_touch of I7154: signal is true;
	signal I7157: std_logic; attribute dont_touch of I7157: signal is true;
	signal I7163: std_logic; attribute dont_touch of I7163: signal is true;
	signal I7166: std_logic; attribute dont_touch of I7166: signal is true;
	signal I7173: std_logic; attribute dont_touch of I7173: signal is true;
	signal I7176: std_logic; attribute dont_touch of I7176: signal is true;
	signal I7182: std_logic; attribute dont_touch of I7182: signal is true;
	signal I7185: std_logic; attribute dont_touch of I7185: signal is true;
	signal I7191: std_logic; attribute dont_touch of I7191: signal is true;
	signal I7194: std_logic; attribute dont_touch of I7194: signal is true;
	signal I7202: std_logic; attribute dont_touch of I7202: signal is true;
	signal I7205: std_logic; attribute dont_touch of I7205: signal is true;
	signal I7210: std_logic; attribute dont_touch of I7210: signal is true;
	signal I7213: std_logic; attribute dont_touch of I7213: signal is true;
	signal I7216: std_logic; attribute dont_touch of I7216: signal is true;
	signal I7220: std_logic; attribute dont_touch of I7220: signal is true;
	signal I7223: std_logic; attribute dont_touch of I7223: signal is true;
	signal I7224: std_logic; attribute dont_touch of I7224: signal is true;
	signal I7225: std_logic; attribute dont_touch of I7225: signal is true;
	signal I7233: std_logic; attribute dont_touch of I7233: signal is true;
	signal I7236: std_logic; attribute dont_touch of I7236: signal is true;
	signal I7240: std_logic; attribute dont_touch of I7240: signal is true;
	signal I7244: std_logic; attribute dont_touch of I7244: signal is true;
	signal I7249: std_logic; attribute dont_touch of I7249: signal is true;
	signal I7255: std_logic; attribute dont_touch of I7255: signal is true;
	signal I7260: std_logic; attribute dont_touch of I7260: signal is true;
	signal I7264: std_logic; attribute dont_touch of I7264: signal is true;
	signal I7269: std_logic; attribute dont_touch of I7269: signal is true;
	signal I7272: std_logic; attribute dont_touch of I7272: signal is true;
	signal I7276: std_logic; attribute dont_touch of I7276: signal is true;
	signal I7280: std_logic; attribute dont_touch of I7280: signal is true;
	signal I7284: std_logic; attribute dont_touch of I7284: signal is true;
	signal I7288: std_logic; attribute dont_touch of I7288: signal is true;
	signal I7291: std_logic; attribute dont_touch of I7291: signal is true;
	signal I7295: std_logic; attribute dont_touch of I7295: signal is true;
	signal I7300: std_logic; attribute dont_touch of I7300: signal is true;
	signal I7303: std_logic; attribute dont_touch of I7303: signal is true;
	signal I7308: std_logic; attribute dont_touch of I7308: signal is true;
	signal I7311: std_logic; attribute dont_touch of I7311: signal is true;
	signal I7315: std_logic; attribute dont_touch of I7315: signal is true;
	signal I7318: std_logic; attribute dont_touch of I7318: signal is true;
	signal I7321: std_logic; attribute dont_touch of I7321: signal is true;
	signal I7322: std_logic; attribute dont_touch of I7322: signal is true;
	signal I7323: std_logic; attribute dont_touch of I7323: signal is true;
	signal I7330: std_logic; attribute dont_touch of I7330: signal is true;
	signal I7333: std_logic; attribute dont_touch of I7333: signal is true;
	signal I7336: std_logic; attribute dont_touch of I7336: signal is true;
	signal I7339: std_logic; attribute dont_touch of I7339: signal is true;
	signal I7342: std_logic; attribute dont_touch of I7342: signal is true;
	signal I7345: std_logic; attribute dont_touch of I7345: signal is true;
	signal I7348: std_logic; attribute dont_touch of I7348: signal is true;
	signal I7351: std_logic; attribute dont_touch of I7351: signal is true;
	signal I7354: std_logic; attribute dont_touch of I7354: signal is true;
	signal I7357: std_logic; attribute dont_touch of I7357: signal is true;
	signal I7360: std_logic; attribute dont_touch of I7360: signal is true;
	signal I7363: std_logic; attribute dont_touch of I7363: signal is true;
	signal I7366: std_logic; attribute dont_touch of I7366: signal is true;
	signal I7369: std_logic; attribute dont_touch of I7369: signal is true;
	signal I7372: std_logic; attribute dont_touch of I7372: signal is true;
	signal I7375: std_logic; attribute dont_touch of I7375: signal is true;
	signal I7378: std_logic; attribute dont_touch of I7378: signal is true;
	signal I7381: std_logic; attribute dont_touch of I7381: signal is true;
	signal I7384: std_logic; attribute dont_touch of I7384: signal is true;
	signal I7387: std_logic; attribute dont_touch of I7387: signal is true;
	signal I7390: std_logic; attribute dont_touch of I7390: signal is true;
	signal I7393: std_logic; attribute dont_touch of I7393: signal is true;
	signal I7396: std_logic; attribute dont_touch of I7396: signal is true;
	signal I7399: std_logic; attribute dont_touch of I7399: signal is true;
	signal I7402: std_logic; attribute dont_touch of I7402: signal is true;
	signal I7405: std_logic; attribute dont_touch of I7405: signal is true;
	signal I7408: std_logic; attribute dont_touch of I7408: signal is true;
	signal I7411: std_logic; attribute dont_touch of I7411: signal is true;
	signal I7414: std_logic; attribute dont_touch of I7414: signal is true;
	signal I7417: std_logic; attribute dont_touch of I7417: signal is true;
	signal I7420: std_logic; attribute dont_touch of I7420: signal is true;
	signal I7423: std_logic; attribute dont_touch of I7423: signal is true;
	signal I7426: std_logic; attribute dont_touch of I7426: signal is true;
	signal I7429: std_logic; attribute dont_touch of I7429: signal is true;
	signal I7432: std_logic; attribute dont_touch of I7432: signal is true;
	signal I7435: std_logic; attribute dont_touch of I7435: signal is true;
	signal I7438: std_logic; attribute dont_touch of I7438: signal is true;
	signal I7441: std_logic; attribute dont_touch of I7441: signal is true;
	signal I7444: std_logic; attribute dont_touch of I7444: signal is true;
	signal I7447: std_logic; attribute dont_touch of I7447: signal is true;
	signal I7450: std_logic; attribute dont_touch of I7450: signal is true;
	signal I7453: std_logic; attribute dont_touch of I7453: signal is true;
	signal I7456: std_logic; attribute dont_touch of I7456: signal is true;
	signal I7459: std_logic; attribute dont_touch of I7459: signal is true;
	signal I7462: std_logic; attribute dont_touch of I7462: signal is true;
	signal I7465: std_logic; attribute dont_touch of I7465: signal is true;
	signal I7468: std_logic; attribute dont_touch of I7468: signal is true;
	signal I7478: std_logic; attribute dont_touch of I7478: signal is true;
	signal I7487: std_logic; attribute dont_touch of I7487: signal is true;
	signal I7509: std_logic; attribute dont_touch of I7509: signal is true;
	signal I7513: std_logic; attribute dont_touch of I7513: signal is true;
	signal I7523: std_logic; attribute dont_touch of I7523: signal is true;
	signal I7536: std_logic; attribute dont_touch of I7536: signal is true;
	signal I7546: std_logic; attribute dont_touch of I7546: signal is true;
	signal I7556: std_logic; attribute dont_touch of I7556: signal is true;
	signal I7559: std_logic; attribute dont_touch of I7559: signal is true;
	signal I7562: std_logic; attribute dont_touch of I7562: signal is true;
	signal I7563: std_logic; attribute dont_touch of I7563: signal is true;
	signal I7564: std_logic; attribute dont_touch of I7564: signal is true;
	signal I7577: std_logic; attribute dont_touch of I7577: signal is true;
	signal I7586: std_logic; attribute dont_touch of I7586: signal is true;
	signal I7593: std_logic; attribute dont_touch of I7593: signal is true;
	signal I7600: std_logic; attribute dont_touch of I7600: signal is true;
	signal I7606: std_logic; attribute dont_touch of I7606: signal is true;
	signal I7612: std_logic; attribute dont_touch of I7612: signal is true;
	signal I7625: std_logic; attribute dont_touch of I7625: signal is true;
	signal I7630: std_logic; attribute dont_touch of I7630: signal is true;
	signal I7633: std_logic; attribute dont_touch of I7633: signal is true;
	signal I7636: std_logic; attribute dont_touch of I7636: signal is true;
	signal I7639: std_logic; attribute dont_touch of I7639: signal is true;
	signal I7642: std_logic; attribute dont_touch of I7642: signal is true;
	signal I7648: std_logic; attribute dont_touch of I7648: signal is true;
	signal I7651: std_logic; attribute dont_touch of I7651: signal is true;
	signal I7654: std_logic; attribute dont_touch of I7654: signal is true;
	signal I7659: std_logic; attribute dont_touch of I7659: signal is true;
	signal I7662: std_logic; attribute dont_touch of I7662: signal is true;
	signal I7665: std_logic; attribute dont_touch of I7665: signal is true;
	signal I7668: std_logic; attribute dont_touch of I7668: signal is true;
	signal I7671: std_logic; attribute dont_touch of I7671: signal is true;
	signal I7674: std_logic; attribute dont_touch of I7674: signal is true;
	signal I7677: std_logic; attribute dont_touch of I7677: signal is true;
	signal I7680: std_logic; attribute dont_touch of I7680: signal is true;
	signal I7683: std_logic; attribute dont_touch of I7683: signal is true;
	signal I7684: std_logic; attribute dont_touch of I7684: signal is true;
	signal I7685: std_logic; attribute dont_touch of I7685: signal is true;
	signal I7691: std_logic; attribute dont_touch of I7691: signal is true;
	signal I7694: std_logic; attribute dont_touch of I7694: signal is true;
	signal I7697: std_logic; attribute dont_touch of I7697: signal is true;
	signal I7701: std_logic; attribute dont_touch of I7701: signal is true;
	signal I7707: std_logic; attribute dont_touch of I7707: signal is true;
	signal I7710: std_logic; attribute dont_touch of I7710: signal is true;
	signal I7713: std_logic; attribute dont_touch of I7713: signal is true;
	signal I7716: std_logic; attribute dont_touch of I7716: signal is true;
	signal I7719: std_logic; attribute dont_touch of I7719: signal is true;
	signal I7726: std_logic; attribute dont_touch of I7726: signal is true;
	signal I7729: std_logic; attribute dont_touch of I7729: signal is true;
	signal I7732: std_logic; attribute dont_touch of I7732: signal is true;
	signal I7735: std_logic; attribute dont_touch of I7735: signal is true;
	signal I7743: std_logic; attribute dont_touch of I7743: signal is true;
	signal I7746: std_logic; attribute dont_touch of I7746: signal is true;
	signal I7749: std_logic; attribute dont_touch of I7749: signal is true;
	signal I7752: std_logic; attribute dont_touch of I7752: signal is true;
	signal I7757: std_logic; attribute dont_touch of I7757: signal is true;
	signal I7760: std_logic; attribute dont_touch of I7760: signal is true;
	signal I7763: std_logic; attribute dont_touch of I7763: signal is true;
	signal I7766: std_logic; attribute dont_touch of I7766: signal is true;
	signal I7771: std_logic; attribute dont_touch of I7771: signal is true;
	signal I7776: std_logic; attribute dont_touch of I7776: signal is true;
	signal I7779: std_logic; attribute dont_touch of I7779: signal is true;
	signal I7782: std_logic; attribute dont_touch of I7782: signal is true;
	signal I7790: std_logic; attribute dont_touch of I7790: signal is true;
	signal I7793: std_logic; attribute dont_touch of I7793: signal is true;
	signal I7800: std_logic; attribute dont_touch of I7800: signal is true;
	signal I7803: std_logic; attribute dont_touch of I7803: signal is true;
	signal I7810: std_logic; attribute dont_touch of I7810: signal is true;
	signal I7817: std_logic; attribute dont_touch of I7817: signal is true;
	signal I7820: std_logic; attribute dont_touch of I7820: signal is true;
	signal I7825: std_logic; attribute dont_touch of I7825: signal is true;
	signal I7829: std_logic; attribute dont_touch of I7829: signal is true;
	signal I7833: std_logic; attribute dont_touch of I7833: signal is true;
	signal I7837: std_logic; attribute dont_touch of I7837: signal is true;
	signal I7840: std_logic; attribute dont_touch of I7840: signal is true;
	signal I7843: std_logic; attribute dont_touch of I7843: signal is true;
	signal I7847: std_logic; attribute dont_touch of I7847: signal is true;
	signal I7852: std_logic; attribute dont_touch of I7852: signal is true;
	signal I7858: std_logic; attribute dont_touch of I7858: signal is true;
	signal I7863: std_logic; attribute dont_touch of I7863: signal is true;
	signal I7864: std_logic; attribute dont_touch of I7864: signal is true;
	signal I7865: std_logic; attribute dont_touch of I7865: signal is true;
	signal I7875: std_logic; attribute dont_touch of I7875: signal is true;
	signal I7876: std_logic; attribute dont_touch of I7876: signal is true;
	signal I7877: std_logic; attribute dont_touch of I7877: signal is true;
	signal I7886: std_logic; attribute dont_touch of I7886: signal is true;
	signal I7889: std_logic; attribute dont_touch of I7889: signal is true;
	signal I7899: std_logic; attribute dont_touch of I7899: signal is true;
	signal I7906: std_logic; attribute dont_touch of I7906: signal is true;
	signal I7909: std_logic; attribute dont_touch of I7909: signal is true;
	signal I7916: std_logic; attribute dont_touch of I7916: signal is true;
	signal I7920: std_logic; attribute dont_touch of I7920: signal is true;
	signal I7923: std_logic; attribute dont_touch of I7923: signal is true;
	signal I7931: std_logic; attribute dont_touch of I7931: signal is true;
	signal I7935: std_logic; attribute dont_touch of I7935: signal is true;
	signal I7938: std_logic; attribute dont_touch of I7938: signal is true;
	signal I7946: std_logic; attribute dont_touch of I7946: signal is true;
	signal I7952: std_logic; attribute dont_touch of I7952: signal is true;
	signal I7956: std_logic; attribute dont_touch of I7956: signal is true;
	signal I7964: std_logic; attribute dont_touch of I7964: signal is true;
	signal I7973: std_logic; attribute dont_touch of I7973: signal is true;
	signal I7984: std_logic; attribute dont_touch of I7984: signal is true;
	signal I7996: std_logic; attribute dont_touch of I7996: signal is true;
	signal I7999: std_logic; attribute dont_touch of I7999: signal is true;
	signal I8004: std_logic; attribute dont_touch of I8004: signal is true;
	signal I8007: std_logic; attribute dont_touch of I8007: signal is true;
	signal I8011: std_logic; attribute dont_touch of I8011: signal is true;
	signal I8024: std_logic; attribute dont_touch of I8024: signal is true;
	signal I8031: std_logic; attribute dont_touch of I8031: signal is true;
	signal I8036: std_logic; attribute dont_touch of I8036: signal is true;
	signal I8039: std_logic; attribute dont_touch of I8039: signal is true;
	signal I8050: std_logic; attribute dont_touch of I8050: signal is true;
	signal I8061: std_logic; attribute dont_touch of I8061: signal is true;
	signal I8080: std_logic; attribute dont_touch of I8080: signal is true;
	signal I8085: std_logic; attribute dont_touch of I8085: signal is true;
	signal I8089: std_logic; attribute dont_touch of I8089: signal is true;
	signal I8098: std_logic; attribute dont_touch of I8098: signal is true;
	signal I8109: std_logic; attribute dont_touch of I8109: signal is true;
	signal I8116: std_logic; attribute dont_touch of I8116: signal is true;
	signal I8123: std_logic; attribute dont_touch of I8123: signal is true;
	signal I8126: std_logic; attribute dont_touch of I8126: signal is true;
	signal I8133: std_logic; attribute dont_touch of I8133: signal is true;
	signal I8136: std_logic; attribute dont_touch of I8136: signal is true;
	signal I8139: std_logic; attribute dont_touch of I8139: signal is true;
	signal I8147: std_logic; attribute dont_touch of I8147: signal is true;
	signal I8154: std_logic; attribute dont_touch of I8154: signal is true;
	signal I8161: std_logic; attribute dont_touch of I8161: signal is true;
	signal I8164: std_logic; attribute dont_touch of I8164: signal is true;
	signal I8178: std_logic; attribute dont_touch of I8178: signal is true;
	signal I8179: std_logic; attribute dont_touch of I8179: signal is true;
	signal I8180: std_logic; attribute dont_touch of I8180: signal is true;
	signal I8192: std_logic; attribute dont_touch of I8192: signal is true;
	signal I8199: std_logic; attribute dont_touch of I8199: signal is true;
	signal I8204: std_logic; attribute dont_touch of I8204: signal is true;
	signal I8211: std_logic; attribute dont_touch of I8211: signal is true;
	signal I8215: std_logic; attribute dont_touch of I8215: signal is true;
	signal I8228: std_logic; attribute dont_touch of I8228: signal is true;
	signal I8231: std_logic; attribute dont_touch of I8231: signal is true;
	signal I8234: std_logic; attribute dont_touch of I8234: signal is true;
	signal I8237: std_logic; attribute dont_touch of I8237: signal is true;
	signal I8240: std_logic; attribute dont_touch of I8240: signal is true;
	signal I8247: std_logic; attribute dont_touch of I8247: signal is true;
	signal I8250: std_logic; attribute dont_touch of I8250: signal is true;
	signal I8253: std_logic; attribute dont_touch of I8253: signal is true;
	signal I8256: std_logic; attribute dont_touch of I8256: signal is true;
	signal I8259: std_logic; attribute dont_touch of I8259: signal is true;
	signal I8262: std_logic; attribute dont_touch of I8262: signal is true;
	signal I8265: std_logic; attribute dont_touch of I8265: signal is true;
	signal I8268: std_logic; attribute dont_touch of I8268: signal is true;
	signal I8275: std_logic; attribute dont_touch of I8275: signal is true;
	signal I8278: std_logic; attribute dont_touch of I8278: signal is true;
	signal I8282: std_logic; attribute dont_touch of I8282: signal is true;
	signal I8285: std_logic; attribute dont_touch of I8285: signal is true;
	signal I8290: std_logic; attribute dont_touch of I8290: signal is true;
	signal I8293: std_logic; attribute dont_touch of I8293: signal is true;
	signal I8298: std_logic; attribute dont_touch of I8298: signal is true;
	signal I8303: std_logic; attribute dont_touch of I8303: signal is true;
	signal I8308: std_logic; attribute dont_touch of I8308: signal is true;
	signal I8311: std_logic; attribute dont_touch of I8311: signal is true;
	signal I8315: std_logic; attribute dont_touch of I8315: signal is true;
	signal I8320: std_logic; attribute dont_touch of I8320: signal is true;
	signal I8324: std_logic; attribute dont_touch of I8324: signal is true;
	signal I8328: std_logic; attribute dont_touch of I8328: signal is true;
	signal I8333: std_logic; attribute dont_touch of I8333: signal is true;
	signal I8337: std_logic; attribute dont_touch of I8337: signal is true;
	signal I8340: std_logic; attribute dont_touch of I8340: signal is true;
	signal I8351: std_logic; attribute dont_touch of I8351: signal is true;
	signal I8358: std_logic; attribute dont_touch of I8358: signal is true;
	signal I8379: std_logic; attribute dont_touch of I8379: signal is true;
	signal I8385: std_logic; attribute dont_touch of I8385: signal is true;
	signal I8388: std_logic; attribute dont_touch of I8388: signal is true;
	signal I8396: std_logic; attribute dont_touch of I8396: signal is true;
	signal I8403: std_logic; attribute dont_touch of I8403: signal is true;
	signal I8406: std_logic; attribute dont_touch of I8406: signal is true;
	signal I8410: std_logic; attribute dont_touch of I8410: signal is true;
	signal I8414: std_logic; attribute dont_touch of I8414: signal is true;
	signal I8418: std_logic; attribute dont_touch of I8418: signal is true;
	signal I8421: std_logic; attribute dont_touch of I8421: signal is true;
	signal I8429: std_logic; attribute dont_touch of I8429: signal is true;
	signal I8436: std_logic; attribute dont_touch of I8436: signal is true;
	signal I8442: std_logic; attribute dont_touch of I8442: signal is true;
	signal I8449: std_logic; attribute dont_touch of I8449: signal is true;
	signal I8456: std_logic; attribute dont_touch of I8456: signal is true;
	signal I8462: std_logic; attribute dont_touch of I8462: signal is true;
	signal I8465: std_logic; attribute dont_touch of I8465: signal is true;
	signal I8473: std_logic; attribute dont_touch of I8473: signal is true;
	signal I8476: std_logic; attribute dont_touch of I8476: signal is true;
	signal I8479: std_logic; attribute dont_touch of I8479: signal is true;
	signal I8480: std_logic; attribute dont_touch of I8480: signal is true;
	signal I8481: std_logic; attribute dont_touch of I8481: signal is true;
	signal I8487: std_logic; attribute dont_touch of I8487: signal is true;
	signal I8490: std_logic; attribute dont_touch of I8490: signal is true;
	signal I8495: std_logic; attribute dont_touch of I8495: signal is true;
	signal I8499: std_logic; attribute dont_touch of I8499: signal is true;
	signal I8503: std_logic; attribute dont_touch of I8503: signal is true;
	signal I8506: std_logic; attribute dont_touch of I8506: signal is true;
	signal I8513: std_logic; attribute dont_touch of I8513: signal is true;
	signal I8514: std_logic; attribute dont_touch of I8514: signal is true;
	signal I8515: std_logic; attribute dont_touch of I8515: signal is true;
	signal I8520: std_logic; attribute dont_touch of I8520: signal is true;
	signal I8527: std_logic; attribute dont_touch of I8527: signal is true;
	signal I8528: std_logic; attribute dont_touch of I8528: signal is true;
	signal I8529: std_logic; attribute dont_touch of I8529: signal is true;
	signal I8535: std_logic; attribute dont_touch of I8535: signal is true;
	signal I8543: std_logic; attribute dont_touch of I8543: signal is true;
	signal I8544: std_logic; attribute dont_touch of I8544: signal is true;
	signal I8545: std_logic; attribute dont_touch of I8545: signal is true;
	signal I8551: std_logic; attribute dont_touch of I8551: signal is true;
	signal I8561: std_logic; attribute dont_touch of I8561: signal is true;
	signal I8562: std_logic; attribute dont_touch of I8562: signal is true;
	signal I8563: std_logic; attribute dont_touch of I8563: signal is true;
	signal I8575: std_logic; attribute dont_touch of I8575: signal is true;
	signal I8576: std_logic; attribute dont_touch of I8576: signal is true;
	signal I8577: std_logic; attribute dont_touch of I8577: signal is true;
	signal I8589: std_logic; attribute dont_touch of I8589: signal is true;
	signal I8590: std_logic; attribute dont_touch of I8590: signal is true;
	signal I8591: std_logic; attribute dont_touch of I8591: signal is true;
	signal I8604: std_logic; attribute dont_touch of I8604: signal is true;
	signal I8605: std_logic; attribute dont_touch of I8605: signal is true;
	signal I8606: std_logic; attribute dont_touch of I8606: signal is true;
	signal I8611: std_logic; attribute dont_touch of I8611: signal is true;
	signal I8614: std_logic; attribute dont_touch of I8614: signal is true;
	signal I8624: std_logic; attribute dont_touch of I8624: signal is true;
	signal I8625: std_logic; attribute dont_touch of I8625: signal is true;
	signal I8626: std_logic; attribute dont_touch of I8626: signal is true;
	signal I8631: std_logic; attribute dont_touch of I8631: signal is true;
	signal I8640: std_logic; attribute dont_touch of I8640: signal is true;
	signal I8641: std_logic; attribute dont_touch of I8641: signal is true;
	signal I8642: std_logic; attribute dont_touch of I8642: signal is true;
	signal I8647: std_logic; attribute dont_touch of I8647: signal is true;
	signal I8650: std_logic; attribute dont_touch of I8650: signal is true;
	signal I8651: std_logic; attribute dont_touch of I8651: signal is true;
	signal I8652: std_logic; attribute dont_touch of I8652: signal is true;
	signal I8662: std_logic; attribute dont_touch of I8662: signal is true;
	signal I8663: std_logic; attribute dont_touch of I8663: signal is true;
	signal I8664: std_logic; attribute dont_touch of I8664: signal is true;
	signal I8669: std_logic; attribute dont_touch of I8669: signal is true;
	signal I8670: std_logic; attribute dont_touch of I8670: signal is true;
	signal I8671: std_logic; attribute dont_touch of I8671: signal is true;
	signal I8676: std_logic; attribute dont_touch of I8676: signal is true;
	signal I8677: std_logic; attribute dont_touch of I8677: signal is true;
	signal I8678: std_logic; attribute dont_touch of I8678: signal is true;
	signal I8711: std_logic; attribute dont_touch of I8711: signal is true;
	signal I8715: std_logic; attribute dont_touch of I8715: signal is true;
	signal I8716: std_logic; attribute dont_touch of I8716: signal is true;
	signal I8717: std_logic; attribute dont_touch of I8717: signal is true;
	signal I8724: std_logic; attribute dont_touch of I8724: signal is true;
	signal I8728: std_logic; attribute dont_touch of I8728: signal is true;
	signal I8729: std_logic; attribute dont_touch of I8729: signal is true;
	signal I8730: std_logic; attribute dont_touch of I8730: signal is true;
	signal I8738: std_logic; attribute dont_touch of I8738: signal is true;
	signal I8739: std_logic; attribute dont_touch of I8739: signal is true;
	signal I8740: std_logic; attribute dont_touch of I8740: signal is true;
	signal I8750: std_logic; attribute dont_touch of I8750: signal is true;
	signal I8751: std_logic; attribute dont_touch of I8751: signal is true;
	signal I8752: std_logic; attribute dont_touch of I8752: signal is true;
	signal I8761: std_logic; attribute dont_touch of I8761: signal is true;
	signal I8762: std_logic; attribute dont_touch of I8762: signal is true;
	signal I8763: std_logic; attribute dont_touch of I8763: signal is true;
	signal I8770: std_logic; attribute dont_touch of I8770: signal is true;
	signal I8771: std_logic; attribute dont_touch of I8771: signal is true;
	signal I8772: std_logic; attribute dont_touch of I8772: signal is true;
	signal I8778: std_logic; attribute dont_touch of I8778: signal is true;
	signal I8779: std_logic; attribute dont_touch of I8779: signal is true;
	signal I8780: std_logic; attribute dont_touch of I8780: signal is true;
	signal I8786: std_logic; attribute dont_touch of I8786: signal is true;
	signal I8787: std_logic; attribute dont_touch of I8787: signal is true;
	signal I8788: std_logic; attribute dont_touch of I8788: signal is true;
	signal I8795: std_logic; attribute dont_touch of I8795: signal is true;
	signal I8796: std_logic; attribute dont_touch of I8796: signal is true;
	signal I8797: std_logic; attribute dont_touch of I8797: signal is true;
	signal I8803: std_logic; attribute dont_touch of I8803: signal is true;
	signal I8804: std_logic; attribute dont_touch of I8804: signal is true;
	signal I8805: std_logic; attribute dont_touch of I8805: signal is true;
	signal I8811: std_logic; attribute dont_touch of I8811: signal is true;
	signal I8815: std_logic; attribute dont_touch of I8815: signal is true;
	signal I8820: std_logic; attribute dont_touch of I8820: signal is true;
	signal I8827: std_logic; attribute dont_touch of I8827: signal is true;
	signal I8831: std_logic; attribute dont_touch of I8831: signal is true;
	signal I8835: std_logic; attribute dont_touch of I8835: signal is true;
	signal I8839: std_logic; attribute dont_touch of I8839: signal is true;
	signal I8842: std_logic; attribute dont_touch of I8842: signal is true;
	signal I8848: std_logic; attribute dont_touch of I8848: signal is true;
	signal I8851: std_logic; attribute dont_touch of I8851: signal is true;
	signal I8854: std_logic; attribute dont_touch of I8854: signal is true;
	signal I8858: std_logic; attribute dont_touch of I8858: signal is true;
	signal I8865: std_logic; attribute dont_touch of I8865: signal is true;
	signal I8869: std_logic; attribute dont_touch of I8869: signal is true;
	signal I8872: std_logic; attribute dont_touch of I8872: signal is true;
	signal I8877: std_logic; attribute dont_touch of I8877: signal is true;
	signal I8880: std_logic; attribute dont_touch of I8880: signal is true;
	signal I8885: std_logic; attribute dont_touch of I8885: signal is true;
	signal I8889: std_logic; attribute dont_touch of I8889: signal is true;
	signal I8892: std_logic; attribute dont_touch of I8892: signal is true;
	signal I8900: std_logic; attribute dont_touch of I8900: signal is true;
	signal I8903: std_logic; attribute dont_touch of I8903: signal is true;
	signal I8911: std_logic; attribute dont_touch of I8911: signal is true;
	signal I8919: std_logic; attribute dont_touch of I8919: signal is true;
	signal I8929: std_logic; attribute dont_touch of I8929: signal is true;
	signal I8934: std_logic; attribute dont_touch of I8934: signal is true;
	signal I8943: std_logic; attribute dont_touch of I8943: signal is true;
	signal I8967: std_logic; attribute dont_touch of I8967: signal is true;
	signal I8973: std_logic; attribute dont_touch of I8973: signal is true;
	signal I8982: std_logic; attribute dont_touch of I8982: signal is true;
	signal I8985: std_logic; attribute dont_touch of I8985: signal is true;
	signal I8989: std_logic; attribute dont_touch of I8989: signal is true;
	signal I8996: std_logic; attribute dont_touch of I8996: signal is true;
	signal I9001: std_logic; attribute dont_touch of I9001: signal is true;
	signal I9006: std_logic; attribute dont_touch of I9006: signal is true;
	signal I9007: std_logic; attribute dont_touch of I9007: signal is true;
	signal I9008: std_logic; attribute dont_touch of I9008: signal is true;
	signal I9013: std_logic; attribute dont_touch of I9013: signal is true;
	signal I9016: std_logic; attribute dont_touch of I9016: signal is true;
	signal I9020: std_logic; attribute dont_touch of I9020: signal is true;
	signal I9023: std_logic; attribute dont_touch of I9023: signal is true;
	signal I9029: std_logic; attribute dont_touch of I9029: signal is true;
	signal I9032: std_logic; attribute dont_touch of I9032: signal is true;
	signal I9040: std_logic; attribute dont_touch of I9040: signal is true;
	signal I9043: std_logic; attribute dont_touch of I9043: signal is true;
	signal I9046: std_logic; attribute dont_touch of I9046: signal is true;
	signal I9053: std_logic; attribute dont_touch of I9053: signal is true;
	signal I9056: std_logic; attribute dont_touch of I9056: signal is true;
	signal I9062: std_logic; attribute dont_touch of I9062: signal is true;
	signal I9065: std_logic; attribute dont_touch of I9065: signal is true;
	signal I9068: std_logic; attribute dont_touch of I9068: signal is true;
	signal I9074: std_logic; attribute dont_touch of I9074: signal is true;
	signal I9077: std_logic; attribute dont_touch of I9077: signal is true;
	signal I9080: std_logic; attribute dont_touch of I9080: signal is true;
	signal I9084: std_logic; attribute dont_touch of I9084: signal is true;
	signal I9087: std_logic; attribute dont_touch of I9087: signal is true;
	signal I9090: std_logic; attribute dont_touch of I9090: signal is true;
	signal I9093: std_logic; attribute dont_touch of I9093: signal is true;
	signal I9096: std_logic; attribute dont_touch of I9096: signal is true;
	signal I9099: std_logic; attribute dont_touch of I9099: signal is true;
	signal I9102: std_logic; attribute dont_touch of I9102: signal is true;
	signal I9105: std_logic; attribute dont_touch of I9105: signal is true;
	signal I9108: std_logic; attribute dont_touch of I9108: signal is true;
	signal I9111: std_logic; attribute dont_touch of I9111: signal is true;
	signal I9114: std_logic; attribute dont_touch of I9114: signal is true;
	signal I9117: std_logic; attribute dont_touch of I9117: signal is true;
	signal I9120: std_logic; attribute dont_touch of I9120: signal is true;
	signal I9123: std_logic; attribute dont_touch of I9123: signal is true;
	signal I9126: std_logic; attribute dont_touch of I9126: signal is true;
	signal I9129: std_logic; attribute dont_touch of I9129: signal is true;
	signal I9132: std_logic; attribute dont_touch of I9132: signal is true;
	signal I9135: std_logic; attribute dont_touch of I9135: signal is true;
	signal I9138: std_logic; attribute dont_touch of I9138: signal is true;
	signal I9141: std_logic; attribute dont_touch of I9141: signal is true;
	signal I9144: std_logic; attribute dont_touch of I9144: signal is true;
	signal I9147: std_logic; attribute dont_touch of I9147: signal is true;
	signal I9150: std_logic; attribute dont_touch of I9150: signal is true;
	signal I9153: std_logic; attribute dont_touch of I9153: signal is true;
	signal I9156: std_logic; attribute dont_touch of I9156: signal is true;
	signal I9159: std_logic; attribute dont_touch of I9159: signal is true;
	signal I9162: std_logic; attribute dont_touch of I9162: signal is true;
	signal I9165: std_logic; attribute dont_touch of I9165: signal is true;
	signal I9168: std_logic; attribute dont_touch of I9168: signal is true;
	signal I9171: std_logic; attribute dont_touch of I9171: signal is true;
	signal I9174: std_logic; attribute dont_touch of I9174: signal is true;
	signal I9177: std_logic; attribute dont_touch of I9177: signal is true;
	signal I9180: std_logic; attribute dont_touch of I9180: signal is true;
	signal I9185: std_logic; attribute dont_touch of I9185: signal is true;
	signal I9188: std_logic; attribute dont_touch of I9188: signal is true;
	signal I9191: std_logic; attribute dont_touch of I9191: signal is true;
	signal I9194: std_logic; attribute dont_touch of I9194: signal is true;
	signal I9199: std_logic; attribute dont_touch of I9199: signal is true;
	signal I9202: std_logic; attribute dont_touch of I9202: signal is true;
	signal I9205: std_logic; attribute dont_touch of I9205: signal is true;
	signal I9208: std_logic; attribute dont_touch of I9208: signal is true;
	signal I9213: std_logic; attribute dont_touch of I9213: signal is true;
	signal I9216: std_logic; attribute dont_touch of I9216: signal is true;
	signal I9221: std_logic; attribute dont_touch of I9221: signal is true;
	signal I9224: std_logic; attribute dont_touch of I9224: signal is true;
	signal I9229: std_logic; attribute dont_touch of I9229: signal is true;
	signal I9232: std_logic; attribute dont_touch of I9232: signal is true;
	signal I9237: std_logic; attribute dont_touch of I9237: signal is true;
	signal I9240: std_logic; attribute dont_touch of I9240: signal is true;
	signal I9243: std_logic; attribute dont_touch of I9243: signal is true;
	signal I9248: std_logic; attribute dont_touch of I9248: signal is true;
	signal I9253: std_logic; attribute dont_touch of I9253: signal is true;
	signal I9256: std_logic; attribute dont_touch of I9256: signal is true;
	signal I9259: std_logic; attribute dont_touch of I9259: signal is true;
	signal I9265: std_logic; attribute dont_touch of I9265: signal is true;
	signal I9268: std_logic; attribute dont_touch of I9268: signal is true;
	signal I9273: std_logic; attribute dont_touch of I9273: signal is true;
	signal I9276: std_logic; attribute dont_touch of I9276: signal is true;
	signal I9279: std_logic; attribute dont_touch of I9279: signal is true;
	signal I9282: std_logic; attribute dont_touch of I9282: signal is true;
	signal I9287: std_logic; attribute dont_touch of I9287: signal is true;
	signal I9290: std_logic; attribute dont_touch of I9290: signal is true;
	signal I9293: std_logic; attribute dont_touch of I9293: signal is true;
	signal I9296: std_logic; attribute dont_touch of I9296: signal is true;
	signal I9302: std_logic; attribute dont_touch of I9302: signal is true;
	signal I9305: std_logic; attribute dont_touch of I9305: signal is true;
	signal I9308: std_logic; attribute dont_touch of I9308: signal is true;
	signal I9311: std_logic; attribute dont_touch of I9311: signal is true;
	signal I9317: std_logic; attribute dont_touch of I9317: signal is true;
	signal I9320: std_logic; attribute dont_touch of I9320: signal is true;
	signal I9323: std_logic; attribute dont_touch of I9323: signal is true;
	signal I9326: std_logic; attribute dont_touch of I9326: signal is true;
	signal I9329: std_logic; attribute dont_touch of I9329: signal is true;
	signal I9332: std_logic; attribute dont_touch of I9332: signal is true;
	signal I9338: std_logic; attribute dont_touch of I9338: signal is true;
	signal I9341: std_logic; attribute dont_touch of I9341: signal is true;
	signal I9346: std_logic; attribute dont_touch of I9346: signal is true;
	signal I9349: std_logic; attribute dont_touch of I9349: signal is true;
	signal I9352: std_logic; attribute dont_touch of I9352: signal is true;
	signal I9359: std_logic; attribute dont_touch of I9359: signal is true;
	signal I9362: std_logic; attribute dont_touch of I9362: signal is true;
	signal I9365: std_logic; attribute dont_touch of I9365: signal is true;
	signal I9368: std_logic; attribute dont_touch of I9368: signal is true;
	signal I9371: std_logic; attribute dont_touch of I9371: signal is true;
	signal I9377: std_logic; attribute dont_touch of I9377: signal is true;
	signal I9380: std_logic; attribute dont_touch of I9380: signal is true;
	signal I9383: std_logic; attribute dont_touch of I9383: signal is true;
	signal I9388: std_logic; attribute dont_touch of I9388: signal is true;
	signal I9391: std_logic; attribute dont_touch of I9391: signal is true;
	signal I9394: std_logic; attribute dont_touch of I9394: signal is true;
	signal I9399: std_logic; attribute dont_touch of I9399: signal is true;
	signal I9402: std_logic; attribute dont_touch of I9402: signal is true;
	signal I9409: std_logic; attribute dont_touch of I9409: signal is true;
	signal I9415: std_logic; attribute dont_touch of I9415: signal is true;
	signal I9421: std_logic; attribute dont_touch of I9421: signal is true;
	signal I9424: std_logic; attribute dont_touch of I9424: signal is true;
	signal I9427: std_logic; attribute dont_touch of I9427: signal is true;
	signal I9433: std_logic; attribute dont_touch of I9433: signal is true;
	signal I9440: std_logic; attribute dont_touch of I9440: signal is true;
	signal I9443: std_logic; attribute dont_touch of I9443: signal is true;
	signal I9446: std_logic; attribute dont_touch of I9446: signal is true;
	signal I9452: std_logic; attribute dont_touch of I9452: signal is true;
	signal I9458: std_logic; attribute dont_touch of I9458: signal is true;
	signal I9461: std_logic; attribute dont_touch of I9461: signal is true;
	signal I9475: std_logic; attribute dont_touch of I9475: signal is true;
	signal I9479: std_logic; attribute dont_touch of I9479: signal is true;
	signal I9483: std_logic; attribute dont_touch of I9483: signal is true;
	signal I9486: std_logic; attribute dont_touch of I9486: signal is true;
	signal I9491: std_logic; attribute dont_touch of I9491: signal is true;
	signal I9498: std_logic; attribute dont_touch of I9498: signal is true;
	signal I9505: std_logic; attribute dont_touch of I9505: signal is true;
	signal I9510: std_logic; attribute dont_touch of I9510: signal is true;
	signal I9514: std_logic; attribute dont_touch of I9514: signal is true;
	signal I9519: std_logic; attribute dont_touch of I9519: signal is true;
	signal I9525: std_logic; attribute dont_touch of I9525: signal is true;
	signal I9531: std_logic; attribute dont_touch of I9531: signal is true;
	signal I9536: std_logic; attribute dont_touch of I9536: signal is true;
	signal I9539: std_logic; attribute dont_touch of I9539: signal is true;
	signal I9544: std_logic; attribute dont_touch of I9544: signal is true;
	signal I9550: std_logic; attribute dont_touch of I9550: signal is true;
	signal I9557: std_logic; attribute dont_touch of I9557: signal is true;
	signal I9558: std_logic; attribute dont_touch of I9558: signal is true;
	signal I9559: std_logic; attribute dont_touch of I9559: signal is true;
	signal I9564: std_logic; attribute dont_touch of I9564: signal is true;
	signal I9567: std_logic; attribute dont_touch of I9567: signal is true;
	signal I9571: std_logic; attribute dont_touch of I9571: signal is true;
	signal I9574: std_logic; attribute dont_touch of I9574: signal is true;
	signal I9575: std_logic; attribute dont_touch of I9575: signal is true;
	signal I9576: std_logic; attribute dont_touch of I9576: signal is true;
	signal I9581: std_logic; attribute dont_touch of I9581: signal is true;
	signal I9585: std_logic; attribute dont_touch of I9585: signal is true;
	signal I9588: std_logic; attribute dont_touch of I9588: signal is true;
	signal I9591: std_logic; attribute dont_touch of I9591: signal is true;
	signal I9594: std_logic; attribute dont_touch of I9594: signal is true;
	signal I9598: std_logic; attribute dont_touch of I9598: signal is true;
	signal I9602: std_logic; attribute dont_touch of I9602: signal is true;
	signal I9605: std_logic; attribute dont_touch of I9605: signal is true;
	signal I9608: std_logic; attribute dont_touch of I9608: signal is true;
	signal I9612: std_logic; attribute dont_touch of I9612: signal is true;
	signal I9617: std_logic; attribute dont_touch of I9617: signal is true;
	signal I9620: std_logic; attribute dont_touch of I9620: signal is true;
	signal I9625: std_logic; attribute dont_touch of I9625: signal is true;
	signal I9632: std_logic; attribute dont_touch of I9632: signal is true;
	signal I9639: std_logic; attribute dont_touch of I9639: signal is true;
	signal I9642: std_logic; attribute dont_touch of I9642: signal is true;
	signal I9647: std_logic; attribute dont_touch of I9647: signal is true;
	signal I9652: std_logic; attribute dont_touch of I9652: signal is true;
	signal I9655: std_logic; attribute dont_touch of I9655: signal is true;
	signal I9658: std_logic; attribute dont_touch of I9658: signal is true;
	signal I9662: std_logic; attribute dont_touch of I9662: signal is true;
	signal I9665: std_logic; attribute dont_touch of I9665: signal is true;
	signal I9669: std_logic; attribute dont_touch of I9669: signal is true;
	signal I9673: std_logic; attribute dont_touch of I9673: signal is true;
	signal I9677: std_logic; attribute dont_touch of I9677: signal is true;
	signal I9680: std_logic; attribute dont_touch of I9680: signal is true;
	signal I9684: std_logic; attribute dont_touch of I9684: signal is true;
	signal I9688: std_logic; attribute dont_touch of I9688: signal is true;
	signal I9695: std_logic; attribute dont_touch of I9695: signal is true;
	signal I9699: std_logic; attribute dont_touch of I9699: signal is true;
	signal I9706: std_logic; attribute dont_touch of I9706: signal is true;
	signal I9712: std_logic; attribute dont_touch of I9712: signal is true;
	signal I9717: std_logic; attribute dont_touch of I9717: signal is true;
	signal I9720: std_logic; attribute dont_touch of I9720: signal is true;
	signal I9727: std_logic; attribute dont_touch of I9727: signal is true;
	signal I9731: std_logic; attribute dont_touch of I9731: signal is true;
	signal I9734: std_logic; attribute dont_touch of I9734: signal is true;
	signal I9737: std_logic; attribute dont_touch of I9737: signal is true;
	signal I9744: std_logic; attribute dont_touch of I9744: signal is true;
	signal I9749: std_logic; attribute dont_touch of I9749: signal is true;
	signal I9754: std_logic; attribute dont_touch of I9754: signal is true;
	signal I9759: std_logic; attribute dont_touch of I9759: signal is true;
	signal I9762: std_logic; attribute dont_touch of I9762: signal is true;
	signal I9766: std_logic; attribute dont_touch of I9766: signal is true;
	signal I9769: std_logic; attribute dont_touch of I9769: signal is true;
	signal I9773: std_logic; attribute dont_touch of I9773: signal is true;
	signal I9776: std_logic; attribute dont_touch of I9776: signal is true;
	signal I9779: std_logic; attribute dont_touch of I9779: signal is true;
	signal I9783: std_logic; attribute dont_touch of I9783: signal is true;
	signal I9786: std_logic; attribute dont_touch of I9786: signal is true;
	signal I9789: std_logic; attribute dont_touch of I9789: signal is true;
	signal I9792: std_logic; attribute dont_touch of I9792: signal is true;
	signal I9795: std_logic; attribute dont_touch of I9795: signal is true;
	signal I9798: std_logic; attribute dont_touch of I9798: signal is true;
	signal I9801: std_logic; attribute dont_touch of I9801: signal is true;
	signal I9804: std_logic; attribute dont_touch of I9804: signal is true;
	signal I9807: std_logic; attribute dont_touch of I9807: signal is true;
	signal I9810: std_logic; attribute dont_touch of I9810: signal is true;
	signal I9813: std_logic; attribute dont_touch of I9813: signal is true;
	signal I9816: std_logic; attribute dont_touch of I9816: signal is true;
	signal I9822: std_logic; attribute dont_touch of I9822: signal is true;
	signal I9826: std_logic; attribute dont_touch of I9826: signal is true;
	signal I9829: std_logic; attribute dont_touch of I9829: signal is true;
	signal I9833: std_logic; attribute dont_touch of I9833: signal is true;
	signal I9836: std_logic; attribute dont_touch of I9836: signal is true;
	signal I9839: std_logic; attribute dont_touch of I9839: signal is true;
	signal I9842: std_logic; attribute dont_touch of I9842: signal is true;
	signal I9845: std_logic; attribute dont_touch of I9845: signal is true;
	signal I9848: std_logic; attribute dont_touch of I9848: signal is true;
	signal I9851: std_logic; attribute dont_touch of I9851: signal is true;
	signal I9854: std_logic; attribute dont_touch of I9854: signal is true;
	signal I9857: std_logic; attribute dont_touch of I9857: signal is true;
	signal I9860: std_logic; attribute dont_touch of I9860: signal is true;
	signal I9863: std_logic; attribute dont_touch of I9863: signal is true;
	signal I9866: std_logic; attribute dont_touch of I9866: signal is true;
	signal I9869: std_logic; attribute dont_touch of I9869: signal is true;
	signal I9872: std_logic; attribute dont_touch of I9872: signal is true;
	signal I9875: std_logic; attribute dont_touch of I9875: signal is true;
	signal I9880: std_logic; attribute dont_touch of I9880: signal is true;
	signal I9883: std_logic; attribute dont_touch of I9883: signal is true;
	signal I9886: std_logic; attribute dont_touch of I9886: signal is true;
	signal I9893: std_logic; attribute dont_touch of I9893: signal is true;
	signal I9896: std_logic; attribute dont_touch of I9896: signal is true;
	signal I9901: std_logic; attribute dont_touch of I9901: signal is true;
	signal I9905: std_logic; attribute dont_touch of I9905: signal is true;
	signal I9915: std_logic; attribute dont_touch of I9915: signal is true;
	signal I9923: std_logic; attribute dont_touch of I9923: signal is true;
	signal I9930: std_logic; attribute dont_touch of I9930: signal is true;
	signal I9935: std_logic; attribute dont_touch of I9935: signal is true;
	signal I9938: std_logic; attribute dont_touch of I9938: signal is true;
	signal I9946: std_logic; attribute dont_touch of I9946: signal is true;
	signal I9947: std_logic; attribute dont_touch of I9947: signal is true;
	signal I9948: std_logic; attribute dont_touch of I9948: signal is true;
	signal I9953: std_logic; attribute dont_touch of I9953: signal is true;
	signal I9956: std_logic; attribute dont_touch of I9956: signal is true;
	signal I9965: std_logic; attribute dont_touch of I9965: signal is true;
	signal I9973: std_logic; attribute dont_touch of I9973: signal is true;
	signal I9981: std_logic; attribute dont_touch of I9981: signal is true;
	signal I9984: std_logic; attribute dont_touch of I9984: signal is true;
	signal I9988: std_logic; attribute dont_touch of I9988: signal is true;
	signal I9992: std_logic; attribute dont_touch of I9992: signal is true;
	signal I9995: std_logic; attribute dont_touch of I9995: signal is true;
	signal I10003: std_logic; attribute dont_touch of I10003: signal is true;
	signal I10006: std_logic; attribute dont_touch of I10006: signal is true;
	signal I10009: std_logic; attribute dont_touch of I10009: signal is true;
	signal I10012: std_logic; attribute dont_touch of I10012: signal is true;
	signal I10015: std_logic; attribute dont_touch of I10015: signal is true;
	signal I10018: std_logic; attribute dont_touch of I10018: signal is true;
	signal I10021: std_logic; attribute dont_touch of I10021: signal is true;
	signal I10024: std_logic; attribute dont_touch of I10024: signal is true;
	signal I10027: std_logic; attribute dont_touch of I10027: signal is true;
	signal I10030: std_logic; attribute dont_touch of I10030: signal is true;
	signal I10033: std_logic; attribute dont_touch of I10033: signal is true;
	signal I10036: std_logic; attribute dont_touch of I10036: signal is true;
	signal I10039: std_logic; attribute dont_touch of I10039: signal is true;
	signal I10042: std_logic; attribute dont_touch of I10042: signal is true;
	signal I10045: std_logic; attribute dont_touch of I10045: signal is true;
	signal I10048: std_logic; attribute dont_touch of I10048: signal is true;
	signal I10051: std_logic; attribute dont_touch of I10051: signal is true;
	signal I10054: std_logic; attribute dont_touch of I10054: signal is true;
	signal I10057: std_logic; attribute dont_touch of I10057: signal is true;
	signal I10060: std_logic; attribute dont_touch of I10060: signal is true;
	signal I10063: std_logic; attribute dont_touch of I10063: signal is true;
	signal I10066: std_logic; attribute dont_touch of I10066: signal is true;
	signal I10069: std_logic; attribute dont_touch of I10069: signal is true;
	signal I10072: std_logic; attribute dont_touch of I10072: signal is true;
	signal I10075: std_logic; attribute dont_touch of I10075: signal is true;
	signal I10078: std_logic; attribute dont_touch of I10078: signal is true;
	signal I10081: std_logic; attribute dont_touch of I10081: signal is true;
	signal I10084: std_logic; attribute dont_touch of I10084: signal is true;
	signal I10087: std_logic; attribute dont_touch of I10087: signal is true;
	signal I10090: std_logic; attribute dont_touch of I10090: signal is true;
	signal I10093: std_logic; attribute dont_touch of I10093: signal is true;
	signal I10096: std_logic; attribute dont_touch of I10096: signal is true;
	signal I10099: std_logic; attribute dont_touch of I10099: signal is true;
	signal I10102: std_logic; attribute dont_touch of I10102: signal is true;
	signal I10105: std_logic; attribute dont_touch of I10105: signal is true;
	signal I10108: std_logic; attribute dont_touch of I10108: signal is true;
	signal I10111: std_logic; attribute dont_touch of I10111: signal is true;
	signal I10114: std_logic; attribute dont_touch of I10114: signal is true;
	signal I10117: std_logic; attribute dont_touch of I10117: signal is true;
	signal I10120: std_logic; attribute dont_touch of I10120: signal is true;
	signal I10123: std_logic; attribute dont_touch of I10123: signal is true;
	signal I10126: std_logic; attribute dont_touch of I10126: signal is true;
	signal I10129: std_logic; attribute dont_touch of I10129: signal is true;
	signal I10132: std_logic; attribute dont_touch of I10132: signal is true;
	signal I10135: std_logic; attribute dont_touch of I10135: signal is true;
	signal I10138: std_logic; attribute dont_touch of I10138: signal is true;
	signal I10141: std_logic; attribute dont_touch of I10141: signal is true;
	signal I10144: std_logic; attribute dont_touch of I10144: signal is true;
	signal I10147: std_logic; attribute dont_touch of I10147: signal is true;
	signal I10150: std_logic; attribute dont_touch of I10150: signal is true;
	signal I10153: std_logic; attribute dont_touch of I10153: signal is true;
	signal I10156: std_logic; attribute dont_touch of I10156: signal is true;
	signal I10159: std_logic; attribute dont_touch of I10159: signal is true;
	signal I10162: std_logic; attribute dont_touch of I10162: signal is true;
	signal I10165: std_logic; attribute dont_touch of I10165: signal is true;
	signal I10168: std_logic; attribute dont_touch of I10168: signal is true;
	signal I10171: std_logic; attribute dont_touch of I10171: signal is true;
	signal I10174: std_logic; attribute dont_touch of I10174: signal is true;
	signal I10177: std_logic; attribute dont_touch of I10177: signal is true;
	signal I10180: std_logic; attribute dont_touch of I10180: signal is true;
	signal I10183: std_logic; attribute dont_touch of I10183: signal is true;
	signal I10186: std_logic; attribute dont_touch of I10186: signal is true;
	signal I10189: std_logic; attribute dont_touch of I10189: signal is true;
	signal I10192: std_logic; attribute dont_touch of I10192: signal is true;
	signal I10195: std_logic; attribute dont_touch of I10195: signal is true;
	signal I10198: std_logic; attribute dont_touch of I10198: signal is true;
	signal I10201: std_logic; attribute dont_touch of I10201: signal is true;
	signal I10204: std_logic; attribute dont_touch of I10204: signal is true;
	signal I10221: std_logic; attribute dont_touch of I10221: signal is true;
	signal I10228: std_logic; attribute dont_touch of I10228: signal is true;
	signal I10231: std_logic; attribute dont_touch of I10231: signal is true;
	signal I10234: std_logic; attribute dont_touch of I10234: signal is true;
	signal I10237: std_logic; attribute dont_touch of I10237: signal is true;
	signal I10240: std_logic; attribute dont_touch of I10240: signal is true;
	signal I10243: std_logic; attribute dont_touch of I10243: signal is true;
	signal I10248: std_logic; attribute dont_touch of I10248: signal is true;
	signal I10251: std_logic; attribute dont_touch of I10251: signal is true;
	signal I10258: std_logic; attribute dont_touch of I10258: signal is true;
	signal I10274: std_logic; attribute dont_touch of I10274: signal is true;
	signal I10278: std_logic; attribute dont_touch of I10278: signal is true;
	signal I10282: std_logic; attribute dont_touch of I10282: signal is true;
	signal I10286: std_logic; attribute dont_touch of I10286: signal is true;
	signal I10289: std_logic; attribute dont_touch of I10289: signal is true;
	signal I10293: std_logic; attribute dont_touch of I10293: signal is true;
	signal I10296: std_logic; attribute dont_touch of I10296: signal is true;
	signal I10299: std_logic; attribute dont_touch of I10299: signal is true;
	signal I10302: std_logic; attribute dont_touch of I10302: signal is true;
	signal I10305: std_logic; attribute dont_touch of I10305: signal is true;
	signal I10308: std_logic; attribute dont_touch of I10308: signal is true;
	signal I10314: std_logic; attribute dont_touch of I10314: signal is true;
	signal I10317: std_logic; attribute dont_touch of I10317: signal is true;
	signal I10322: std_logic; attribute dont_touch of I10322: signal is true;
	signal I10325: std_logic; attribute dont_touch of I10325: signal is true;
	signal I10331: std_logic; attribute dont_touch of I10331: signal is true;
	signal I10334: std_logic; attribute dont_touch of I10334: signal is true;
	signal I10340: std_logic; attribute dont_touch of I10340: signal is true;
	signal I10343: std_logic; attribute dont_touch of I10343: signal is true;
	signal I10349: std_logic; attribute dont_touch of I10349: signal is true;
	signal I10352: std_logic; attribute dont_touch of I10352: signal is true;
	signal I10355: std_logic; attribute dont_touch of I10355: signal is true;
	signal I10362: std_logic; attribute dont_touch of I10362: signal is true;
	signal I10367: std_logic; attribute dont_touch of I10367: signal is true;
	signal I10370: std_logic; attribute dont_touch of I10370: signal is true;
	signal I10374: std_logic; attribute dont_touch of I10374: signal is true;
	signal I10378: std_logic; attribute dont_touch of I10378: signal is true;
	signal I10381: std_logic; attribute dont_touch of I10381: signal is true;
	signal I10384: std_logic; attribute dont_touch of I10384: signal is true;
	signal I10388: std_logic; attribute dont_touch of I10388: signal is true;
	signal I10391: std_logic; attribute dont_touch of I10391: signal is true;
	signal I10394: std_logic; attribute dont_touch of I10394: signal is true;
	signal I10398: std_logic; attribute dont_touch of I10398: signal is true;
	signal I10412: std_logic; attribute dont_touch of I10412: signal is true;
	signal I10421: std_logic; attribute dont_touch of I10421: signal is true;
	signal I10427: std_logic; attribute dont_touch of I10427: signal is true;
	signal I10434: std_logic; attribute dont_touch of I10434: signal is true;
	signal I10437: std_logic; attribute dont_touch of I10437: signal is true;
	signal I10445: std_logic; attribute dont_touch of I10445: signal is true;
	signal I10456: std_logic; attribute dont_touch of I10456: signal is true;
	signal I10461: std_logic; attribute dont_touch of I10461: signal is true;
	signal I10477: std_logic; attribute dont_touch of I10477: signal is true;
	signal I10484: std_logic; attribute dont_touch of I10484: signal is true;
	signal I10495: std_logic; attribute dont_touch of I10495: signal is true;
	signal I10499: std_logic; attribute dont_touch of I10499: signal is true;
	signal I10503: std_logic; attribute dont_touch of I10503: signal is true;
	signal I10507: std_logic; attribute dont_touch of I10507: signal is true;
	signal I10508: std_logic; attribute dont_touch of I10508: signal is true;
	signal I10509: std_logic; attribute dont_touch of I10509: signal is true;
	signal I10514: std_logic; attribute dont_touch of I10514: signal is true;
	signal I10519: std_logic; attribute dont_touch of I10519: signal is true;
	signal I10520: std_logic; attribute dont_touch of I10520: signal is true;
	signal I10521: std_logic; attribute dont_touch of I10521: signal is true;
	signal I10526: std_logic; attribute dont_touch of I10526: signal is true;
	signal I10531: std_logic; attribute dont_touch of I10531: signal is true;
	signal I10535: std_logic; attribute dont_touch of I10535: signal is true;
	signal I10538: std_logic; attribute dont_touch of I10538: signal is true;
	signal I10541: std_logic; attribute dont_touch of I10541: signal is true;
	signal I10546: std_logic; attribute dont_touch of I10546: signal is true;
	signal I10549: std_logic; attribute dont_touch of I10549: signal is true;
	signal I10553: std_logic; attribute dont_touch of I10553: signal is true;
	signal I10557: std_logic; attribute dont_touch of I10557: signal is true;
	signal I10560: std_logic; attribute dont_touch of I10560: signal is true;
	signal I10563: std_logic; attribute dont_touch of I10563: signal is true;
	signal I10566: std_logic; attribute dont_touch of I10566: signal is true;
	signal I10573: std_logic; attribute dont_touch of I10573: signal is true;
	signal I10584: std_logic; attribute dont_touch of I10584: signal is true;
	signal I10589: std_logic; attribute dont_touch of I10589: signal is true;
	signal I10592: std_logic; attribute dont_touch of I10592: signal is true;
	signal I10598: std_logic; attribute dont_touch of I10598: signal is true;
	signal I10601: std_logic; attribute dont_touch of I10601: signal is true;
	signal I10607: std_logic; attribute dont_touch of I10607: signal is true;
	signal I10610: std_logic; attribute dont_touch of I10610: signal is true;
	signal I10613: std_logic; attribute dont_touch of I10613: signal is true;
	signal I10620: std_logic; attribute dont_touch of I10620: signal is true;
	signal I10623: std_logic; attribute dont_touch of I10623: signal is true;
	signal I10630: std_logic; attribute dont_touch of I10630: signal is true;
	signal I10633: std_logic; attribute dont_touch of I10633: signal is true;
	signal I10639: std_logic; attribute dont_touch of I10639: signal is true;
	signal I10643: std_logic; attribute dont_touch of I10643: signal is true;
	signal I10648: std_logic; attribute dont_touch of I10648: signal is true;
	signal I10651: std_logic; attribute dont_touch of I10651: signal is true;
	signal I10655: std_logic; attribute dont_touch of I10655: signal is true;
	signal I10659: std_logic; attribute dont_touch of I10659: signal is true;
	signal I10663: std_logic; attribute dont_touch of I10663: signal is true;
	signal I10666: std_logic; attribute dont_touch of I10666: signal is true;
	signal I10671: std_logic; attribute dont_touch of I10671: signal is true;
	signal I10678: std_logic; attribute dont_touch of I10678: signal is true;
	signal I10682: std_logic; attribute dont_touch of I10682: signal is true;
	signal I10685: std_logic; attribute dont_touch of I10685: signal is true;
	signal I10689: std_logic; attribute dont_touch of I10689: signal is true;
	signal I10693: std_logic; attribute dont_touch of I10693: signal is true;
	signal I10698: std_logic; attribute dont_touch of I10698: signal is true;
	signal I10702: std_logic; attribute dont_touch of I10702: signal is true;
	signal I10706: std_logic; attribute dont_touch of I10706: signal is true;
	signal I10710: std_logic; attribute dont_touch of I10710: signal is true;
	signal I10713: std_logic; attribute dont_touch of I10713: signal is true;
	signal I10716: std_logic; attribute dont_touch of I10716: signal is true;
	signal I10719: std_logic; attribute dont_touch of I10719: signal is true;
	signal I10724: std_logic; attribute dont_touch of I10724: signal is true;
	signal I10729: std_logic; attribute dont_touch of I10729: signal is true;
	signal I10733: std_logic; attribute dont_touch of I10733: signal is true;
	signal I10736: std_logic; attribute dont_touch of I10736: signal is true;
	signal I10739: std_logic; attribute dont_touch of I10739: signal is true;
	signal I10753: std_logic; attribute dont_touch of I10753: signal is true;
	signal I10756: std_logic; attribute dont_touch of I10756: signal is true;
	signal I10759: std_logic; attribute dont_touch of I10759: signal is true;
	signal I10762: std_logic; attribute dont_touch of I10762: signal is true;
	signal I10769: std_logic; attribute dont_touch of I10769: signal is true;
	signal I10770: std_logic; attribute dont_touch of I10770: signal is true;
	signal I10771: std_logic; attribute dont_touch of I10771: signal is true;
	signal I10789: std_logic; attribute dont_touch of I10789: signal is true;
	signal I10795: std_logic; attribute dont_touch of I10795: signal is true;
	signal I10801: std_logic; attribute dont_touch of I10801: signal is true;
	signal I10804: std_logic; attribute dont_touch of I10804: signal is true;
	signal I10807: std_logic; attribute dont_touch of I10807: signal is true;
	signal I10810: std_logic; attribute dont_touch of I10810: signal is true;
	signal I10813: std_logic; attribute dont_touch of I10813: signal is true;
	signal I10816: std_logic; attribute dont_touch of I10816: signal is true;
	signal I10819: std_logic; attribute dont_touch of I10819: signal is true;
	signal I10822: std_logic; attribute dont_touch of I10822: signal is true;
	signal I10825: std_logic; attribute dont_touch of I10825: signal is true;
	signal I10828: std_logic; attribute dont_touch of I10828: signal is true;
	signal I10831: std_logic; attribute dont_touch of I10831: signal is true;
	signal I10834: std_logic; attribute dont_touch of I10834: signal is true;
	signal I10837: std_logic; attribute dont_touch of I10837: signal is true;
	signal I10840: std_logic; attribute dont_touch of I10840: signal is true;
	signal I10843: std_logic; attribute dont_touch of I10843: signal is true;
	signal I10846: std_logic; attribute dont_touch of I10846: signal is true;
	signal I10849: std_logic; attribute dont_touch of I10849: signal is true;
	signal I10852: std_logic; attribute dont_touch of I10852: signal is true;
	signal I10855: std_logic; attribute dont_touch of I10855: signal is true;
	signal I10858: std_logic; attribute dont_touch of I10858: signal is true;
	signal I10861: std_logic; attribute dont_touch of I10861: signal is true;
	signal I10864: std_logic; attribute dont_touch of I10864: signal is true;
	signal I10873: std_logic; attribute dont_touch of I10873: signal is true;
	signal I10885: std_logic; attribute dont_touch of I10885: signal is true;
	signal I10888: std_logic; attribute dont_touch of I10888: signal is true;
	signal I10891: std_logic; attribute dont_touch of I10891: signal is true;
	signal I10898: std_logic; attribute dont_touch of I10898: signal is true;
	signal I10901: std_logic; attribute dont_touch of I10901: signal is true;
	signal I10904: std_logic; attribute dont_touch of I10904: signal is true;
	signal I10907: std_logic; attribute dont_touch of I10907: signal is true;
	signal I10910: std_logic; attribute dont_touch of I10910: signal is true;
	signal I10914: std_logic; attribute dont_touch of I10914: signal is true;
	signal I10917: std_logic; attribute dont_touch of I10917: signal is true;
	signal I10920: std_logic; attribute dont_touch of I10920: signal is true;
	signal I10924: std_logic; attribute dont_touch of I10924: signal is true;
	signal I10927: std_logic; attribute dont_touch of I10927: signal is true;
	signal I10930: std_logic; attribute dont_touch of I10930: signal is true;
	signal I10931: std_logic; attribute dont_touch of I10931: signal is true;
	signal I10932: std_logic; attribute dont_touch of I10932: signal is true;
	signal I10937: std_logic; attribute dont_touch of I10937: signal is true;
	signal I10941: std_logic; attribute dont_touch of I10941: signal is true;
	signal I10946: std_logic; attribute dont_touch of I10946: signal is true;
	signal I10949: std_logic; attribute dont_touch of I10949: signal is true;
	signal I10952: std_logic; attribute dont_touch of I10952: signal is true;
	signal I10958: std_logic; attribute dont_touch of I10958: signal is true;
	signal I10963: std_logic; attribute dont_touch of I10963: signal is true;
	signal I10966: std_logic; attribute dont_touch of I10966: signal is true;
	signal I10971: std_logic; attribute dont_touch of I10971: signal is true;
	signal I10974: std_logic; attribute dont_touch of I10974: signal is true;
	signal I10979: std_logic; attribute dont_touch of I10979: signal is true;
	signal I10984: std_logic; attribute dont_touch of I10984: signal is true;
	signal I10991: std_logic; attribute dont_touch of I10991: signal is true;
	signal I10996: std_logic; attribute dont_touch of I10996: signal is true;
	signal I11005: std_logic; attribute dont_touch of I11005: signal is true;
	signal I11008: std_logic; attribute dont_touch of I11008: signal is true;
	signal I11011: std_logic; attribute dont_touch of I11011: signal is true;
	signal I11021: std_logic; attribute dont_touch of I11021: signal is true;
	signal I11024: std_logic; attribute dont_touch of I11024: signal is true;
	signal I11029: std_logic; attribute dont_touch of I11029: signal is true;
	signal I11034: std_logic; attribute dont_touch of I11034: signal is true;
	signal I11037: std_logic; attribute dont_touch of I11037: signal is true;
	signal I11043: std_logic; attribute dont_touch of I11043: signal is true;
	signal I11046: std_logic; attribute dont_touch of I11046: signal is true;
	signal I11049: std_logic; attribute dont_touch of I11049: signal is true;
	signal I11055: std_logic; attribute dont_touch of I11055: signal is true;
	signal I11058: std_logic; attribute dont_touch of I11058: signal is true;
	signal I11061: std_logic; attribute dont_touch of I11061: signal is true;
	signal I11065: std_logic; attribute dont_touch of I11065: signal is true;
	signal I11068: std_logic; attribute dont_touch of I11068: signal is true;
	signal I11071: std_logic; attribute dont_touch of I11071: signal is true;
	signal I11076: std_logic; attribute dont_touch of I11076: signal is true;
	signal I11079: std_logic; attribute dont_touch of I11079: signal is true;
	signal I11082: std_logic; attribute dont_touch of I11082: signal is true;
	signal I11085: std_logic; attribute dont_touch of I11085: signal is true;
	signal I11088: std_logic; attribute dont_touch of I11088: signal is true;
	signal I11091: std_logic; attribute dont_touch of I11091: signal is true;
	signal I11094: std_logic; attribute dont_touch of I11094: signal is true;
	signal I11097: std_logic; attribute dont_touch of I11097: signal is true;
	signal I11100: std_logic; attribute dont_touch of I11100: signal is true;
	signal I11103: std_logic; attribute dont_touch of I11103: signal is true;
	signal I11106: std_logic; attribute dont_touch of I11106: signal is true;
	signal I11109: std_logic; attribute dont_touch of I11109: signal is true;
	signal I11112: std_logic; attribute dont_touch of I11112: signal is true;
	signal I11115: std_logic; attribute dont_touch of I11115: signal is true;
	signal I11119: std_logic; attribute dont_touch of I11119: signal is true;
	signal I11122: std_logic; attribute dont_touch of I11122: signal is true;
	signal I11127: std_logic; attribute dont_touch of I11127: signal is true;
	signal I11132: std_logic; attribute dont_touch of I11132: signal is true;
	signal I11135: std_logic; attribute dont_touch of I11135: signal is true;
	signal I11140: std_logic; attribute dont_touch of I11140: signal is true;
	signal I11143: std_logic; attribute dont_touch of I11143: signal is true;
	signal I11146: std_logic; attribute dont_touch of I11146: signal is true;
	signal I11149: std_logic; attribute dont_touch of I11149: signal is true;
	signal I11152: std_logic; attribute dont_touch of I11152: signal is true;
	signal I11155: std_logic; attribute dont_touch of I11155: signal is true;
	signal I11159: std_logic; attribute dont_touch of I11159: signal is true;
	signal I11162: std_logic; attribute dont_touch of I11162: signal is true;
	signal I11166: std_logic; attribute dont_touch of I11166: signal is true;
	signal I11169: std_logic; attribute dont_touch of I11169: signal is true;
	signal I11173: std_logic; attribute dont_touch of I11173: signal is true;
	signal I11176: std_logic; attribute dont_touch of I11176: signal is true;
	signal I11180: std_logic; attribute dont_touch of I11180: signal is true;
	signal I11183: std_logic; attribute dont_touch of I11183: signal is true;
	signal I11188: std_logic; attribute dont_touch of I11188: signal is true;
	signal I11191: std_logic; attribute dont_touch of I11191: signal is true;
	signal I11194: std_logic; attribute dont_touch of I11194: signal is true;
	signal I11198: std_logic; attribute dont_touch of I11198: signal is true;
	signal I11201: std_logic; attribute dont_touch of I11201: signal is true;
	signal I11204: std_logic; attribute dont_touch of I11204: signal is true;
	signal I11207: std_logic; attribute dont_touch of I11207: signal is true;
	signal I11211: std_logic; attribute dont_touch of I11211: signal is true;
	signal I11214: std_logic; attribute dont_touch of I11214: signal is true;
	signal I11217: std_logic; attribute dont_touch of I11217: signal is true;
	signal I11222: std_logic; attribute dont_touch of I11222: signal is true;
	signal I11225: std_logic; attribute dont_touch of I11225: signal is true;
	signal I11228: std_logic; attribute dont_touch of I11228: signal is true;
	signal I11232: std_logic; attribute dont_touch of I11232: signal is true;
	signal I11235: std_logic; attribute dont_touch of I11235: signal is true;
	signal I11238: std_logic; attribute dont_touch of I11238: signal is true;
	signal I11241: std_logic; attribute dont_touch of I11241: signal is true;
	signal I11242: std_logic; attribute dont_touch of I11242: signal is true;
	signal I11243: std_logic; attribute dont_touch of I11243: signal is true;
	signal I11249: std_logic; attribute dont_touch of I11249: signal is true;
	signal I11252: std_logic; attribute dont_touch of I11252: signal is true;
	signal I11255: std_logic; attribute dont_touch of I11255: signal is true;
	signal I11261: std_logic; attribute dont_touch of I11261: signal is true;
	signal I11262: std_logic; attribute dont_touch of I11262: signal is true;
	signal I11263: std_logic; attribute dont_touch of I11263: signal is true;
	signal I11269: std_logic; attribute dont_touch of I11269: signal is true;
	signal I11272: std_logic; attribute dont_touch of I11272: signal is true;
	signal I11275: std_logic; attribute dont_touch of I11275: signal is true;
	signal I11278: std_logic; attribute dont_touch of I11278: signal is true;
	signal I11279: std_logic; attribute dont_touch of I11279: signal is true;
	signal I11280: std_logic; attribute dont_touch of I11280: signal is true;
	signal I11286: std_logic; attribute dont_touch of I11286: signal is true;
	signal I11289: std_logic; attribute dont_touch of I11289: signal is true;
	signal I11293: std_logic; attribute dont_touch of I11293: signal is true;
	signal I11296: std_logic; attribute dont_touch of I11296: signal is true;
	signal I11299: std_logic; attribute dont_touch of I11299: signal is true;
	signal I11303: std_logic; attribute dont_touch of I11303: signal is true;
	signal I11306: std_logic; attribute dont_touch of I11306: signal is true;
	signal I11309: std_logic; attribute dont_touch of I11309: signal is true;
	signal I11312: std_logic; attribute dont_touch of I11312: signal is true;
	signal I11315: std_logic; attribute dont_touch of I11315: signal is true;
	signal I11318: std_logic; attribute dont_touch of I11318: signal is true;
	signal I11322: std_logic; attribute dont_touch of I11322: signal is true;
	signal I11326: std_logic; attribute dont_touch of I11326: signal is true;
	signal I11330: std_logic; attribute dont_touch of I11330: signal is true;
	signal I11333: std_logic; attribute dont_touch of I11333: signal is true;
	signal I11338: std_logic; attribute dont_touch of I11338: signal is true;
	signal I11342: std_logic; attribute dont_touch of I11342: signal is true;
	signal I11345: std_logic; attribute dont_touch of I11345: signal is true;
	signal I11348: std_logic; attribute dont_touch of I11348: signal is true;
	signal I11351: std_logic; attribute dont_touch of I11351: signal is true;
	signal I11354: std_logic; attribute dont_touch of I11354: signal is true;
	signal I11357: std_logic; attribute dont_touch of I11357: signal is true;
	signal I11360: std_logic; attribute dont_touch of I11360: signal is true;
	signal I11363: std_logic; attribute dont_touch of I11363: signal is true;
	signal I11367: std_logic; attribute dont_touch of I11367: signal is true;
	signal I11383: std_logic; attribute dont_touch of I11383: signal is true;
	signal I11387: std_logic; attribute dont_touch of I11387: signal is true;
	signal I11391: std_logic; attribute dont_touch of I11391: signal is true;
	signal I11394: std_logic; attribute dont_touch of I11394: signal is true;
	signal I11397: std_logic; attribute dont_touch of I11397: signal is true;
	signal I11405: std_logic; attribute dont_touch of I11405: signal is true;
	signal I11408: std_logic; attribute dont_touch of I11408: signal is true;
	signal I11412: std_logic; attribute dont_touch of I11412: signal is true;
	signal I11417: std_logic; attribute dont_touch of I11417: signal is true;
	signal I11420: std_logic; attribute dont_touch of I11420: signal is true;
	signal I11423: std_logic; attribute dont_touch of I11423: signal is true;
	signal I11427: std_logic; attribute dont_touch of I11427: signal is true;
	signal I11433: std_logic; attribute dont_touch of I11433: signal is true;
	signal I11436: std_logic; attribute dont_touch of I11436: signal is true;
	signal I11440: std_logic; attribute dont_touch of I11440: signal is true;
	signal I11444: std_logic; attribute dont_touch of I11444: signal is true;
	signal I11447: std_logic; attribute dont_touch of I11447: signal is true;
	signal I11450: std_logic; attribute dont_touch of I11450: signal is true;
	signal I11456: std_logic; attribute dont_touch of I11456: signal is true;
	signal I11459: std_logic; attribute dont_touch of I11459: signal is true;
	signal I11464: std_logic; attribute dont_touch of I11464: signal is true;
	signal I11467: std_logic; attribute dont_touch of I11467: signal is true;
	signal I11472: std_logic; attribute dont_touch of I11472: signal is true;
	signal I11477: std_logic; attribute dont_touch of I11477: signal is true;
	signal I11483: std_logic; attribute dont_touch of I11483: signal is true;
	signal I11489: std_logic; attribute dont_touch of I11489: signal is true;
	signal I11494: std_logic; attribute dont_touch of I11494: signal is true;
	signal I11498: std_logic; attribute dont_touch of I11498: signal is true;
	signal I11501: std_logic; attribute dont_touch of I11501: signal is true;
	signal I11505: std_logic; attribute dont_touch of I11505: signal is true;
	signal I11508: std_logic; attribute dont_touch of I11508: signal is true;
	signal I11509: std_logic; attribute dont_touch of I11509: signal is true;
	signal I11510: std_logic; attribute dont_touch of I11510: signal is true;
	signal I11515: std_logic; attribute dont_touch of I11515: signal is true;
	signal I11519: std_logic; attribute dont_touch of I11519: signal is true;
	signal I11524: std_logic; attribute dont_touch of I11524: signal is true;
	signal I11528: std_logic; attribute dont_touch of I11528: signal is true;
	signal I11531: std_logic; attribute dont_touch of I11531: signal is true;
	signal I11534: std_logic; attribute dont_touch of I11534: signal is true;
	signal I11537: std_logic; attribute dont_touch of I11537: signal is true;
	signal I11540: std_logic; attribute dont_touch of I11540: signal is true;
	signal I11543: std_logic; attribute dont_touch of I11543: signal is true;
	signal I11560: std_logic; attribute dont_touch of I11560: signal is true;
	signal I11563: std_logic; attribute dont_touch of I11563: signal is true;
	signal I11566: std_logic; attribute dont_touch of I11566: signal is true;
	signal I11569: std_logic; attribute dont_touch of I11569: signal is true;
	signal I11572: std_logic; attribute dont_touch of I11572: signal is true;
	signal I11575: std_logic; attribute dont_touch of I11575: signal is true;
	signal I11578: std_logic; attribute dont_touch of I11578: signal is true;
	signal I11581: std_logic; attribute dont_touch of I11581: signal is true;
	signal I11584: std_logic; attribute dont_touch of I11584: signal is true;
	signal I11587: std_logic; attribute dont_touch of I11587: signal is true;
	signal I11590: std_logic; attribute dont_touch of I11590: signal is true;
	signal I11593: std_logic; attribute dont_touch of I11593: signal is true;
	signal I11596: std_logic; attribute dont_touch of I11596: signal is true;
	signal I11599: std_logic; attribute dont_touch of I11599: signal is true;
	signal I11602: std_logic; attribute dont_touch of I11602: signal is true;
	signal I11605: std_logic; attribute dont_touch of I11605: signal is true;
	signal I11608: std_logic; attribute dont_touch of I11608: signal is true;
	signal I11611: std_logic; attribute dont_touch of I11611: signal is true;
	signal I11614: std_logic; attribute dont_touch of I11614: signal is true;
	signal I11617: std_logic; attribute dont_touch of I11617: signal is true;
	signal I11620: std_logic; attribute dont_touch of I11620: signal is true;
	signal I11623: std_logic; attribute dont_touch of I11623: signal is true;
	signal I11626: std_logic; attribute dont_touch of I11626: signal is true;
	signal I11629: std_logic; attribute dont_touch of I11629: signal is true;
	signal I11632: std_logic; attribute dont_touch of I11632: signal is true;
	signal I11635: std_logic; attribute dont_touch of I11635: signal is true;
	signal I11638: std_logic; attribute dont_touch of I11638: signal is true;
	signal I11641: std_logic; attribute dont_touch of I11641: signal is true;
	signal I11644: std_logic; attribute dont_touch of I11644: signal is true;
	signal I11647: std_logic; attribute dont_touch of I11647: signal is true;
	signal I11650: std_logic; attribute dont_touch of I11650: signal is true;
	signal I11653: std_logic; attribute dont_touch of I11653: signal is true;
	signal I11656: std_logic; attribute dont_touch of I11656: signal is true;
	signal I11659: std_logic; attribute dont_touch of I11659: signal is true;
	signal I11662: std_logic; attribute dont_touch of I11662: signal is true;
	signal I11665: std_logic; attribute dont_touch of I11665: signal is true;
	signal I11668: std_logic; attribute dont_touch of I11668: signal is true;
	signal I11671: std_logic; attribute dont_touch of I11671: signal is true;
	signal I11674: std_logic; attribute dont_touch of I11674: signal is true;
	signal I11677: std_logic; attribute dont_touch of I11677: signal is true;
	signal I11680: std_logic; attribute dont_touch of I11680: signal is true;
	signal I11683: std_logic; attribute dont_touch of I11683: signal is true;
	signal I11686: std_logic; attribute dont_touch of I11686: signal is true;
	signal I11689: std_logic; attribute dont_touch of I11689: signal is true;
	signal I11692: std_logic; attribute dont_touch of I11692: signal is true;
	signal I11695: std_logic; attribute dont_touch of I11695: signal is true;
	signal I11698: std_logic; attribute dont_touch of I11698: signal is true;
	signal I11701: std_logic; attribute dont_touch of I11701: signal is true;
	signal I11704: std_logic; attribute dont_touch of I11704: signal is true;
	signal I11707: std_logic; attribute dont_touch of I11707: signal is true;
	signal I11710: std_logic; attribute dont_touch of I11710: signal is true;
	signal I11713: std_logic; attribute dont_touch of I11713: signal is true;
	signal I11716: std_logic; attribute dont_touch of I11716: signal is true;
	signal I11719: std_logic; attribute dont_touch of I11719: signal is true;
	signal I11722: std_logic; attribute dont_touch of I11722: signal is true;
	signal I11725: std_logic; attribute dont_touch of I11725: signal is true;
	signal I11728: std_logic; attribute dont_touch of I11728: signal is true;
	signal I11731: std_logic; attribute dont_touch of I11731: signal is true;
	signal I11734: std_logic; attribute dont_touch of I11734: signal is true;
	signal I11737: std_logic; attribute dont_touch of I11737: signal is true;
	signal I11740: std_logic; attribute dont_touch of I11740: signal is true;
	signal I11743: std_logic; attribute dont_touch of I11743: signal is true;
	signal I11746: std_logic; attribute dont_touch of I11746: signal is true;
	signal I11752: std_logic; attribute dont_touch of I11752: signal is true;
	signal I11756: std_logic; attribute dont_touch of I11756: signal is true;
	signal I11759: std_logic; attribute dont_touch of I11759: signal is true;
	signal I11767: std_logic; attribute dont_touch of I11767: signal is true;
	signal I11770: std_logic; attribute dont_touch of I11770: signal is true;
	signal I11773: std_logic; attribute dont_touch of I11773: signal is true;
	signal I11778: std_logic; attribute dont_touch of I11778: signal is true;
	signal I11783: std_logic; attribute dont_touch of I11783: signal is true;
	signal I11786: std_logic; attribute dont_touch of I11786: signal is true;
	signal I11790: std_logic; attribute dont_touch of I11790: signal is true;
	signal I11794: std_logic; attribute dont_touch of I11794: signal is true;
	signal I11797: std_logic; attribute dont_touch of I11797: signal is true;
	signal I11800: std_logic; attribute dont_touch of I11800: signal is true;
	signal I11804: std_logic; attribute dont_touch of I11804: signal is true;
	signal I11807: std_logic; attribute dont_touch of I11807: signal is true;
	signal I11810: std_logic; attribute dont_touch of I11810: signal is true;
	signal I11814: std_logic; attribute dont_touch of I11814: signal is true;
	signal I11817: std_logic; attribute dont_touch of I11817: signal is true;
	signal I11821: std_logic; attribute dont_touch of I11821: signal is true;
	signal I11824: std_logic; attribute dont_touch of I11824: signal is true;
	signal I11829: std_logic; attribute dont_touch of I11829: signal is true;
	signal I11833: std_logic; attribute dont_touch of I11833: signal is true;
	signal I11836: std_logic; attribute dont_touch of I11836: signal is true;
	signal I11841: std_logic; attribute dont_touch of I11841: signal is true;
	signal I11845: std_logic; attribute dont_touch of I11845: signal is true;
	signal I11858: std_logic; attribute dont_touch of I11858: signal is true;
	signal I11869: std_logic; attribute dont_touch of I11869: signal is true;
	signal I11873: std_logic; attribute dont_touch of I11873: signal is true;
	signal I11879: std_logic; attribute dont_touch of I11879: signal is true;
	signal I11882: std_logic; attribute dont_touch of I11882: signal is true;
	signal I11889: std_logic; attribute dont_touch of I11889: signal is true;
	signal I11898: std_logic; attribute dont_touch of I11898: signal is true;
	signal I11901: std_logic; attribute dont_touch of I11901: signal is true;
	signal I11904: std_logic; attribute dont_touch of I11904: signal is true;
	signal I11907: std_logic; attribute dont_touch of I11907: signal is true;
	signal I11908: std_logic; attribute dont_touch of I11908: signal is true;
	signal I11909: std_logic; attribute dont_touch of I11909: signal is true;
	signal I11914: std_logic; attribute dont_touch of I11914: signal is true;
	signal I11915: std_logic; attribute dont_touch of I11915: signal is true;
	signal I11916: std_logic; attribute dont_touch of I11916: signal is true;
	signal I11921: std_logic; attribute dont_touch of I11921: signal is true;
	signal I11926: std_logic; attribute dont_touch of I11926: signal is true;
	signal I11929: std_logic; attribute dont_touch of I11929: signal is true;
	signal I11932: std_logic; attribute dont_touch of I11932: signal is true;
	signal I11935: std_logic; attribute dont_touch of I11935: signal is true;
	signal I11936: std_logic; attribute dont_touch of I11936: signal is true;
	signal I11937: std_logic; attribute dont_touch of I11937: signal is true;
	signal I11942: std_logic; attribute dont_touch of I11942: signal is true;
	signal I11947: std_logic; attribute dont_touch of I11947: signal is true;
	signal I11950: std_logic; attribute dont_touch of I11950: signal is true;
	signal I11953: std_logic; attribute dont_touch of I11953: signal is true;
	signal I11956: std_logic; attribute dont_touch of I11956: signal is true;
	signal I11961: std_logic; attribute dont_touch of I11961: signal is true;
	signal I11964: std_logic; attribute dont_touch of I11964: signal is true;
	signal I11967: std_logic; attribute dont_touch of I11967: signal is true;
	signal I11970: std_logic; attribute dont_touch of I11970: signal is true;
	signal I11973: std_logic; attribute dont_touch of I11973: signal is true;
	signal I11974: std_logic; attribute dont_touch of I11974: signal is true;
	signal I11975: std_logic; attribute dont_touch of I11975: signal is true;
	signal I11980: std_logic; attribute dont_touch of I11980: signal is true;
	signal I11981: std_logic; attribute dont_touch of I11981: signal is true;
	signal I11982: std_logic; attribute dont_touch of I11982: signal is true;
	signal I11989: std_logic; attribute dont_touch of I11989: signal is true;
	signal I11992: std_logic; attribute dont_touch of I11992: signal is true;
	signal I11995: std_logic; attribute dont_touch of I11995: signal is true;
	signal I11996: std_logic; attribute dont_touch of I11996: signal is true;
	signal I11997: std_logic; attribute dont_touch of I11997: signal is true;
	signal I12002: std_logic; attribute dont_touch of I12002: signal is true;
	signal I12003: std_logic; attribute dont_touch of I12003: signal is true;
	signal I12004: std_logic; attribute dont_touch of I12004: signal is true;
	signal I12009: std_logic; attribute dont_touch of I12009: signal is true;
	signal I12012: std_logic; attribute dont_touch of I12012: signal is true;
	signal I12015: std_logic; attribute dont_touch of I12015: signal is true;
	signal I12019: std_logic; attribute dont_touch of I12019: signal is true;
	signal I12020: std_logic; attribute dont_touch of I12020: signal is true;
	signal I12021: std_logic; attribute dont_touch of I12021: signal is true;
	signal I12026: std_logic; attribute dont_touch of I12026: signal is true;
	signal I12029: std_logic; attribute dont_touch of I12029: signal is true;
	signal I12032: std_logic; attribute dont_touch of I12032: signal is true;
	signal I12035: std_logic; attribute dont_touch of I12035: signal is true;
	signal I12038: std_logic; attribute dont_touch of I12038: signal is true;
	signal I12039: std_logic; attribute dont_touch of I12039: signal is true;
	signal I12040: std_logic; attribute dont_touch of I12040: signal is true;
	signal I12045: std_logic; attribute dont_touch of I12045: signal is true;
	signal I12046: std_logic; attribute dont_touch of I12046: signal is true;
	signal I12047: std_logic; attribute dont_touch of I12047: signal is true;
	signal I12053: std_logic; attribute dont_touch of I12053: signal is true;
	signal I12056: std_logic; attribute dont_touch of I12056: signal is true;
	signal I12060: std_logic; attribute dont_touch of I12060: signal is true;
	signal I12061: std_logic; attribute dont_touch of I12061: signal is true;
	signal I12062: std_logic; attribute dont_touch of I12062: signal is true;
	signal I12067: std_logic; attribute dont_touch of I12067: signal is true;
	signal I12068: std_logic; attribute dont_touch of I12068: signal is true;
	signal I12069: std_logic; attribute dont_touch of I12069: signal is true;
	signal I12074: std_logic; attribute dont_touch of I12074: signal is true;
	signal I12075: std_logic; attribute dont_touch of I12075: signal is true;
	signal I12076: std_logic; attribute dont_touch of I12076: signal is true;
	signal I12081: std_logic; attribute dont_touch of I12081: signal is true;
	signal I12085: std_logic; attribute dont_touch of I12085: signal is true;
	signal I12086: std_logic; attribute dont_touch of I12086: signal is true;
	signal I12087: std_logic; attribute dont_touch of I12087: signal is true;
	signal I12092: std_logic; attribute dont_touch of I12092: signal is true;
	signal I12093: std_logic; attribute dont_touch of I12093: signal is true;
	signal I12094: std_logic; attribute dont_touch of I12094: signal is true;
	signal I12099: std_logic; attribute dont_touch of I12099: signal is true;
	signal I12103: std_logic; attribute dont_touch of I12103: signal is true;
	signal I12106: std_logic; attribute dont_touch of I12106: signal is true;
	signal I12107: std_logic; attribute dont_touch of I12107: signal is true;
	signal I12108: std_logic; attribute dont_touch of I12108: signal is true;
	signal I12113: std_logic; attribute dont_touch of I12113: signal is true;
	signal I12114: std_logic; attribute dont_touch of I12114: signal is true;
	signal I12115: std_logic; attribute dont_touch of I12115: signal is true;
	signal I12120: std_logic; attribute dont_touch of I12120: signal is true;
	signal I12123: std_logic; attribute dont_touch of I12123: signal is true;
	signal I12126: std_logic; attribute dont_touch of I12126: signal is true;
	signal I12127: std_logic; attribute dont_touch of I12127: signal is true;
	signal I12128: std_logic; attribute dont_touch of I12128: signal is true;
	signal I12133: std_logic; attribute dont_touch of I12133: signal is true;
	signal I12136: std_logic; attribute dont_touch of I12136: signal is true;
	signal I12137: std_logic; attribute dont_touch of I12137: signal is true;
	signal I12138: std_logic; attribute dont_touch of I12138: signal is true;
	signal I12143: std_logic; attribute dont_touch of I12143: signal is true;
	signal I12144: std_logic; attribute dont_touch of I12144: signal is true;
	signal I12145: std_logic; attribute dont_touch of I12145: signal is true;
	signal I12150: std_logic; attribute dont_touch of I12150: signal is true;
	signal I12153: std_logic; attribute dont_touch of I12153: signal is true;
	signal I12156: std_logic; attribute dont_touch of I12156: signal is true;
	signal I12159: std_logic; attribute dont_touch of I12159: signal is true;
	signal I12162: std_logic; attribute dont_touch of I12162: signal is true;
	signal I12165: std_logic; attribute dont_touch of I12165: signal is true;
	signal I12168: std_logic; attribute dont_touch of I12168: signal is true;
	signal I12171: std_logic; attribute dont_touch of I12171: signal is true;
	signal I12174: std_logic; attribute dont_touch of I12174: signal is true;
	signal I12177: std_logic; attribute dont_touch of I12177: signal is true;
	signal I12180: std_logic; attribute dont_touch of I12180: signal is true;
	signal I12183: std_logic; attribute dont_touch of I12183: signal is true;
	signal I12186: std_logic; attribute dont_touch of I12186: signal is true;
	signal I12190: std_logic; attribute dont_touch of I12190: signal is true;
	signal I12193: std_logic; attribute dont_touch of I12193: signal is true;
	signal I12196: std_logic; attribute dont_touch of I12196: signal is true;
	signal I12199: std_logic; attribute dont_touch of I12199: signal is true;
	signal I12202: std_logic; attribute dont_touch of I12202: signal is true;
	signal I12205: std_logic; attribute dont_touch of I12205: signal is true;
	signal I12208: std_logic; attribute dont_touch of I12208: signal is true;
	signal I12214: std_logic; attribute dont_touch of I12214: signal is true;
	signal I12215: std_logic; attribute dont_touch of I12215: signal is true;
	signal I12216: std_logic; attribute dont_touch of I12216: signal is true;
	signal I12223: std_logic; attribute dont_touch of I12223: signal is true;
	signal I12226: std_logic; attribute dont_touch of I12226: signal is true;
	signal I12229: std_logic; attribute dont_touch of I12229: signal is true;
	signal I12232: std_logic; attribute dont_touch of I12232: signal is true;
	signal I12235: std_logic; attribute dont_touch of I12235: signal is true;
	signal I12239: std_logic; attribute dont_touch of I12239: signal is true;
	signal I12242: std_logic; attribute dont_touch of I12242: signal is true;
	signal I12245: std_logic; attribute dont_touch of I12245: signal is true;
	signal I12248: std_logic; attribute dont_touch of I12248: signal is true;
	signal I12251: std_logic; attribute dont_touch of I12251: signal is true;
	signal I12255: std_logic; attribute dont_touch of I12255: signal is true;
	signal I12258: std_logic; attribute dont_touch of I12258: signal is true;
	signal I12261: std_logic; attribute dont_touch of I12261: signal is true;
	signal I12265: std_logic; attribute dont_touch of I12265: signal is true;
	signal I12268: std_logic; attribute dont_touch of I12268: signal is true;
	signal I12271: std_logic; attribute dont_touch of I12271: signal is true;
	signal I12274: std_logic; attribute dont_touch of I12274: signal is true;
	signal I12279: std_logic; attribute dont_touch of I12279: signal is true;
	signal I12282: std_logic; attribute dont_touch of I12282: signal is true;
	signal I12286: std_logic; attribute dont_touch of I12286: signal is true;
	signal I12289: std_logic; attribute dont_touch of I12289: signal is true;
	signal I12293: std_logic; attribute dont_touch of I12293: signal is true;
	signal I12296: std_logic; attribute dont_touch of I12296: signal is true;
	signal I12300: std_logic; attribute dont_touch of I12300: signal is true;
	signal I12303: std_logic; attribute dont_touch of I12303: signal is true;
	signal I12307: std_logic; attribute dont_touch of I12307: signal is true;
	signal I12318: std_logic; attribute dont_touch of I12318: signal is true;
	signal I12322: std_logic; attribute dont_touch of I12322: signal is true;
	signal I12326: std_logic; attribute dont_touch of I12326: signal is true;
	signal I12335: std_logic; attribute dont_touch of I12335: signal is true;
	signal I12339: std_logic; attribute dont_touch of I12339: signal is true;
	signal I12344: std_logic; attribute dont_touch of I12344: signal is true;
	signal I12354: std_logic; attribute dont_touch of I12354: signal is true;
	signal I12357: std_logic; attribute dont_touch of I12357: signal is true;
	signal I12360: std_logic; attribute dont_touch of I12360: signal is true;
	signal I12363: std_logic; attribute dont_touch of I12363: signal is true;
	signal I12366: std_logic; attribute dont_touch of I12366: signal is true;
	signal I12369: std_logic; attribute dont_touch of I12369: signal is true;
	signal I12372: std_logic; attribute dont_touch of I12372: signal is true;
	signal I12376: std_logic; attribute dont_touch of I12376: signal is true;
	signal I12380: std_logic; attribute dont_touch of I12380: signal is true;
	signal I12384: std_logic; attribute dont_touch of I12384: signal is true;
	signal I12388: std_logic; attribute dont_touch of I12388: signal is true;
	signal I12397: std_logic; attribute dont_touch of I12397: signal is true;
	signal I12400: std_logic; attribute dont_touch of I12400: signal is true;
	signal I12403: std_logic; attribute dont_touch of I12403: signal is true;
	signal I12406: std_logic; attribute dont_touch of I12406: signal is true;
	signal I12409: std_logic; attribute dont_touch of I12409: signal is true;
	signal I12412: std_logic; attribute dont_touch of I12412: signal is true;
	signal I12415: std_logic; attribute dont_touch of I12415: signal is true;
	signal I12418: std_logic; attribute dont_touch of I12418: signal is true;
	signal I12421: std_logic; attribute dont_touch of I12421: signal is true;
	signal I12424: std_logic; attribute dont_touch of I12424: signal is true;
	signal I12427: std_logic; attribute dont_touch of I12427: signal is true;
	signal I12430: std_logic; attribute dont_touch of I12430: signal is true;
	signal I12433: std_logic; attribute dont_touch of I12433: signal is true;
	signal I12436: std_logic; attribute dont_touch of I12436: signal is true;
	signal I12439: std_logic; attribute dont_touch of I12439: signal is true;
	signal I12442: std_logic; attribute dont_touch of I12442: signal is true;
	signal I12445: std_logic; attribute dont_touch of I12445: signal is true;
	signal I12448: std_logic; attribute dont_touch of I12448: signal is true;
	signal I12451: std_logic; attribute dont_touch of I12451: signal is true;
	signal I12454: std_logic; attribute dont_touch of I12454: signal is true;
	signal I12457: std_logic; attribute dont_touch of I12457: signal is true;
	signal I12460: std_logic; attribute dont_touch of I12460: signal is true;
	signal I12463: std_logic; attribute dont_touch of I12463: signal is true;
	signal I12466: std_logic; attribute dont_touch of I12466: signal is true;
	signal I12469: std_logic; attribute dont_touch of I12469: signal is true;
	signal I12472: std_logic; attribute dont_touch of I12472: signal is true;
	signal I12475: std_logic; attribute dont_touch of I12475: signal is true;
	signal I12478: std_logic; attribute dont_touch of I12478: signal is true;
	signal I12481: std_logic; attribute dont_touch of I12481: signal is true;
	signal I12484: std_logic; attribute dont_touch of I12484: signal is true;
	signal I12487: std_logic; attribute dont_touch of I12487: signal is true;
	signal I12490: std_logic; attribute dont_touch of I12490: signal is true;
	signal I12493: std_logic; attribute dont_touch of I12493: signal is true;
	signal I12496: std_logic; attribute dont_touch of I12496: signal is true;
	signal I12499: std_logic; attribute dont_touch of I12499: signal is true;
	signal I12502: std_logic; attribute dont_touch of I12502: signal is true;
	signal I12505: std_logic; attribute dont_touch of I12505: signal is true;
	signal I12508: std_logic; attribute dont_touch of I12508: signal is true;
	signal I12511: std_logic; attribute dont_touch of I12511: signal is true;
	signal I12514: std_logic; attribute dont_touch of I12514: signal is true;
	signal I12517: std_logic; attribute dont_touch of I12517: signal is true;
	signal I12520: std_logic; attribute dont_touch of I12520: signal is true;
	signal I12523: std_logic; attribute dont_touch of I12523: signal is true;
	signal I12526: std_logic; attribute dont_touch of I12526: signal is true;
	signal I12529: std_logic; attribute dont_touch of I12529: signal is true;
	signal I12532: std_logic; attribute dont_touch of I12532: signal is true;
	signal I12535: std_logic; attribute dont_touch of I12535: signal is true;
	signal I12538: std_logic; attribute dont_touch of I12538: signal is true;
	signal I12541: std_logic; attribute dont_touch of I12541: signal is true;
	signal I12544: std_logic; attribute dont_touch of I12544: signal is true;
	signal I12547: std_logic; attribute dont_touch of I12547: signal is true;
	signal I12550: std_logic; attribute dont_touch of I12550: signal is true;
	signal I12553: std_logic; attribute dont_touch of I12553: signal is true;
	signal I12556: std_logic; attribute dont_touch of I12556: signal is true;
	signal I12559: std_logic; attribute dont_touch of I12559: signal is true;
	signal I12562: std_logic; attribute dont_touch of I12562: signal is true;
	signal I12565: std_logic; attribute dont_touch of I12565: signal is true;
	signal I12568: std_logic; attribute dont_touch of I12568: signal is true;
	signal I12571: std_logic; attribute dont_touch of I12571: signal is true;
	signal I12574: std_logic; attribute dont_touch of I12574: signal is true;
	signal I12577: std_logic; attribute dont_touch of I12577: signal is true;
	signal I12580: std_logic; attribute dont_touch of I12580: signal is true;
	signal I12583: std_logic; attribute dont_touch of I12583: signal is true;
	signal I12586: std_logic; attribute dont_touch of I12586: signal is true;
	signal I12589: std_logic; attribute dont_touch of I12589: signal is true;
	signal I12592: std_logic; attribute dont_touch of I12592: signal is true;
	signal I12595: std_logic; attribute dont_touch of I12595: signal is true;
	signal I12598: std_logic; attribute dont_touch of I12598: signal is true;
	signal I12601: std_logic; attribute dont_touch of I12601: signal is true;
	signal I12604: std_logic; attribute dont_touch of I12604: signal is true;
	signal I12607: std_logic; attribute dont_touch of I12607: signal is true;
	signal I12610: std_logic; attribute dont_touch of I12610: signal is true;
	signal I12613: std_logic; attribute dont_touch of I12613: signal is true;
	signal I12616: std_logic; attribute dont_touch of I12616: signal is true;
	signal I12627: std_logic; attribute dont_touch of I12627: signal is true;
	signal I12631: std_logic; attribute dont_touch of I12631: signal is true;
	signal I12634: std_logic; attribute dont_touch of I12634: signal is true;
	signal I12638: std_logic; attribute dont_touch of I12638: signal is true;
	signal I12641: std_logic; attribute dont_touch of I12641: signal is true;
	signal I12644: std_logic; attribute dont_touch of I12644: signal is true;
	signal I12647: std_logic; attribute dont_touch of I12647: signal is true;
	signal I12652: std_logic; attribute dont_touch of I12652: signal is true;
	signal I12655: std_logic; attribute dont_touch of I12655: signal is true;
	signal I12678: std_logic; attribute dont_touch of I12678: signal is true;
	signal I12683: std_logic; attribute dont_touch of I12683: signal is true;
	signal I12690: std_logic; attribute dont_touch of I12690: signal is true;
	signal I12694: std_logic; attribute dont_touch of I12694: signal is true;
	signal I12712: std_logic; attribute dont_touch of I12712: signal is true;
	signal I12751: std_logic; attribute dont_touch of I12751: signal is true;
	signal I12759: std_logic; attribute dont_touch of I12759: signal is true;
	signal I12762: std_logic; attribute dont_touch of I12762: signal is true;
	signal I12765: std_logic; attribute dont_touch of I12765: signal is true;
	signal I12770: std_logic; attribute dont_touch of I12770: signal is true;
	signal I12773: std_logic; attribute dont_touch of I12773: signal is true;
	signal I12776: std_logic; attribute dont_touch of I12776: signal is true;
	signal I12779: std_logic; attribute dont_touch of I12779: signal is true;
	signal I12783: std_logic; attribute dont_touch of I12783: signal is true;
	signal I12786: std_logic; attribute dont_touch of I12786: signal is true;
	signal I12790: std_logic; attribute dont_touch of I12790: signal is true;
	signal I12793: std_logic; attribute dont_touch of I12793: signal is true;
	signal I12796: std_logic; attribute dont_touch of I12796: signal is true;
	signal I12799: std_logic; attribute dont_touch of I12799: signal is true;
	signal I12805: std_logic; attribute dont_touch of I12805: signal is true;
	signal I12809: std_logic; attribute dont_touch of I12809: signal is true;
	signal I12813: std_logic; attribute dont_touch of I12813: signal is true;
	signal I12817: std_logic; attribute dont_touch of I12817: signal is true;
	signal I12822: std_logic; attribute dont_touch of I12822: signal is true;
	signal I12825: std_logic; attribute dont_touch of I12825: signal is true;
	signal I12829: std_logic; attribute dont_touch of I12829: signal is true;
	signal I12832: std_logic; attribute dont_touch of I12832: signal is true;
	signal I12835: std_logic; attribute dont_touch of I12835: signal is true;
	signal I12838: std_logic; attribute dont_touch of I12838: signal is true;
	signal I12843: std_logic; attribute dont_touch of I12843: signal is true;
	signal I12846: std_logic; attribute dont_touch of I12846: signal is true;
	signal I12849: std_logic; attribute dont_touch of I12849: signal is true;
	signal I12853: std_logic; attribute dont_touch of I12853: signal is true;
	signal I12857: std_logic; attribute dont_touch of I12857: signal is true;
	signal I12862: std_logic; attribute dont_touch of I12862: signal is true;
	signal I12867: std_logic; attribute dont_touch of I12867: signal is true;
	signal I12871: std_logic; attribute dont_touch of I12871: signal is true;
	signal I12875: std_logic; attribute dont_touch of I12875: signal is true;
	signal I12878: std_logic; attribute dont_touch of I12878: signal is true;
	signal I12901: std_logic; attribute dont_touch of I12901: signal is true;
	signal I12904: std_logic; attribute dont_touch of I12904: signal is true;
	signal I12907: std_logic; attribute dont_touch of I12907: signal is true;
	signal I12910: std_logic; attribute dont_touch of I12910: signal is true;
	signal I12913: std_logic; attribute dont_touch of I12913: signal is true;
	signal I12916: std_logic; attribute dont_touch of I12916: signal is true;
	signal I12919: std_logic; attribute dont_touch of I12919: signal is true;
	signal I12930: std_logic; attribute dont_touch of I12930: signal is true;
	signal I12933: std_logic; attribute dont_touch of I12933: signal is true;
	signal I12936: std_logic; attribute dont_touch of I12936: signal is true;
	signal I12939: std_logic; attribute dont_touch of I12939: signal is true;
	signal I12942: std_logic; attribute dont_touch of I12942: signal is true;
	signal I12948: std_logic; attribute dont_touch of I12948: signal is true;
	signal I12953: std_logic; attribute dont_touch of I12953: signal is true;
	signal I12971: std_logic; attribute dont_touch of I12971: signal is true;
	signal I12978: std_logic; attribute dont_touch of I12978: signal is true;
	signal I12981: std_logic; attribute dont_touch of I12981: signal is true;
	signal I12986: std_logic; attribute dont_touch of I12986: signal is true;
	signal I12989: std_logic; attribute dont_touch of I12989: signal is true;
	signal I12993: std_logic; attribute dont_touch of I12993: signal is true;
	signal I12999: std_logic; attribute dont_touch of I12999: signal is true;
	signal I13002: std_logic; attribute dont_touch of I13002: signal is true;
	signal I13005: std_logic; attribute dont_touch of I13005: signal is true;
	signal I13010: std_logic; attribute dont_touch of I13010: signal is true;
	signal I13013: std_logic; attribute dont_touch of I13013: signal is true;
	signal I13017: std_logic; attribute dont_touch of I13017: signal is true;
	signal I13020: std_logic; attribute dont_touch of I13020: signal is true;
	signal I13023: std_logic; attribute dont_touch of I13023: signal is true;
	signal I13027: std_logic; attribute dont_touch of I13027: signal is true;
	signal I13030: std_logic; attribute dont_touch of I13030: signal is true;
	signal I13036: std_logic; attribute dont_touch of I13036: signal is true;
	signal I13039: std_logic; attribute dont_touch of I13039: signal is true;
	signal I13043: std_logic; attribute dont_touch of I13043: signal is true;
	signal I13048: std_logic; attribute dont_touch of I13048: signal is true;
	signal I13051: std_logic; attribute dont_touch of I13051: signal is true;
	signal I13057: std_logic; attribute dont_touch of I13057: signal is true;
	signal I13068: std_logic; attribute dont_touch of I13068: signal is true;
	signal I13076: std_logic; attribute dont_touch of I13076: signal is true;
	signal I13077: std_logic; attribute dont_touch of I13077: signal is true;
	signal I13078: std_logic; attribute dont_touch of I13078: signal is true;
	signal I13083: std_logic; attribute dont_touch of I13083: signal is true;
	signal I13086: std_logic; attribute dont_touch of I13086: signal is true;
	signal I13089: std_logic; attribute dont_touch of I13089: signal is true;
	signal I13090: std_logic; attribute dont_touch of I13090: signal is true;
	signal I13091: std_logic; attribute dont_touch of I13091: signal is true;
	signal I13096: std_logic; attribute dont_touch of I13096: signal is true;
	signal I13099: std_logic; attribute dont_touch of I13099: signal is true;
	signal I13102: std_logic; attribute dont_touch of I13102: signal is true;
	signal I13105: std_logic; attribute dont_touch of I13105: signal is true;
	signal I13109: std_logic; attribute dont_touch of I13109: signal is true;
	signal I13114: std_logic; attribute dont_touch of I13114: signal is true;
	signal I13117: std_logic; attribute dont_touch of I13117: signal is true;
	signal I13122: std_logic; attribute dont_touch of I13122: signal is true;
	signal I13125: std_logic; attribute dont_touch of I13125: signal is true;
	signal I13128: std_logic; attribute dont_touch of I13128: signal is true;
	signal I13131: std_logic; attribute dont_touch of I13131: signal is true;
	signal I13166: std_logic; attribute dont_touch of I13166: signal is true;
	signal I13185: std_logic; attribute dont_touch of I13185: signal is true;
	signal I13188: std_logic; attribute dont_touch of I13188: signal is true;
	signal I13191: std_logic; attribute dont_touch of I13191: signal is true;
	signal I13194: std_logic; attribute dont_touch of I13194: signal is true;
	signal I13197: std_logic; attribute dont_touch of I13197: signal is true;
	signal I13200: std_logic; attribute dont_touch of I13200: signal is true;
	signal I13203: std_logic; attribute dont_touch of I13203: signal is true;
	signal I13206: std_logic; attribute dont_touch of I13206: signal is true;
	signal I13209: std_logic; attribute dont_touch of I13209: signal is true;
	signal I13212: std_logic; attribute dont_touch of I13212: signal is true;
	signal I13224: std_logic; attribute dont_touch of I13224: signal is true;
	signal I13227: std_logic; attribute dont_touch of I13227: signal is true;
	signal I13230: std_logic; attribute dont_touch of I13230: signal is true;
	signal I13233: std_logic; attribute dont_touch of I13233: signal is true;
	signal I13236: std_logic; attribute dont_touch of I13236: signal is true;
	signal I13239: std_logic; attribute dont_touch of I13239: signal is true;
	signal I13242: std_logic; attribute dont_touch of I13242: signal is true;
	signal I13245: std_logic; attribute dont_touch of I13245: signal is true;
	signal I13248: std_logic; attribute dont_touch of I13248: signal is true;
	signal I13249: std_logic; attribute dont_touch of I13249: signal is true;
	signal I13250: std_logic; attribute dont_touch of I13250: signal is true;
	signal I13255: std_logic; attribute dont_touch of I13255: signal is true;
	signal I13258: std_logic; attribute dont_touch of I13258: signal is true;
	signal I13259: std_logic; attribute dont_touch of I13259: signal is true;
	signal I13260: std_logic; attribute dont_touch of I13260: signal is true;
	signal I13265: std_logic; attribute dont_touch of I13265: signal is true;
	signal I13266: std_logic; attribute dont_touch of I13266: signal is true;
	signal I13267: std_logic; attribute dont_touch of I13267: signal is true;
	signal I13272: std_logic; attribute dont_touch of I13272: signal is true;
	signal I13273: std_logic; attribute dont_touch of I13273: signal is true;
	signal I13274: std_logic; attribute dont_touch of I13274: signal is true;
	signal I13280: std_logic; attribute dont_touch of I13280: signal is true;
	signal I13283: std_logic; attribute dont_touch of I13283: signal is true;
	signal I13284: std_logic; attribute dont_touch of I13284: signal is true;
	signal I13285: std_logic; attribute dont_touch of I13285: signal is true;
	signal I13290: std_logic; attribute dont_touch of I13290: signal is true;
	signal I13293: std_logic; attribute dont_touch of I13293: signal is true;
	signal I13294: std_logic; attribute dont_touch of I13294: signal is true;
	signal I13295: std_logic; attribute dont_touch of I13295: signal is true;
	signal I13300: std_logic; attribute dont_touch of I13300: signal is true;
	signal I13301: std_logic; attribute dont_touch of I13301: signal is true;
	signal I13302: std_logic; attribute dont_touch of I13302: signal is true;
	signal I13307: std_logic; attribute dont_touch of I13307: signal is true;
	signal I13308: std_logic; attribute dont_touch of I13308: signal is true;
	signal I13309: std_logic; attribute dont_touch of I13309: signal is true;
	signal I13314: std_logic; attribute dont_touch of I13314: signal is true;
	signal I13317: std_logic; attribute dont_touch of I13317: signal is true;
	signal I13320: std_logic; attribute dont_touch of I13320: signal is true;
	signal I13323: std_logic; attribute dont_touch of I13323: signal is true;
	signal I13326: std_logic; attribute dont_touch of I13326: signal is true;
	signal I13329: std_logic; attribute dont_touch of I13329: signal is true;
	signal I13332: std_logic; attribute dont_touch of I13332: signal is true;
	signal I13335: std_logic; attribute dont_touch of I13335: signal is true;
	signal I13338: std_logic; attribute dont_touch of I13338: signal is true;
	signal I13341: std_logic; attribute dont_touch of I13341: signal is true;
	signal I13344: std_logic; attribute dont_touch of I13344: signal is true;
	signal I13347: std_logic; attribute dont_touch of I13347: signal is true;
	signal I13351: std_logic; attribute dont_touch of I13351: signal is true;
	signal I13354: std_logic; attribute dont_touch of I13354: signal is true;
	signal I13357: std_logic; attribute dont_touch of I13357: signal is true;
	signal I13360: std_logic; attribute dont_touch of I13360: signal is true;
	signal I13364: std_logic; attribute dont_touch of I13364: signal is true;
	signal I13367: std_logic; attribute dont_touch of I13367: signal is true;
	signal I13370: std_logic; attribute dont_touch of I13370: signal is true;
	signal I13373: std_logic; attribute dont_touch of I13373: signal is true;
	signal I13376: std_logic; attribute dont_touch of I13376: signal is true;
	signal I13379: std_logic; attribute dont_touch of I13379: signal is true;
	signal I13382: std_logic; attribute dont_touch of I13382: signal is true;
	signal I13385: std_logic; attribute dont_touch of I13385: signal is true;
	signal I13388: std_logic; attribute dont_touch of I13388: signal is true;
	signal I13391: std_logic; attribute dont_touch of I13391: signal is true;
	signal I13394: std_logic; attribute dont_touch of I13394: signal is true;
	signal I13397: std_logic; attribute dont_touch of I13397: signal is true;
	signal I13400: std_logic; attribute dont_touch of I13400: signal is true;
	signal I13403: std_logic; attribute dont_touch of I13403: signal is true;
	signal I13406: std_logic; attribute dont_touch of I13406: signal is true;
	signal I13409: std_logic; attribute dont_touch of I13409: signal is true;
	signal I13412: std_logic; attribute dont_touch of I13412: signal is true;
	signal I13415: std_logic; attribute dont_touch of I13415: signal is true;
	signal I13418: std_logic; attribute dont_touch of I13418: signal is true;
	signal I13421: std_logic; attribute dont_touch of I13421: signal is true;
	signal I13424: std_logic; attribute dont_touch of I13424: signal is true;
	signal I13427: std_logic; attribute dont_touch of I13427: signal is true;
	signal I13430: std_logic; attribute dont_touch of I13430: signal is true;
	signal I13433: std_logic; attribute dont_touch of I13433: signal is true;
	signal I13436: std_logic; attribute dont_touch of I13436: signal is true;
	signal I13439: std_logic; attribute dont_touch of I13439: signal is true;
	signal I13442: std_logic; attribute dont_touch of I13442: signal is true;
	signal I13445: std_logic; attribute dont_touch of I13445: signal is true;
	signal I13448: std_logic; attribute dont_touch of I13448: signal is true;
	signal I13451: std_logic; attribute dont_touch of I13451: signal is true;
	signal I13454: std_logic; attribute dont_touch of I13454: signal is true;
	signal I13457: std_logic; attribute dont_touch of I13457: signal is true;
	signal I13460: std_logic; attribute dont_touch of I13460: signal is true;
	signal I13463: std_logic; attribute dont_touch of I13463: signal is true;
	signal I13466: std_logic; attribute dont_touch of I13466: signal is true;
	signal I13469: std_logic; attribute dont_touch of I13469: signal is true;
	signal I13475: std_logic; attribute dont_touch of I13475: signal is true;
	signal I13478: std_logic; attribute dont_touch of I13478: signal is true;
	signal I13482: std_logic; attribute dont_touch of I13482: signal is true;
	signal I13485: std_logic; attribute dont_touch of I13485: signal is true;
	signal I13489: std_logic; attribute dont_touch of I13489: signal is true;
	signal I13504: std_logic; attribute dont_touch of I13504: signal is true;
	signal I13505: std_logic; attribute dont_touch of I13505: signal is true;
	signal I13506: std_logic; attribute dont_touch of I13506: signal is true;
	signal I13513: std_logic; attribute dont_touch of I13513: signal is true;
	signal I13514: std_logic; attribute dont_touch of I13514: signal is true;
	signal I13515: std_logic; attribute dont_touch of I13515: signal is true;
	signal I13521: std_logic; attribute dont_touch of I13521: signal is true;
	signal I13522: std_logic; attribute dont_touch of I13522: signal is true;
	signal I13523: std_logic; attribute dont_touch of I13523: signal is true;
	signal I13529: std_logic; attribute dont_touch of I13529: signal is true;
	signal I13530: std_logic; attribute dont_touch of I13530: signal is true;
	signal I13531: std_logic; attribute dont_touch of I13531: signal is true;
	signal I13537: std_logic; attribute dont_touch of I13537: signal is true;
	signal I13538: std_logic; attribute dont_touch of I13538: signal is true;
	signal I13539: std_logic; attribute dont_touch of I13539: signal is true;
	signal I13544: std_logic; attribute dont_touch of I13544: signal is true;
	signal I13545: std_logic; attribute dont_touch of I13545: signal is true;
	signal I13546: std_logic; attribute dont_touch of I13546: signal is true;
	signal I13552: std_logic; attribute dont_touch of I13552: signal is true;
	signal I13553: std_logic; attribute dont_touch of I13553: signal is true;
	signal I13554: std_logic; attribute dont_touch of I13554: signal is true;
	signal I13559: std_logic; attribute dont_touch of I13559: signal is true;
	signal I13560: std_logic; attribute dont_touch of I13560: signal is true;
	signal I13561: std_logic; attribute dont_touch of I13561: signal is true;
	signal I13568: std_logic; attribute dont_touch of I13568: signal is true;
	signal I13571: std_logic; attribute dont_touch of I13571: signal is true;
	signal I13574: std_logic; attribute dont_touch of I13574: signal is true;
	signal I13577: std_logic; attribute dont_touch of I13577: signal is true;
	signal I13580: std_logic; attribute dont_touch of I13580: signal is true;
	signal I13583: std_logic; attribute dont_touch of I13583: signal is true;
	signal I13586: std_logic; attribute dont_touch of I13586: signal is true;
	signal I13589: std_logic; attribute dont_touch of I13589: signal is true;
	signal I13592: std_logic; attribute dont_touch of I13592: signal is true;
	signal I13595: std_logic; attribute dont_touch of I13595: signal is true;
	signal I13606: std_logic; attribute dont_touch of I13606: signal is true;
	signal I13609: std_logic; attribute dont_touch of I13609: signal is true;
	signal I13612: std_logic; attribute dont_touch of I13612: signal is true;
	signal I13615: std_logic; attribute dont_touch of I13615: signal is true;
	signal I13618: std_logic; attribute dont_touch of I13618: signal is true;
	signal I13621: std_logic; attribute dont_touch of I13621: signal is true;
	signal I13624: std_logic; attribute dont_touch of I13624: signal is true;
	signal I13627: std_logic; attribute dont_touch of I13627: signal is true;
	signal I13630: std_logic; attribute dont_touch of I13630: signal is true;
	signal I13633: std_logic; attribute dont_touch of I13633: signal is true;
	signal I13636: std_logic; attribute dont_touch of I13636: signal is true;
	signal I13639: std_logic; attribute dont_touch of I13639: signal is true;
	signal I13642: std_logic; attribute dont_touch of I13642: signal is true;
	signal I13645: std_logic; attribute dont_touch of I13645: signal is true;
	signal I13648: std_logic; attribute dont_touch of I13648: signal is true;
	signal I13659: std_logic; attribute dont_touch of I13659: signal is true;
	signal I13660: std_logic; attribute dont_touch of I13660: signal is true;
	signal I13661: std_logic; attribute dont_touch of I13661: signal is true;
	signal I13666: std_logic; attribute dont_touch of I13666: signal is true;
	signal I13669: std_logic; attribute dont_touch of I13669: signal is true;
	signal I13674: std_logic; attribute dont_touch of I13674: signal is true;
	signal I13678: std_logic; attribute dont_touch of I13678: signal is true;
	signal I13682: std_logic; attribute dont_touch of I13682: signal is true;
	signal I13695: std_logic; attribute dont_touch of I13695: signal is true;
	signal I13708: std_logic; attribute dont_touch of I13708: signal is true;
	signal I13711: std_logic; attribute dont_touch of I13711: signal is true;
	signal I13714: std_logic; attribute dont_touch of I13714: signal is true;
	signal I13717: std_logic; attribute dont_touch of I13717: signal is true;
	signal I13720: std_logic; attribute dont_touch of I13720: signal is true;
	signal I13723: std_logic; attribute dont_touch of I13723: signal is true;
	signal I13726: std_logic; attribute dont_touch of I13726: signal is true;
	signal I13729: std_logic; attribute dont_touch of I13729: signal is true;
	signal I13732: std_logic; attribute dont_touch of I13732: signal is true;
	signal I13735: std_logic; attribute dont_touch of I13735: signal is true;
	signal I13738: std_logic; attribute dont_touch of I13738: signal is true;
	signal I13741: std_logic; attribute dont_touch of I13741: signal is true;
	signal I13744: std_logic; attribute dont_touch of I13744: signal is true;
	signal I13747: std_logic; attribute dont_touch of I13747: signal is true;
	signal I13765: std_logic; attribute dont_touch of I13765: signal is true;
	signal I13766: std_logic; attribute dont_touch of I13766: signal is true;
	signal I13767: std_logic; attribute dont_touch of I13767: signal is true;
	signal I13773: std_logic; attribute dont_touch of I13773: signal is true;
	signal I13776: std_logic; attribute dont_touch of I13776: signal is true;
	signal I13779: std_logic; attribute dont_touch of I13779: signal is true;
	signal I13782: std_logic; attribute dont_touch of I13782: signal is true;
	signal I13785: std_logic; attribute dont_touch of I13785: signal is true;
	signal I13788: std_logic; attribute dont_touch of I13788: signal is true;
	signal I13791: std_logic; attribute dont_touch of I13791: signal is true;
	signal I13794: std_logic; attribute dont_touch of I13794: signal is true;
	signal I13797: std_logic; attribute dont_touch of I13797: signal is true;
	signal I13800: std_logic; attribute dont_touch of I13800: signal is true;
	signal I13803: std_logic; attribute dont_touch of I13803: signal is true;
	signal I13806: std_logic; attribute dont_touch of I13806: signal is true;
	signal I13809: std_logic; attribute dont_touch of I13809: signal is true;
	signal I13812: std_logic; attribute dont_touch of I13812: signal is true;
	signal I13816: std_logic; attribute dont_touch of I13816: signal is true;
	signal I13819: std_logic; attribute dont_touch of I13819: signal is true;
	signal I13822: std_logic; attribute dont_touch of I13822: signal is true;
	signal I13825: std_logic; attribute dont_touch of I13825: signal is true;
	signal I13828: std_logic; attribute dont_touch of I13828: signal is true;
	signal I13831: std_logic; attribute dont_touch of I13831: signal is true;
	signal I13834: std_logic; attribute dont_touch of I13834: signal is true;
	signal I13837: std_logic; attribute dont_touch of I13837: signal is true;
	signal I13840: std_logic; attribute dont_touch of I13840: signal is true;
	signal I13857: std_logic; attribute dont_touch of I13857: signal is true;
	signal I13858: std_logic; attribute dont_touch of I13858: signal is true;
	signal I13859: std_logic; attribute dont_touch of I13859: signal is true;
	signal I13867: std_logic; attribute dont_touch of I13867: signal is true;
	signal I13868: std_logic; attribute dont_touch of I13868: signal is true;
	signal I13869: std_logic; attribute dont_touch of I13869: signal is true;
	signal I13876: std_logic; attribute dont_touch of I13876: signal is true;
	signal I13877: std_logic; attribute dont_touch of I13877: signal is true;
	signal I13878: std_logic; attribute dont_touch of I13878: signal is true;
	signal I13886: std_logic; attribute dont_touch of I13886: signal is true;
	signal I13887: std_logic; attribute dont_touch of I13887: signal is true;
	signal I13888: std_logic; attribute dont_touch of I13888: signal is true;
	signal I13893: std_logic; attribute dont_touch of I13893: signal is true;
	signal I13894: std_logic; attribute dont_touch of I13894: signal is true;
	signal I13895: std_logic; attribute dont_touch of I13895: signal is true;
	signal I13900: std_logic; attribute dont_touch of I13900: signal is true;
	signal I13901: std_logic; attribute dont_touch of I13901: signal is true;
	signal I13902: std_logic; attribute dont_touch of I13902: signal is true;
	signal I13907: std_logic; attribute dont_touch of I13907: signal is true;
	signal I13908: std_logic; attribute dont_touch of I13908: signal is true;
	signal I13909: std_logic; attribute dont_touch of I13909: signal is true;
	signal I13915: std_logic; attribute dont_touch of I13915: signal is true;
	signal I13918: std_logic; attribute dont_touch of I13918: signal is true;
	signal I13933: std_logic; attribute dont_touch of I13933: signal is true;
	signal I13941: std_logic; attribute dont_touch of I13941: signal is true;
	signal I13945: std_logic; attribute dont_touch of I13945: signal is true;
	signal I13949: std_logic; attribute dont_touch of I13949: signal is true;
	signal I13952: std_logic; attribute dont_touch of I13952: signal is true;
	signal I13956: std_logic; attribute dont_touch of I13956: signal is true;
	signal I13959: std_logic; attribute dont_touch of I13959: signal is true;
	signal I13962: std_logic; attribute dont_touch of I13962: signal is true;
	signal I13965: std_logic; attribute dont_touch of I13965: signal is true;
	signal I13969: std_logic; attribute dont_touch of I13969: signal is true;
	signal I13975: std_logic; attribute dont_touch of I13975: signal is true;
	signal I13978: std_logic; attribute dont_touch of I13978: signal is true;
	signal I13990: std_logic; attribute dont_touch of I13990: signal is true;
	signal I13991: std_logic; attribute dont_touch of I13991: signal is true;
	signal I13992: std_logic; attribute dont_touch of I13992: signal is true;
	signal I14005: std_logic; attribute dont_touch of I14005: signal is true;
	signal I14010: std_logic; attribute dont_touch of I14010: signal is true;
	signal I14040: std_logic; attribute dont_touch of I14040: signal is true;
	signal I14045: std_logic; attribute dont_touch of I14045: signal is true;
	signal I14055: std_logic; attribute dont_touch of I14055: signal is true;
	signal I14077: std_logic; attribute dont_touch of I14077: signal is true;
	signal I14080: std_logic; attribute dont_touch of I14080: signal is true;
	signal I14083: std_logic; attribute dont_touch of I14083: signal is true;
	signal I14087: std_logic; attribute dont_touch of I14087: signal is true;
	signal I14090: std_logic; attribute dont_touch of I14090: signal is true;
	signal I14094: std_logic; attribute dont_touch of I14094: signal is true;
	signal I14097: std_logic; attribute dont_touch of I14097: signal is true;
	signal I14101: std_logic; attribute dont_touch of I14101: signal is true;
	signal I14105: std_logic; attribute dont_touch of I14105: signal is true;
	signal I14109: std_logic; attribute dont_touch of I14109: signal is true;
	signal I14112: std_logic; attribute dont_touch of I14112: signal is true;
	signal I14116: std_logic; attribute dont_touch of I14116: signal is true;
	signal I14119: std_logic; attribute dont_touch of I14119: signal is true;
	signal I14123: std_logic; attribute dont_touch of I14123: signal is true;
	signal I14127: std_logic; attribute dont_touch of I14127: signal is true;
	signal I14130: std_logic; attribute dont_touch of I14130: signal is true;
	signal I14133: std_logic; attribute dont_touch of I14133: signal is true;
	signal I14136: std_logic; attribute dont_touch of I14136: signal is true;
	signal I14140: std_logic; attribute dont_touch of I14140: signal is true;
	signal I14176: std_logic; attribute dont_touch of I14176: signal is true;
	signal I14179: std_logic; attribute dont_touch of I14179: signal is true;
	signal I14182: std_logic; attribute dont_touch of I14182: signal is true;
	signal I14185: std_logic; attribute dont_touch of I14185: signal is true;
	signal I14188: std_logic; attribute dont_touch of I14188: signal is true;
	signal I14191: std_logic; attribute dont_touch of I14191: signal is true;
	signal I14194: std_logic; attribute dont_touch of I14194: signal is true;
	signal I14202: std_logic; attribute dont_touch of I14202: signal is true;
	signal I14203: std_logic; attribute dont_touch of I14203: signal is true;
	signal I14204: std_logic; attribute dont_touch of I14204: signal is true;
	signal I14209: std_logic; attribute dont_touch of I14209: signal is true;
	signal I14210: std_logic; attribute dont_touch of I14210: signal is true;
	signal I14211: std_logic; attribute dont_touch of I14211: signal is true;
	signal I14216: std_logic; attribute dont_touch of I14216: signal is true;
	signal I14217: std_logic; attribute dont_touch of I14217: signal is true;
	signal I14218: std_logic; attribute dont_touch of I14218: signal is true;
	signal I14224: std_logic; attribute dont_touch of I14224: signal is true;
	signal I14228: std_logic; attribute dont_touch of I14228: signal is true;
	signal I14232: std_logic; attribute dont_touch of I14232: signal is true;
	signal I14236: std_logic; attribute dont_touch of I14236: signal is true;
	signal I14239: std_logic; attribute dont_touch of I14239: signal is true;
	signal I14242: std_logic; attribute dont_touch of I14242: signal is true;
	signal I14249: std_logic; attribute dont_touch of I14249: signal is true;
	signal I14252: std_logic; attribute dont_touch of I14252: signal is true;
	signal I14257: std_logic; attribute dont_touch of I14257: signal is true;
	signal I14263: std_logic; attribute dont_touch of I14263: signal is true;
	signal I14264: std_logic; attribute dont_touch of I14264: signal is true;
	signal I14265: std_logic; attribute dont_touch of I14265: signal is true;
	signal I14270: std_logic; attribute dont_touch of I14270: signal is true;
	signal I14271: std_logic; attribute dont_touch of I14271: signal is true;
	signal I14272: std_logic; attribute dont_touch of I14272: signal is true;
	signal I14277: std_logic; attribute dont_touch of I14277: signal is true;
	signal I14278: std_logic; attribute dont_touch of I14278: signal is true;
	signal I14279: std_logic; attribute dont_touch of I14279: signal is true;
	signal I14295: std_logic; attribute dont_touch of I14295: signal is true;
	signal I14299: std_logic; attribute dont_touch of I14299: signal is true;
	signal I14303: std_logic; attribute dont_touch of I14303: signal is true;
	signal I14306: std_logic; attribute dont_touch of I14306: signal is true;
	signal I14309: std_logic; attribute dont_touch of I14309: signal is true;
	signal I14312: std_logic; attribute dont_touch of I14312: signal is true;
	signal I14315: std_logic; attribute dont_touch of I14315: signal is true;
	signal I14319: std_logic; attribute dont_touch of I14319: signal is true;
	signal I14323: std_logic; attribute dont_touch of I14323: signal is true;
	signal I14326: std_logic; attribute dont_touch of I14326: signal is true;
	signal I14330: std_logic; attribute dont_touch of I14330: signal is true;
	signal I14340: std_logic; attribute dont_touch of I14340: signal is true;
	signal I14349: std_logic; attribute dont_touch of I14349: signal is true;
	signal I14352: std_logic; attribute dont_touch of I14352: signal is true;
	signal I14355: std_logic; attribute dont_touch of I14355: signal is true;
	signal I14358: std_logic; attribute dont_touch of I14358: signal is true;
	signal I14361: std_logic; attribute dont_touch of I14361: signal is true;
	signal I14364: std_logic; attribute dont_touch of I14364: signal is true;
	signal I14367: std_logic; attribute dont_touch of I14367: signal is true;
	signal I14370: std_logic; attribute dont_touch of I14370: signal is true;
	signal I14373: std_logic; attribute dont_touch of I14373: signal is true;
	signal I14376: std_logic; attribute dont_touch of I14376: signal is true;
	signal I14379: std_logic; attribute dont_touch of I14379: signal is true;
	signal I14382: std_logic; attribute dont_touch of I14382: signal is true;
	signal I14385: std_logic; attribute dont_touch of I14385: signal is true;
	signal I14388: std_logic; attribute dont_touch of I14388: signal is true;
	signal I14391: std_logic; attribute dont_touch of I14391: signal is true;
	signal I14394: std_logic; attribute dont_touch of I14394: signal is true;
	signal I14397: std_logic; attribute dont_touch of I14397: signal is true;
	signal I14400: std_logic; attribute dont_touch of I14400: signal is true;
	signal I14405: std_logic; attribute dont_touch of I14405: signal is true;
	signal I14409: std_logic; attribute dont_touch of I14409: signal is true;
	signal I14412: std_logic; attribute dont_touch of I14412: signal is true;
	signal I14415: std_logic; attribute dont_touch of I14415: signal is true;
	signal I14418: std_logic; attribute dont_touch of I14418: signal is true;
	signal I14421: std_logic; attribute dont_touch of I14421: signal is true;
	signal I14424: std_logic; attribute dont_touch of I14424: signal is true;
	signal I14439: std_logic; attribute dont_touch of I14439: signal is true;
	signal I14442: std_logic; attribute dont_touch of I14442: signal is true;
	signal I14443: std_logic; attribute dont_touch of I14443: signal is true;
	signal I14444: std_logic; attribute dont_touch of I14444: signal is true;
	signal I14449: std_logic; attribute dont_touch of I14449: signal is true;
	signal I14452: std_logic; attribute dont_touch of I14452: signal is true;
	signal I14473: std_logic; attribute dont_touch of I14473: signal is true;
	signal I14477: std_logic; attribute dont_touch of I14477: signal is true;
	signal I14485: std_logic; attribute dont_touch of I14485: signal is true;
	signal I14490: std_logic; attribute dont_touch of I14490: signal is true;
	signal I14494: std_logic; attribute dont_touch of I14494: signal is true;
	signal I14499: std_logic; attribute dont_touch of I14499: signal is true;
	signal I14503: std_logic; attribute dont_touch of I14503: signal is true;
	signal I14506: std_logic; attribute dont_touch of I14506: signal is true;
	signal I14509: std_logic; attribute dont_touch of I14509: signal is true;
	signal I14519: std_logic; attribute dont_touch of I14519: signal is true;
	signal I14522: std_logic; attribute dont_touch of I14522: signal is true;
	signal I14525: std_logic; attribute dont_touch of I14525: signal is true;
	signal I14528: std_logic; attribute dont_touch of I14528: signal is true;
	signal I14531: std_logic; attribute dont_touch of I14531: signal is true;
	signal I14534: std_logic; attribute dont_touch of I14534: signal is true;
	signal I14537: std_logic; attribute dont_touch of I14537: signal is true;
	signal I14540: std_logic; attribute dont_touch of I14540: signal is true;
	signal I14543: std_logic; attribute dont_touch of I14543: signal is true;
	signal I14546: std_logic; attribute dont_touch of I14546: signal is true;
	signal I14549: std_logic; attribute dont_touch of I14549: signal is true;
	signal I14552: std_logic; attribute dont_touch of I14552: signal is true;
	signal I14555: std_logic; attribute dont_touch of I14555: signal is true;
	signal I14558: std_logic; attribute dont_touch of I14558: signal is true;
	signal I14561: std_logic; attribute dont_touch of I14561: signal is true;
	signal I14564: std_logic; attribute dont_touch of I14564: signal is true;
	signal I14567: std_logic; attribute dont_touch of I14567: signal is true;
	signal I14570: std_logic; attribute dont_touch of I14570: signal is true;
	signal I14573: std_logic; attribute dont_touch of I14573: signal is true;
	signal I14579: std_logic; attribute dont_touch of I14579: signal is true;
	signal I14582: std_logic; attribute dont_touch of I14582: signal is true;
	signal I14585: std_logic; attribute dont_touch of I14585: signal is true;
	signal I14596: std_logic; attribute dont_touch of I14596: signal is true;
	signal I14602: std_logic; attribute dont_touch of I14602: signal is true;
	signal I14607: std_logic; attribute dont_touch of I14607: signal is true;
	signal I14612: std_logic; attribute dont_touch of I14612: signal is true;
	signal I14613: std_logic; attribute dont_touch of I14613: signal is true;
	signal I14614: std_logic; attribute dont_touch of I14614: signal is true;
	signal I14642: std_logic; attribute dont_touch of I14642: signal is true;
	signal I14645: std_logic; attribute dont_touch of I14645: signal is true;
	signal I14668: std_logic; attribute dont_touch of I14668: signal is true;
	signal I14672: std_logic; attribute dont_touch of I14672: signal is true;
	signal I14675: std_logic; attribute dont_touch of I14675: signal is true;
	signal I14678: std_logic; attribute dont_touch of I14678: signal is true;
	signal I14681: std_logic; attribute dont_touch of I14681: signal is true;
	signal I14684: std_logic; attribute dont_touch of I14684: signal is true;
	signal I14687: std_logic; attribute dont_touch of I14687: signal is true;
	signal I14690: std_logic; attribute dont_touch of I14690: signal is true;
	signal I14694: std_logic; attribute dont_touch of I14694: signal is true;
	signal I14697: std_logic; attribute dont_touch of I14697: signal is true;
	signal I14701: std_logic; attribute dont_touch of I14701: signal is true;
	signal I14709: std_logic; attribute dont_touch of I14709: signal is true;
	signal I14713: std_logic; attribute dont_touch of I14713: signal is true;
	signal I14751: std_logic; attribute dont_touch of I14751: signal is true;
	signal I14776: std_logic; attribute dont_touch of I14776: signal is true;
	signal I14779: std_logic; attribute dont_touch of I14779: signal is true;
	signal I14786: std_logic; attribute dont_touch of I14786: signal is true;
	signal I14793: std_logic; attribute dont_touch of I14793: signal is true;
	signal I14799: std_logic; attribute dont_touch of I14799: signal is true;
	signal I14802: std_logic; attribute dont_touch of I14802: signal is true;
	signal I14805: std_logic; attribute dont_touch of I14805: signal is true;
	signal I14822: std_logic; attribute dont_touch of I14822: signal is true;
	signal I14827: std_logic; attribute dont_touch of I14827: signal is true;
	signal I14831: std_logic; attribute dont_touch of I14831: signal is true;
	signal I14835: std_logic; attribute dont_touch of I14835: signal is true;
	signal I14855: std_logic; attribute dont_touch of I14855: signal is true;
	signal I14858: std_logic; attribute dont_touch of I14858: signal is true;
	signal I14862: std_logic; attribute dont_touch of I14862: signal is true;
	signal I14866: std_logic; attribute dont_touch of I14866: signal is true;
	signal I14873: std_logic; attribute dont_touch of I14873: signal is true;
	signal I14876: std_logic; attribute dont_touch of I14876: signal is true;
	signal I14884: std_logic; attribute dont_touch of I14884: signal is true;
	signal I14888: std_logic; attribute dont_touch of I14888: signal is true;
	signal I14903: std_logic; attribute dont_touch of I14903: signal is true;
	signal I14906: std_logic; attribute dont_touch of I14906: signal is true;
	signal I14910: std_logic; attribute dont_touch of I14910: signal is true;
	signal I14914: std_logic; attribute dont_touch of I14914: signal is true;
	signal I14918: std_logic; attribute dont_touch of I14918: signal is true;
	signal I14933: std_logic; attribute dont_touch of I14933: signal is true;
	signal I14939: std_logic; attribute dont_touch of I14939: signal is true;
	signal I14944: std_logic; attribute dont_touch of I14944: signal is true;
	signal I14948: std_logic; attribute dont_touch of I14948: signal is true;
	signal I14955: std_logic; attribute dont_touch of I14955: signal is true;
	signal I14958: std_logic; attribute dont_touch of I14958: signal is true;
	signal I14961: std_logic; attribute dont_touch of I14961: signal is true;
	signal I14964: std_logic; attribute dont_touch of I14964: signal is true;
	signal I14967: std_logic; attribute dont_touch of I14967: signal is true;
	signal I14970: std_logic; attribute dont_touch of I14970: signal is true;
	signal I14973: std_logic; attribute dont_touch of I14973: signal is true;
	signal I14976: std_logic; attribute dont_touch of I14976: signal is true;
	signal I14979: std_logic; attribute dont_touch of I14979: signal is true;
	signal I14982: std_logic; attribute dont_touch of I14982: signal is true;
	signal I14989: std_logic; attribute dont_touch of I14989: signal is true;
	signal I15033: std_logic; attribute dont_touch of I15033: signal is true;
	signal I15036: std_logic; attribute dont_touch of I15036: signal is true;
	signal I15039: std_logic; attribute dont_touch of I15039: signal is true;
	signal I15042: std_logic; attribute dont_touch of I15042: signal is true;
	signal I15045: std_logic; attribute dont_touch of I15045: signal is true;
	signal I15048: std_logic; attribute dont_touch of I15048: signal is true;
	signal I15051: std_logic; attribute dont_touch of I15051: signal is true;
	signal I15054: std_logic; attribute dont_touch of I15054: signal is true;
	signal I15057: std_logic; attribute dont_touch of I15057: signal is true;
	signal I15060: std_logic; attribute dont_touch of I15060: signal is true;
	signal I15063: std_logic; attribute dont_touch of I15063: signal is true;
	signal I15068: std_logic; attribute dont_touch of I15068: signal is true;
	signal I15072: std_logic; attribute dont_touch of I15072: signal is true;
	signal I15075: std_logic; attribute dont_touch of I15075: signal is true;
	signal I15079: std_logic; attribute dont_touch of I15079: signal is true;
	signal I15082: std_logic; attribute dont_touch of I15082: signal is true;
	signal I15085: std_logic; attribute dont_touch of I15085: signal is true;
	signal I15088: std_logic; attribute dont_touch of I15088: signal is true;
	signal I15114: std_logic; attribute dont_touch of I15114: signal is true;
	signal I15127: std_logic; attribute dont_touch of I15127: signal is true;
	signal I15157: std_logic; attribute dont_touch of I15157: signal is true;
	signal I15162: std_logic; attribute dont_touch of I15162: signal is true;
	signal I15171: std_logic; attribute dont_touch of I15171: signal is true;
	signal I15172: std_logic; attribute dont_touch of I15172: signal is true;
	signal I15176: std_logic; attribute dont_touch of I15176: signal is true;
	signal I15177: std_logic; attribute dont_touch of I15177: signal is true;
	signal I15181: std_logic; attribute dont_touch of I15181: signal is true;
	signal I15184: std_logic; attribute dont_touch of I15184: signal is true;
	signal I15187: std_logic; attribute dont_touch of I15187: signal is true;
	signal I15190: std_logic; attribute dont_touch of I15190: signal is true;
	signal I15193: std_logic; attribute dont_touch of I15193: signal is true;
	signal I15196: std_logic; attribute dont_touch of I15196: signal is true;
	signal I15199: std_logic; attribute dont_touch of I15199: signal is true;
	signal I15200: std_logic; attribute dont_touch of I15200: signal is true;
	signal I15204: std_logic; attribute dont_touch of I15204: signal is true;
	signal I15205: std_logic; attribute dont_touch of I15205: signal is true;
	signal I15209: std_logic; attribute dont_touch of I15209: signal is true;
	signal I15210: std_logic; attribute dont_touch of I15210: signal is true;
	signal I15214: std_logic; attribute dont_touch of I15214: signal is true;
	signal I15215: std_logic; attribute dont_touch of I15215: signal is true;
	signal I15219: std_logic; attribute dont_touch of I15219: signal is true;
	signal I15220: std_logic; attribute dont_touch of I15220: signal is true;
	signal I15224: std_logic; attribute dont_touch of I15224: signal is true;
	signal I15225: std_logic; attribute dont_touch of I15225: signal is true;
	signal I15229: std_logic; attribute dont_touch of I15229: signal is true;
	signal I15232: std_logic; attribute dont_touch of I15232: signal is true;
	signal I15235: std_logic; attribute dont_touch of I15235: signal is true;
	signal I15238: std_logic; attribute dont_touch of I15238: signal is true;
	signal I15241: std_logic; attribute dont_touch of I15241: signal is true;
	signal I15244: std_logic; attribute dont_touch of I15244: signal is true;
	signal I15247: std_logic; attribute dont_touch of I15247: signal is true;
	signal I15250: std_logic; attribute dont_touch of I15250: signal is true;
	signal I15253: std_logic; attribute dont_touch of I15253: signal is true;
	signal I15256: std_logic; attribute dont_touch of I15256: signal is true;
	signal I15257: std_logic; attribute dont_touch of I15257: signal is true;
	signal I15258: std_logic; attribute dont_touch of I15258: signal is true;
	signal I15263: std_logic; attribute dont_touch of I15263: signal is true;
	signal I15266: std_logic; attribute dont_touch of I15266: signal is true;
	signal I15269: std_logic; attribute dont_touch of I15269: signal is true;
	signal I15272: std_logic; attribute dont_touch of I15272: signal is true;
	signal I15275: std_logic; attribute dont_touch of I15275: signal is true;
	signal I15278: std_logic; attribute dont_touch of I15278: signal is true;
	signal I15281: std_logic; attribute dont_touch of I15281: signal is true;
	signal I15284: std_logic; attribute dont_touch of I15284: signal is true;
	signal I15287: std_logic; attribute dont_touch of I15287: signal is true;
	signal I15290: std_logic; attribute dont_touch of I15290: signal is true;
	signal I15293: std_logic; attribute dont_touch of I15293: signal is true;
	signal I15296: std_logic; attribute dont_touch of I15296: signal is true;
	signal I15299: std_logic; attribute dont_touch of I15299: signal is true;
	signal I15302: std_logic; attribute dont_touch of I15302: signal is true;
	signal I15305: std_logic; attribute dont_touch of I15305: signal is true;
	signal I15308: std_logic; attribute dont_touch of I15308: signal is true;
	signal I15311: std_logic; attribute dont_touch of I15311: signal is true;
	signal I15314: std_logic; attribute dont_touch of I15314: signal is true;
	signal I15317: std_logic; attribute dont_touch of I15317: signal is true;
	signal I15320: std_logic; attribute dont_touch of I15320: signal is true;
	signal I15323: std_logic; attribute dont_touch of I15323: signal is true;
	signal I15326: std_logic; attribute dont_touch of I15326: signal is true;
	signal I15329: std_logic; attribute dont_touch of I15329: signal is true;
	signal I15332: std_logic; attribute dont_touch of I15332: signal is true;
	signal I15335: std_logic; attribute dont_touch of I15335: signal is true;
	signal I15338: std_logic; attribute dont_touch of I15338: signal is true;
	signal I15341: std_logic; attribute dont_touch of I15341: signal is true;
	signal I15344: std_logic; attribute dont_touch of I15344: signal is true;
	signal I15347: std_logic; attribute dont_touch of I15347: signal is true;
	signal I15350: std_logic; attribute dont_touch of I15350: signal is true;
	signal I15353: std_logic; attribute dont_touch of I15353: signal is true;
	signal I15356: std_logic; attribute dont_touch of I15356: signal is true;
	signal I15359: std_logic; attribute dont_touch of I15359: signal is true;
	signal I15362: std_logic; attribute dont_touch of I15362: signal is true;
	signal I15365: std_logic; attribute dont_touch of I15365: signal is true;
	signal I15368: std_logic; attribute dont_touch of I15368: signal is true;
	signal I15371: std_logic; attribute dont_touch of I15371: signal is true;
	signal I15374: std_logic; attribute dont_touch of I15374: signal is true;
	signal I15377: std_logic; attribute dont_touch of I15377: signal is true;
	signal I15380: std_logic; attribute dont_touch of I15380: signal is true;
	signal I15383: std_logic; attribute dont_touch of I15383: signal is true;
	signal I15386: std_logic; attribute dont_touch of I15386: signal is true;
	signal I15389: std_logic; attribute dont_touch of I15389: signal is true;
	signal I15392: std_logic; attribute dont_touch of I15392: signal is true;
	signal I15395: std_logic; attribute dont_touch of I15395: signal is true;
	signal I15400: std_logic; attribute dont_touch of I15400: signal is true;
	signal I15403: std_logic; attribute dont_touch of I15403: signal is true;
	signal I15406: std_logic; attribute dont_touch of I15406: signal is true;
	signal I15409: std_logic; attribute dont_touch of I15409: signal is true;
	signal I15412: std_logic; attribute dont_touch of I15412: signal is true;
	signal I15415: std_logic; attribute dont_touch of I15415: signal is true;
	signal I15418: std_logic; attribute dont_touch of I15418: signal is true;
	signal I15421: std_logic; attribute dont_touch of I15421: signal is true;
	signal I15424: std_logic; attribute dont_touch of I15424: signal is true;
	signal I15427: std_logic; attribute dont_touch of I15427: signal is true;
	signal I15430: std_logic; attribute dont_touch of I15430: signal is true;
	signal I15431: std_logic; attribute dont_touch of I15431: signal is true;
	signal I15432: std_logic; attribute dont_touch of I15432: signal is true;
	signal I15437: std_logic; attribute dont_touch of I15437: signal is true;
	signal I15441: std_logic; attribute dont_touch of I15441: signal is true;
	signal I15442: std_logic; attribute dont_touch of I15442: signal is true;
	signal I15443: std_logic; attribute dont_touch of I15443: signal is true;
	signal I15448: std_logic; attribute dont_touch of I15448: signal is true;
	signal I15451: std_logic; attribute dont_touch of I15451: signal is true;
	signal I15452: std_logic; attribute dont_touch of I15452: signal is true;
	signal I15453: std_logic; attribute dont_touch of I15453: signal is true;
	signal I15458: std_logic; attribute dont_touch of I15458: signal is true;
	signal I15461: std_logic; attribute dont_touch of I15461: signal is true;
	signal I15464: std_logic; attribute dont_touch of I15464: signal is true;
	signal I15467: std_logic; attribute dont_touch of I15467: signal is true;
	signal I15470: std_logic; attribute dont_touch of I15470: signal is true;
	signal I15473: std_logic; attribute dont_touch of I15473: signal is true;
	signal I15476: std_logic; attribute dont_touch of I15476: signal is true;
	signal I15479: std_logic; attribute dont_touch of I15479: signal is true;
	signal I15482: std_logic; attribute dont_touch of I15482: signal is true;
	signal I15485: std_logic; attribute dont_touch of I15485: signal is true;
	signal I15488: std_logic; attribute dont_touch of I15488: signal is true;
	signal I15491: std_logic; attribute dont_touch of I15491: signal is true;
	signal I15494: std_logic; attribute dont_touch of I15494: signal is true;
	signal I15497: std_logic; attribute dont_touch of I15497: signal is true;
	signal I15500: std_logic; attribute dont_touch of I15500: signal is true;
	signal I15503: std_logic; attribute dont_touch of I15503: signal is true;
	signal I15507: std_logic; attribute dont_touch of I15507: signal is true;
	signal I15510: std_logic; attribute dont_touch of I15510: signal is true;
	signal I15514: std_logic; attribute dont_touch of I15514: signal is true;
	signal I15517: std_logic; attribute dont_touch of I15517: signal is true;
	signal I15520: std_logic; attribute dont_touch of I15520: signal is true;
	signal I15523: std_logic; attribute dont_touch of I15523: signal is true;
	signal I15526: std_logic; attribute dont_touch of I15526: signal is true;
	signal I15530: std_logic; attribute dont_touch of I15530: signal is true;
	signal I15536: std_logic; attribute dont_touch of I15536: signal is true;
	signal I15539: std_logic; attribute dont_touch of I15539: signal is true;
	signal I15542: std_logic; attribute dont_touch of I15542: signal is true;
	signal I15545: std_logic; attribute dont_touch of I15545: signal is true;
	signal I15548: std_logic; attribute dont_touch of I15548: signal is true;
	signal I15551: std_logic; attribute dont_touch of I15551: signal is true;
	signal I15554: std_logic; attribute dont_touch of I15554: signal is true;
	signal I15559: std_logic; attribute dont_touch of I15559: signal is true;
	signal I15562: std_logic; attribute dont_touch of I15562: signal is true;
	signal I15565: std_logic; attribute dont_touch of I15565: signal is true;
	signal I15568: std_logic; attribute dont_touch of I15568: signal is true;
	signal I15580: std_logic; attribute dont_touch of I15580: signal is true;
	signal I15583: std_logic; attribute dont_touch of I15583: signal is true;
	signal I15586: std_logic; attribute dont_touch of I15586: signal is true;
	signal I15589: std_logic; attribute dont_touch of I15589: signal is true;
	signal I15592: std_logic; attribute dont_touch of I15592: signal is true;
	signal I15595: std_logic; attribute dont_touch of I15595: signal is true;
	signal I15598: std_logic; attribute dont_touch of I15598: signal is true;
	signal I15601: std_logic; attribute dont_touch of I15601: signal is true;
	signal I15604: std_logic; attribute dont_touch of I15604: signal is true;
	signal I15607: std_logic; attribute dont_touch of I15607: signal is true;
	signal I15608: std_logic; attribute dont_touch of I15608: signal is true;
	signal I15609: std_logic; attribute dont_touch of I15609: signal is true;
	signal I15615: std_logic; attribute dont_touch of I15615: signal is true;
	signal I15616: std_logic; attribute dont_touch of I15616: signal is true;
	signal I15617: std_logic; attribute dont_touch of I15617: signal is true;
	signal I15632: std_logic; attribute dont_touch of I15632: signal is true;
	signal I15635: std_logic; attribute dont_touch of I15635: signal is true;
	signal I15639: std_logic; attribute dont_touch of I15639: signal is true;
	signal I15665: std_logic; attribute dont_touch of I15665: signal is true;
	signal I15669: std_logic; attribute dont_touch of I15669: signal is true;
	signal I15672: std_logic; attribute dont_touch of I15672: signal is true;
	signal I15675: std_logic; attribute dont_touch of I15675: signal is true;
	signal I15688: std_logic; attribute dont_touch of I15688: signal is true;
	signal I15691: std_logic; attribute dont_touch of I15691: signal is true;
	signal I15694: std_logic; attribute dont_touch of I15694: signal is true;
	signal I15698: std_logic; attribute dont_touch of I15698: signal is true;
	signal I15701: std_logic; attribute dont_touch of I15701: signal is true;
	signal I15704: std_logic; attribute dont_touch of I15704: signal is true;
	signal I15708: std_logic; attribute dont_touch of I15708: signal is true;
	signal I15716: std_logic; attribute dont_touch of I15716: signal is true;
	signal I15717: std_logic; attribute dont_touch of I15717: signal is true;
	signal I15718: std_logic; attribute dont_touch of I15718: signal is true;
	signal I15725: std_logic; attribute dont_touch of I15725: signal is true;
	signal I15729: std_logic; attribute dont_touch of I15729: signal is true;
	signal I15733: std_logic; attribute dont_touch of I15733: signal is true;
	signal I15736: std_logic; attribute dont_touch of I15736: signal is true;
	signal I15741: std_logic; attribute dont_touch of I15741: signal is true;
	signal I15744: std_logic; attribute dont_touch of I15744: signal is true;
	signal I15749: std_logic; attribute dont_touch of I15749: signal is true;
	signal I15752: std_logic; attribute dont_touch of I15752: signal is true;
	signal I15756: std_logic; attribute dont_touch of I15756: signal is true;
	signal I15759: std_logic; attribute dont_touch of I15759: signal is true;
	signal I15763: std_logic; attribute dont_touch of I15763: signal is true;
	signal I15768: std_logic; attribute dont_touch of I15768: signal is true;
	signal I15771: std_logic; attribute dont_touch of I15771: signal is true;
	signal I15775: std_logic; attribute dont_touch of I15775: signal is true;
	signal I15778: std_logic; attribute dont_touch of I15778: signal is true;
	signal I15782: std_logic; attribute dont_touch of I15782: signal is true;
	signal I15787: std_logic; attribute dont_touch of I15787: signal is true;
	signal I15792: std_logic; attribute dont_touch of I15792: signal is true;
	signal I15795: std_logic; attribute dont_touch of I15795: signal is true;
	signal I15798: std_logic; attribute dont_touch of I15798: signal is true;
	signal I15801: std_logic; attribute dont_touch of I15801: signal is true;
	signal I15804: std_logic; attribute dont_touch of I15804: signal is true;
	signal I15807: std_logic; attribute dont_touch of I15807: signal is true;
	signal I15811: std_logic; attribute dont_touch of I15811: signal is true;
	signal I15814: std_logic; attribute dont_touch of I15814: signal is true;
	signal I15817: std_logic; attribute dont_touch of I15817: signal is true;
	signal I15820: std_logic; attribute dont_touch of I15820: signal is true;
	signal I15823: std_logic; attribute dont_touch of I15823: signal is true;
	signal I15826: std_logic; attribute dont_touch of I15826: signal is true;
	signal I15829: std_logic; attribute dont_touch of I15829: signal is true;
	signal I15832: std_logic; attribute dont_touch of I15832: signal is true;
	signal I15855: std_logic; attribute dont_touch of I15855: signal is true;
	signal I15858: std_logic; attribute dont_touch of I15858: signal is true;
	signal I15861: std_logic; attribute dont_touch of I15861: signal is true;
	signal I15864: std_logic; attribute dont_touch of I15864: signal is true;
	signal I15870: std_logic; attribute dont_touch of I15870: signal is true;
	signal I15871: std_logic; attribute dont_touch of I15871: signal is true;
	signal I15872: std_logic; attribute dont_touch of I15872: signal is true;
	signal I15878: std_logic; attribute dont_touch of I15878: signal is true;
	signal I15879: std_logic; attribute dont_touch of I15879: signal is true;
	signal I15880: std_logic; attribute dont_touch of I15880: signal is true;
	signal I15890: std_logic; attribute dont_touch of I15890: signal is true;
	signal I15891: std_logic; attribute dont_touch of I15891: signal is true;
	signal I15892: std_logic; attribute dont_touch of I15892: signal is true;
	signal I15898: std_logic; attribute dont_touch of I15898: signal is true;
	signal I15899: std_logic; attribute dont_touch of I15899: signal is true;
	signal I15900: std_logic; attribute dont_touch of I15900: signal is true;
	signal I15906: std_logic; attribute dont_touch of I15906: signal is true;
	signal I15907: std_logic; attribute dont_touch of I15907: signal is true;
	signal I15908: std_logic; attribute dont_touch of I15908: signal is true;
	signal I15956: std_logic; attribute dont_touch of I15956: signal is true;
	signal I15959: std_logic; attribute dont_touch of I15959: signal is true;
	signal I15962: std_logic; attribute dont_touch of I15962: signal is true;
	signal I15965: std_logic; attribute dont_touch of I15965: signal is true;
	signal I15968: std_logic; attribute dont_touch of I15968: signal is true;
	signal I15971: std_logic; attribute dont_touch of I15971: signal is true;
	signal I15974: std_logic; attribute dont_touch of I15974: signal is true;
	signal I15977: std_logic; attribute dont_touch of I15977: signal is true;
	signal I15980: std_logic; attribute dont_touch of I15980: signal is true;
	signal I15983: std_logic; attribute dont_touch of I15983: signal is true;
	signal I15986: std_logic; attribute dont_touch of I15986: signal is true;
	signal I15989: std_logic; attribute dont_touch of I15989: signal is true;
	signal I15992: std_logic; attribute dont_touch of I15992: signal is true;
	signal I15993: std_logic; attribute dont_touch of I15993: signal is true;
	signal I15994: std_logic; attribute dont_touch of I15994: signal is true;
	signal I15999: std_logic; attribute dont_touch of I15999: signal is true;
	signal I16000: std_logic; attribute dont_touch of I16000: signal is true;
	signal I16001: std_logic; attribute dont_touch of I16001: signal is true;
	signal I16007: std_logic; attribute dont_touch of I16007: signal is true;
	signal I16008: std_logic; attribute dont_touch of I16008: signal is true;
	signal I16009: std_logic; attribute dont_touch of I16009: signal is true;
	signal I16015: std_logic; attribute dont_touch of I16015: signal is true;
	signal I16016: std_logic; attribute dont_touch of I16016: signal is true;
	signal I16017: std_logic; attribute dont_touch of I16017: signal is true;
	signal I16023: std_logic; attribute dont_touch of I16023: signal is true;
	signal I16024: std_logic; attribute dont_touch of I16024: signal is true;
	signal I16025: std_logic; attribute dont_touch of I16025: signal is true;
	signal I16030: std_logic; attribute dont_touch of I16030: signal is true;
	signal I16031: std_logic; attribute dont_touch of I16031: signal is true;
	signal I16032: std_logic; attribute dont_touch of I16032: signal is true;
	signal I16037: std_logic; attribute dont_touch of I16037: signal is true;
	signal I16038: std_logic; attribute dont_touch of I16038: signal is true;
	signal I16039: std_logic; attribute dont_touch of I16039: signal is true;
	signal I16044: std_logic; attribute dont_touch of I16044: signal is true;
	signal I16045: std_logic; attribute dont_touch of I16045: signal is true;
	signal I16046: std_logic; attribute dont_touch of I16046: signal is true;
	signal I16051: std_logic; attribute dont_touch of I16051: signal is true;
	signal I16052: std_logic; attribute dont_touch of I16052: signal is true;
	signal I16053: std_logic; attribute dont_touch of I16053: signal is true;
	signal I16058: std_logic; attribute dont_touch of I16058: signal is true;
	signal I16059: std_logic; attribute dont_touch of I16059: signal is true;
	signal I16060: std_logic; attribute dont_touch of I16060: signal is true;
	signal I16065: std_logic; attribute dont_touch of I16065: signal is true;
	signal I16066: std_logic; attribute dont_touch of I16066: signal is true;
	signal I16067: std_logic; attribute dont_touch of I16067: signal is true;
	signal I16072: std_logic; attribute dont_touch of I16072: signal is true;
	signal I16073: std_logic; attribute dont_touch of I16073: signal is true;
	signal I16074: std_logic; attribute dont_touch of I16074: signal is true;
	signal I16079: std_logic; attribute dont_touch of I16079: signal is true;
	signal I16080: std_logic; attribute dont_touch of I16080: signal is true;
	signal I16081: std_logic; attribute dont_touch of I16081: signal is true;
	signal I16086: std_logic; attribute dont_touch of I16086: signal is true;
	signal I16087: std_logic; attribute dont_touch of I16087: signal is true;
	signal I16088: std_logic; attribute dont_touch of I16088: signal is true;
	signal I16095: std_logic; attribute dont_touch of I16095: signal is true;
	signal I16098: std_logic; attribute dont_touch of I16098: signal is true;
	signal I16101: std_logic; attribute dont_touch of I16101: signal is true;
	signal I16105: std_logic; attribute dont_touch of I16105: signal is true;
	signal I16108: std_logic; attribute dont_touch of I16108: signal is true;
	signal I16111: std_logic; attribute dont_touch of I16111: signal is true;
	signal I16114: std_logic; attribute dont_touch of I16114: signal is true;
	signal I16121: std_logic; attribute dont_touch of I16121: signal is true;
	signal I16124: std_logic; attribute dont_touch of I16124: signal is true;
	signal I16142: std_logic; attribute dont_touch of I16142: signal is true;
	signal I16145: std_logic; attribute dont_touch of I16145: signal is true;
	signal I16148: std_logic; attribute dont_touch of I16148: signal is true;
	signal I16149: std_logic; attribute dont_touch of I16149: signal is true;
	signal I16160: std_logic; attribute dont_touch of I16160: signal is true;
	signal I16161: std_logic; attribute dont_touch of I16161: signal is true;
	signal I16169: std_logic; attribute dont_touch of I16169: signal is true;
	signal I16172: std_logic; attribute dont_touch of I16172: signal is true;
	signal I16175: std_logic; attribute dont_touch of I16175: signal is true;
	signal I16178: std_logic; attribute dont_touch of I16178: signal is true;
	signal I16181: std_logic; attribute dont_touch of I16181: signal is true;
	signal I16184: std_logic; attribute dont_touch of I16184: signal is true;
	signal I16187: std_logic; attribute dont_touch of I16187: signal is true;
	signal I16190: std_logic; attribute dont_touch of I16190: signal is true;
	signal I16193: std_logic; attribute dont_touch of I16193: signal is true;
	signal I16196: std_logic; attribute dont_touch of I16196: signal is true;
	signal I16200: std_logic; attribute dont_touch of I16200: signal is true;
	signal I16203: std_logic; attribute dont_touch of I16203: signal is true;
	signal I16206: std_logic; attribute dont_touch of I16206: signal is true;
	signal I16209: std_logic; attribute dont_touch of I16209: signal is true;
	signal I16214: std_logic; attribute dont_touch of I16214: signal is true;
	signal I16217: std_logic; attribute dont_touch of I16217: signal is true;
	signal I16220: std_logic; attribute dont_touch of I16220: signal is true;
	signal I16236: std_logic; attribute dont_touch of I16236: signal is true;
	signal I16239: std_logic; attribute dont_touch of I16239: signal is true;
	signal I16252: std_logic; attribute dont_touch of I16252: signal is true;
	signal I16255: std_logic; attribute dont_touch of I16255: signal is true;
	signal I16258: std_logic; attribute dont_touch of I16258: signal is true;
	signal I16261: std_logic; attribute dont_touch of I16261: signal is true;
	signal I16264: std_logic; attribute dont_touch of I16264: signal is true;
	signal I16269: std_logic; attribute dont_touch of I16269: signal is true;
	signal I16273: std_logic; attribute dont_touch of I16273: signal is true;
	signal I16277: std_logic; attribute dont_touch of I16277: signal is true;
	signal I16280: std_logic; attribute dont_touch of I16280: signal is true;
	signal I16283: std_logic; attribute dont_touch of I16283: signal is true;
	signal I16286: std_logic; attribute dont_touch of I16286: signal is true;
	signal I16289: std_logic; attribute dont_touch of I16289: signal is true;
	signal I16292: std_logic; attribute dont_touch of I16292: signal is true;
	signal I16295: std_logic; attribute dont_touch of I16295: signal is true;
	signal I16298: std_logic; attribute dont_touch of I16298: signal is true;
	signal I16307: std_logic; attribute dont_touch of I16307: signal is true;
	signal I16311: std_logic; attribute dont_touch of I16311: signal is true;
	signal I16330: std_logic; attribute dont_touch of I16330: signal is true;
	signal I16331: std_logic; attribute dont_touch of I16331: signal is true;
	signal I16332: std_logic; attribute dont_touch of I16332: signal is true;
	signal I16356: std_logic; attribute dont_touch of I16356: signal is true;
	signal I16360: std_logic; attribute dont_touch of I16360: signal is true;
	signal I16363: std_logic; attribute dont_touch of I16363: signal is true;
	signal I16366: std_logic; attribute dont_touch of I16366: signal is true;
	signal I16370: std_logic; attribute dont_touch of I16370: signal is true;
	signal I16373: std_logic; attribute dont_touch of I16373: signal is true;
	signal I16376: std_logic; attribute dont_touch of I16376: signal is true;
	signal I16379: std_logic; attribute dont_touch of I16379: signal is true;
	signal I16387: std_logic; attribute dont_touch of I16387: signal is true;
	signal I16407: std_logic; attribute dont_touch of I16407: signal is true;
	signal I16413: std_logic; attribute dont_touch of I16413: signal is true;
	signal I16416: std_logic; attribute dont_touch of I16416: signal is true;
	signal I16427: std_logic; attribute dont_touch of I16427: signal is true;
	signal I16432: std_logic; attribute dont_touch of I16432: signal is true;
	signal I16439: std_logic; attribute dont_touch of I16439: signal is true;
	signal I16458: std_logic; attribute dont_touch of I16458: signal is true;
	signal I16461: std_logic; attribute dont_touch of I16461: signal is true;
	signal I16467: std_logic; attribute dont_touch of I16467: signal is true;
	signal I16468: std_logic; attribute dont_touch of I16468: signal is true;
	signal I16469: std_logic; attribute dont_touch of I16469: signal is true;
	signal I16475: std_logic; attribute dont_touch of I16475: signal is true;
	signal I16479: std_logic; attribute dont_touch of I16479: signal is true;
	signal I16484: std_logic; attribute dont_touch of I16484: signal is true;
	signal I16487: std_logic; attribute dont_touch of I16487: signal is true;
	signal I16492: std_logic; attribute dont_touch of I16492: signal is true;
	signal I16496: std_logic; attribute dont_touch of I16496: signal is true;
	signal I16500: std_logic; attribute dont_touch of I16500: signal is true;
	signal I16507: std_logic; attribute dont_touch of I16507: signal is true;
	signal I16510: std_logic; attribute dont_touch of I16510: signal is true;
	signal I16514: std_logic; attribute dont_touch of I16514: signal is true;
	signal I16518: std_logic; attribute dont_touch of I16518: signal is true;
	signal I16525: std_logic; attribute dont_touch of I16525: signal is true;
	signal I16528: std_logic; attribute dont_touch of I16528: signal is true;
	signal I16531: std_logic; attribute dont_touch of I16531: signal is true;
	signal I16534: std_logic; attribute dont_touch of I16534: signal is true;
	signal I16537: std_logic; attribute dont_touch of I16537: signal is true;
	signal I16540: std_logic; attribute dont_touch of I16540: signal is true;
	signal I16543: std_logic; attribute dont_touch of I16543: signal is true;
	signal I16546: std_logic; attribute dont_touch of I16546: signal is true;
	signal I16550: std_logic; attribute dont_touch of I16550: signal is true;
	signal I16553: std_logic; attribute dont_touch of I16553: signal is true;
	signal I16571: std_logic; attribute dont_touch of I16571: signal is true;
	signal I16574: std_logic; attribute dont_touch of I16574: signal is true;
	signal I16577: std_logic; attribute dont_touch of I16577: signal is true;
	signal I16580: std_logic; attribute dont_touch of I16580: signal is true;
	signal I16583: std_logic; attribute dont_touch of I16583: signal is true;
	signal I16586: std_logic; attribute dont_touch of I16586: signal is true;
	signal I16589: std_logic; attribute dont_touch of I16589: signal is true;
	signal I16592: std_logic; attribute dont_touch of I16592: signal is true;
	signal I16595: std_logic; attribute dont_touch of I16595: signal is true;
	signal I16598: std_logic; attribute dont_touch of I16598: signal is true;
	signal I16601: std_logic; attribute dont_touch of I16601: signal is true;
	signal I16604: std_logic; attribute dont_touch of I16604: signal is true;
	signal I16607: std_logic; attribute dont_touch of I16607: signal is true;
	signal I16610: std_logic; attribute dont_touch of I16610: signal is true;
	signal I16613: std_logic; attribute dont_touch of I16613: signal is true;
	signal I16616: std_logic; attribute dont_touch of I16616: signal is true;
	signal I16623: std_logic; attribute dont_touch of I16623: signal is true;
	signal I16626: std_logic; attribute dont_touch of I16626: signal is true;
	signal I16629: std_logic; attribute dont_touch of I16629: signal is true;
	signal I16632: std_logic; attribute dont_touch of I16632: signal is true;
	signal I16635: std_logic; attribute dont_touch of I16635: signal is true;
	signal I16638: std_logic; attribute dont_touch of I16638: signal is true;
	signal I16641: std_logic; attribute dont_touch of I16641: signal is true;
	signal I16644: std_logic; attribute dont_touch of I16644: signal is true;
	signal I16647: std_logic; attribute dont_touch of I16647: signal is true;
	signal I16650: std_logic; attribute dont_touch of I16650: signal is true;
	signal I16656: std_logic; attribute dont_touch of I16656: signal is true;
	signal I16660: std_logic; attribute dont_touch of I16660: signal is true;
	signal I16664: std_logic; attribute dont_touch of I16664: signal is true;
	signal I16667: std_logic; attribute dont_touch of I16667: signal is true;
	signal I16670: std_logic; attribute dont_touch of I16670: signal is true;
	signal I16673: std_logic; attribute dont_touch of I16673: signal is true;
	signal I16676: std_logic; attribute dont_touch of I16676: signal is true;
	signal I16679: std_logic; attribute dont_touch of I16679: signal is true;
	signal I16682: std_logic; attribute dont_touch of I16682: signal is true;
	signal I16685: std_logic; attribute dont_touch of I16685: signal is true;
	signal I16688: std_logic; attribute dont_touch of I16688: signal is true;
	signal I16691: std_logic; attribute dont_touch of I16691: signal is true;
	signal I16708: std_logic; attribute dont_touch of I16708: signal is true;
	signal I16717: std_logic; attribute dont_touch of I16717: signal is true;
	signal I16720: std_logic; attribute dont_touch of I16720: signal is true;
	signal I16723: std_logic; attribute dont_touch of I16723: signal is true;
	signal I16735: std_logic; attribute dont_touch of I16735: signal is true;
	signal I16739: std_logic; attribute dont_touch of I16739: signal is true;
	signal I16742: std_logic; attribute dont_touch of I16742: signal is true;
	signal I16760: std_logic; attribute dont_touch of I16760: signal is true;
	signal I16763: std_logic; attribute dont_touch of I16763: signal is true;
	signal I16766: std_logic; attribute dont_touch of I16766: signal is true;
	signal I16769: std_logic; attribute dont_touch of I16769: signal is true;
	signal I16772: std_logic; attribute dont_touch of I16772: signal is true;
	signal I16775: std_logic; attribute dont_touch of I16775: signal is true;
	signal I16778: std_logic; attribute dont_touch of I16778: signal is true;
	signal I16781: std_logic; attribute dont_touch of I16781: signal is true;
	signal I16784: std_logic; attribute dont_touch of I16784: signal is true;
	signal I16787: std_logic; attribute dont_touch of I16787: signal is true;
	signal I16790: std_logic; attribute dont_touch of I16790: signal is true;
	signal I16793: std_logic; attribute dont_touch of I16793: signal is true;
	signal I16796: std_logic; attribute dont_touch of I16796: signal is true;
	signal I16799: std_logic; attribute dont_touch of I16799: signal is true;
	signal I16802: std_logic; attribute dont_touch of I16802: signal is true;
	signal I16805: std_logic; attribute dont_touch of I16805: signal is true;
	signal I16808: std_logic; attribute dont_touch of I16808: signal is true;
	signal I16811: std_logic; attribute dont_touch of I16811: signal is true;
	signal I16814: std_logic; attribute dont_touch of I16814: signal is true;
	signal I16817: std_logic; attribute dont_touch of I16817: signal is true;
	signal I16843: std_logic; attribute dont_touch of I16843: signal is true;
	signal I16847: std_logic; attribute dont_touch of I16847: signal is true;
	signal I16850: std_logic; attribute dont_touch of I16850: signal is true;
	signal I16853: std_logic; attribute dont_touch of I16853: signal is true;
	signal I16856: std_logic; attribute dont_touch of I16856: signal is true;
	signal I16859: std_logic; attribute dont_touch of I16859: signal is true;
	signal I16863: std_logic; attribute dont_touch of I16863: signal is true;
	signal I16867: std_logic; attribute dont_touch of I16867: signal is true;
	signal I16871: std_logic; attribute dont_touch of I16871: signal is true;
	signal I16879: std_logic; attribute dont_touch of I16879: signal is true;
	signal I16897: std_logic; attribute dont_touch of I16897: signal is true;
	signal I16920: std_logic; attribute dont_touch of I16920: signal is true;
	signal I16938: std_logic; attribute dont_touch of I16938: signal is true;
	signal I16941: std_logic; attribute dont_touch of I16941: signal is true;
	signal I16944: std_logic; attribute dont_touch of I16944: signal is true;
	signal I16947: std_logic; attribute dont_touch of I16947: signal is true;
	signal I16950: std_logic; attribute dont_touch of I16950: signal is true;
	signal I16953: std_logic; attribute dont_touch of I16953: signal is true;
	signal I16956: std_logic; attribute dont_touch of I16956: signal is true;
	signal I16979: std_logic; attribute dont_touch of I16979: signal is true;
	signal I16982: std_logic; attribute dont_touch of I16982: signal is true;
	signal I17051: std_logic; attribute dont_touch of I17051: signal is true;
	signal I17052: std_logic; attribute dont_touch of I17052: signal is true;
	signal I17053: std_logic; attribute dont_touch of I17053: signal is true;
	signal I17070: std_logic; attribute dont_touch of I17070: signal is true;
	signal I17084: std_logic; attribute dont_touch of I17084: signal is true;
	signal I17092: std_logic; attribute dont_touch of I17092: signal is true;
	signal I17096: std_logic; attribute dont_touch of I17096: signal is true;
	signal I17100: std_logic; attribute dont_touch of I17100: signal is true;
	signal I17104: std_logic; attribute dont_touch of I17104: signal is true;
	signal I17108: std_logic; attribute dont_touch of I17108: signal is true;
	signal I17112: std_logic; attribute dont_touch of I17112: signal is true;
	signal I17116: std_logic; attribute dont_touch of I17116: signal is true;
	signal I17121: std_logic; attribute dont_touch of I17121: signal is true;
	signal I17124: std_logic; attribute dont_touch of I17124: signal is true;
	signal I17142: std_logic; attribute dont_touch of I17142: signal is true;
	signal I17146: std_logic; attribute dont_touch of I17146: signal is true;
	signal I17149: std_logic; attribute dont_touch of I17149: signal is true;
	signal I17152: std_logic; attribute dont_touch of I17152: signal is true;
	signal I17155: std_logic; attribute dont_touch of I17155: signal is true;
	signal I17158: std_logic; attribute dont_touch of I17158: signal is true;
	signal I17161: std_logic; attribute dont_touch of I17161: signal is true;
	signal I17164: std_logic; attribute dont_touch of I17164: signal is true;
	signal I17170: std_logic; attribute dont_touch of I17170: signal is true;
	signal I17173: std_logic; attribute dont_touch of I17173: signal is true;
	signal I17176: std_logic; attribute dont_touch of I17176: signal is true;
	signal I17179: std_logic; attribute dont_touch of I17179: signal is true;
	signal I17182: std_logic; attribute dont_touch of I17182: signal is true;
	signal I17185: std_logic; attribute dont_touch of I17185: signal is true;
	signal I17188: std_logic; attribute dont_touch of I17188: signal is true;
	signal I17191: std_logic; attribute dont_touch of I17191: signal is true;
	signal I17194: std_logic; attribute dont_touch of I17194: signal is true;
	signal I17198: std_logic; attribute dont_touch of I17198: signal is true;
	signal I17202: std_logic; attribute dont_touch of I17202: signal is true;
	signal I17206: std_logic; attribute dont_touch of I17206: signal is true;
	signal I17209: std_logic; attribute dont_touch of I17209: signal is true;
	signal I17213: std_logic; attribute dont_touch of I17213: signal is true;
	signal I17216: std_logic; attribute dont_touch of I17216: signal is true;
	signal I17219: std_logic; attribute dont_touch of I17219: signal is true;
	signal I17225: std_logic; attribute dont_touch of I17225: signal is true;
	signal I17228: std_logic; attribute dont_touch of I17228: signal is true;
	signal I17231: std_logic; attribute dont_touch of I17231: signal is true;
	signal I17234: std_logic; attribute dont_touch of I17234: signal is true;
	signal I17237: std_logic; attribute dont_touch of I17237: signal is true;
	signal I17240: std_logic; attribute dont_touch of I17240: signal is true;
	signal I17243: std_logic; attribute dont_touch of I17243: signal is true;
	signal I17246: std_logic; attribute dont_touch of I17246: signal is true;
	signal I17249: std_logic; attribute dont_touch of I17249: signal is true;
	signal I17252: std_logic; attribute dont_touch of I17252: signal is true;
	signal I17255: std_logic; attribute dont_touch of I17255: signal is true;
	signal I17258: std_logic; attribute dont_touch of I17258: signal is true;
	signal I17261: std_logic; attribute dont_touch of I17261: signal is true;
	signal I17265: std_logic; attribute dont_touch of I17265: signal is true;
	signal I17268: std_logic; attribute dont_touch of I17268: signal is true;
	signal I17271: std_logic; attribute dont_touch of I17271: signal is true;
	signal I17274: std_logic; attribute dont_touch of I17274: signal is true;
	signal I17277: std_logic; attribute dont_touch of I17277: signal is true;
	signal I17281: std_logic; attribute dont_touch of I17281: signal is true;
	signal I17282: std_logic; attribute dont_touch of I17282: signal is true;
	signal I17283: std_logic; attribute dont_touch of I17283: signal is true;
	signal I17288: std_logic; attribute dont_touch of I17288: signal is true;
	signal I17289: std_logic; attribute dont_touch of I17289: signal is true;
	signal I17290: std_logic; attribute dont_touch of I17290: signal is true;
	signal I17295: std_logic; attribute dont_touch of I17295: signal is true;
	signal I17296: std_logic; attribute dont_touch of I17296: signal is true;
	signal I17297: std_logic; attribute dont_touch of I17297: signal is true;
	signal I17302: std_logic; attribute dont_touch of I17302: signal is true;
	signal I17305: std_logic; attribute dont_touch of I17305: signal is true;
	signal I17306: std_logic; attribute dont_touch of I17306: signal is true;
	signal I17307: std_logic; attribute dont_touch of I17307: signal is true;
	signal I17312: std_logic; attribute dont_touch of I17312: signal is true;
	signal I17315: std_logic; attribute dont_touch of I17315: signal is true;
	signal I17318: std_logic; attribute dont_touch of I17318: signal is true;
	signal I17321: std_logic; attribute dont_touch of I17321: signal is true;
	signal I17324: std_logic; attribute dont_touch of I17324: signal is true;
	signal I17327: std_logic; attribute dont_touch of I17327: signal is true;
	signal I17331: std_logic; attribute dont_touch of I17331: signal is true;
	signal I17334: std_logic; attribute dont_touch of I17334: signal is true;
	signal I17337: std_logic; attribute dont_touch of I17337: signal is true;
	signal I17340: std_logic; attribute dont_touch of I17340: signal is true;
	signal I17344: std_logic; attribute dont_touch of I17344: signal is true;
	signal I17347: std_logic; attribute dont_touch of I17347: signal is true;
	signal I17350: std_logic; attribute dont_touch of I17350: signal is true;
	signal I17353: std_logic; attribute dont_touch of I17353: signal is true;
	signal I17356: std_logic; attribute dont_touch of I17356: signal is true;
	signal I17359: std_logic; attribute dont_touch of I17359: signal is true;
	signal I17362: std_logic; attribute dont_touch of I17362: signal is true;
	signal I17365: std_logic; attribute dont_touch of I17365: signal is true;
	signal I17368: std_logic; attribute dont_touch of I17368: signal is true;
	signal I17371: std_logic; attribute dont_touch of I17371: signal is true;
	signal I17374: std_logic; attribute dont_touch of I17374: signal is true;
	signal I17377: std_logic; attribute dont_touch of I17377: signal is true;
	signal I17381: std_logic; attribute dont_touch of I17381: signal is true;
	signal I17384: std_logic; attribute dont_touch of I17384: signal is true;
	signal I17387: std_logic; attribute dont_touch of I17387: signal is true;
	signal I17390: std_logic; attribute dont_touch of I17390: signal is true;
	signal I17393: std_logic; attribute dont_touch of I17393: signal is true;
	signal I17394: std_logic; attribute dont_touch of I17394: signal is true;
	signal I17395: std_logic; attribute dont_touch of I17395: signal is true;
	signal I17400: std_logic; attribute dont_touch of I17400: signal is true;
	signal I17401: std_logic; attribute dont_touch of I17401: signal is true;
	signal I17402: std_logic; attribute dont_touch of I17402: signal is true;
	signal I17407: std_logic; attribute dont_touch of I17407: signal is true;
	signal I17410: std_logic; attribute dont_touch of I17410: signal is true;
	signal I17413: std_logic; attribute dont_touch of I17413: signal is true;
	signal I17416: std_logic; attribute dont_touch of I17416: signal is true;
	signal I17419: std_logic; attribute dont_touch of I17419: signal is true;
	signal I17424: std_logic; attribute dont_touch of I17424: signal is true;
	signal I17435: std_logic; attribute dont_touch of I17435: signal is true;
	signal I17438: std_logic; attribute dont_touch of I17438: signal is true;
	signal I17441: std_logic; attribute dont_touch of I17441: signal is true;
	signal I17444: std_logic; attribute dont_touch of I17444: signal is true;
	signal I17447: std_logic; attribute dont_touch of I17447: signal is true;
	signal I17450: std_logic; attribute dont_touch of I17450: signal is true;
	signal I17453: std_logic; attribute dont_touch of I17453: signal is true;
	signal I17456: std_logic; attribute dont_touch of I17456: signal is true;
	signal I17459: std_logic; attribute dont_touch of I17459: signal is true;
	signal I17460: std_logic; attribute dont_touch of I17460: signal is true;
	signal I17461: std_logic; attribute dont_touch of I17461: signal is true;
	signal I17466: std_logic; attribute dont_touch of I17466: signal is true;
	signal I17470: std_logic; attribute dont_touch of I17470: signal is true;
	signal I17482: std_logic; attribute dont_touch of I17482: signal is true;
	signal I17485: std_logic; attribute dont_touch of I17485: signal is true;
	signal I17486: std_logic; attribute dont_touch of I17486: signal is true;
	signal I17487: std_logic; attribute dont_touch of I17487: signal is true;
	signal I17492: std_logic; attribute dont_touch of I17492: signal is true;
	signal I17493: std_logic; attribute dont_touch of I17493: signal is true;
	signal I17494: std_logic; attribute dont_touch of I17494: signal is true;
	signal I17500: std_logic; attribute dont_touch of I17500: signal is true;
	signal I17503: std_logic; attribute dont_touch of I17503: signal is true;
	signal I17504: std_logic; attribute dont_touch of I17504: signal is true;
	signal I17505: std_logic; attribute dont_touch of I17505: signal is true;
	signal I17510: std_logic; attribute dont_touch of I17510: signal is true;
	signal I17513: std_logic; attribute dont_touch of I17513: signal is true;
	signal I17516: std_logic; attribute dont_touch of I17516: signal is true;
	signal I17519: std_logic; attribute dont_touch of I17519: signal is true;
	signal I17522: std_logic; attribute dont_touch of I17522: signal is true;
	signal I17525: std_logic; attribute dont_touch of I17525: signal is true;
	signal I17528: std_logic; attribute dont_touch of I17528: signal is true;
	signal I17531: std_logic; attribute dont_touch of I17531: signal is true;
	signal I17534: std_logic; attribute dont_touch of I17534: signal is true;
	signal I17537: std_logic; attribute dont_touch of I17537: signal is true;
	signal I17540: std_logic; attribute dont_touch of I17540: signal is true;
	signal I17543: std_logic; attribute dont_touch of I17543: signal is true;
	signal I17546: std_logic; attribute dont_touch of I17546: signal is true;
	signal I17549: std_logic; attribute dont_touch of I17549: signal is true;
	signal I17552: std_logic; attribute dont_touch of I17552: signal is true;
	signal I17555: std_logic; attribute dont_touch of I17555: signal is true;
	signal I17558: std_logic; attribute dont_touch of I17558: signal is true;
	signal I17563: std_logic; attribute dont_touch of I17563: signal is true;
	signal I17567: std_logic; attribute dont_touch of I17567: signal is true;
	signal I17568: std_logic; attribute dont_touch of I17568: signal is true;
	signal I17569: std_logic; attribute dont_touch of I17569: signal is true;
	signal I17584: std_logic; attribute dont_touch of I17584: signal is true;
	signal I17585: std_logic; attribute dont_touch of I17585: signal is true;
	signal I17586: std_logic; attribute dont_touch of I17586: signal is true;
	signal I17591: std_logic; attribute dont_touch of I17591: signal is true;
	signal I17610: std_logic; attribute dont_touch of I17610: signal is true;
	signal I17613: std_logic; attribute dont_touch of I17613: signal is true;
	signal I17616: std_logic; attribute dont_touch of I17616: signal is true;
	signal I17633: std_logic; attribute dont_touch of I17633: signal is true;
	signal I17636: std_logic; attribute dont_touch of I17636: signal is true;
	signal I17642: std_logic; attribute dont_touch of I17642: signal is true;
	signal I17657: std_logic; attribute dont_touch of I17657: signal is true;
	signal I17662: std_logic; attribute dont_touch of I17662: signal is true;
	signal I17666: std_logic; attribute dont_touch of I17666: signal is true;
	signal I17669: std_logic; attribute dont_touch of I17669: signal is true;
	signal I17672: std_logic; attribute dont_touch of I17672: signal is true;
	signal I17675: std_logic; attribute dont_touch of I17675: signal is true;
	signal I17678: std_logic; attribute dont_touch of I17678: signal is true;
	signal I17681: std_logic; attribute dont_touch of I17681: signal is true;
	signal I17684: std_logic; attribute dont_touch of I17684: signal is true;
	signal I17687: std_logic; attribute dont_touch of I17687: signal is true;
	signal I17692: std_logic; attribute dont_touch of I17692: signal is true;
	signal I17695: std_logic; attribute dont_touch of I17695: signal is true;
	signal I17698: std_logic; attribute dont_touch of I17698: signal is true;
	signal I17701: std_logic; attribute dont_touch of I17701: signal is true;
	signal I17704: std_logic; attribute dont_touch of I17704: signal is true;
	signal I17707: std_logic; attribute dont_touch of I17707: signal is true;
	signal I17710: std_logic; attribute dont_touch of I17710: signal is true;
	signal I17713: std_logic; attribute dont_touch of I17713: signal is true;
	signal I17716: std_logic; attribute dont_touch of I17716: signal is true;
	signal I17719: std_logic; attribute dont_touch of I17719: signal is true;
	signal I17724: std_logic; attribute dont_touch of I17724: signal is true;
	signal I17730: std_logic; attribute dont_touch of I17730: signal is true;
	signal I17733: std_logic; attribute dont_touch of I17733: signal is true;
	signal I17736: std_logic; attribute dont_touch of I17736: signal is true;
	signal I17739: std_logic; attribute dont_touch of I17739: signal is true;
	signal I17742: std_logic; attribute dont_touch of I17742: signal is true;
	signal I17746: std_logic; attribute dont_touch of I17746: signal is true;
	signal I17749: std_logic; attribute dont_touch of I17749: signal is true;
	signal I17752: std_logic; attribute dont_touch of I17752: signal is true;
	signal I17755: std_logic; attribute dont_touch of I17755: signal is true;
	signal I17758: std_logic; attribute dont_touch of I17758: signal is true;
	signal I17761: std_logic; attribute dont_touch of I17761: signal is true;
	signal I17764: std_logic; attribute dont_touch of I17764: signal is true;
	signal I17767: std_logic; attribute dont_touch of I17767: signal is true;
	signal I17770: std_logic; attribute dont_touch of I17770: signal is true;
	signal I17773: std_logic; attribute dont_touch of I17773: signal is true;
begin
	process(CLK)
	begin
		if(rising_edge(CLK)) then
			G1<=G8078;
			G4<=G8079;
			G7<=G2731;
			G8<=G2613;
			G9<=G7336;
			G12<=G7337;
			G16<=G4906;
			G17<=G4894;
			G26<=G4885;
			G32<=G11397;
			G33<=G10867;
			G34<=G10868;
			G35<=G10869;
			G36<=G10870;
			G37<=G10871;
			G38<=G10872;
			G39<=G10774;
			G40<=G10775;
			G49<=G7774;
			G52<=G7777;
			G55<=G7778;
			G58<=G7779;
			G61<=G7780;
			G64<=G7781;
			G67<=G7782;
			G70<=G7783;
			G73<=G7784;
			G76<=G7775;
			G79<=G7776;
			G105<=G11180;
			G108<=G11593;
			G113<=G7285;
			G114<=G113;
			G115<=G7321;
			G119<=G7745;
			G123<=G8272;
			G126<=G5642;
			G127<=G8421;
			G131<=G8420;
			G135<=G8419;
			G139<=G8418;
			G143<=G7746;
			G148<=G8427;
			G153<=G8426;
			G158<=G8425;
			G162<=G8424;
			G166<=G7747;
			G170<=G8422;
			G174<=G8423;
			G178<=G7748;
			G182<=G7749;
			G186<=G7317;
			G192<=G6837;
			G197<=G6835;
			G201<=G7304;
			G207<=G7315;
			G213<=G7313;
			G219<=G7310;
			G225<=G7309;
			G231<=G7319;
			G237<=G7306;
			G243<=G7325;
			G248<=G7323;
			G253<=G7750;
			G254<=G7759;
			G255<=G7751;
			G256<=G7752;
			G257<=G7753;
			G258<=G7754;
			G259<=G7755;
			G260<=G7756;
			G261<=G7757;
			G262<=G7758;
			G263<=G7760;
			G266<=G7761;
			G269<=G7762;
			G272<=G7763;
			G275<=G7764;
			G278<=G7765;
			G281<=G7766;
			G284<=G7767;
			G287<=G7768;
			G290<=G7769;
			G293<=G7770;
			G296<=G7771;
			G299<=G7772;
			G302<=G7773;
			G305<=G5643;
			G309<=G5652;
			G312<=G5644;
			G315<=G5645;
			G318<=G5646;
			G321<=G5647;
			G324<=G5648;
			G327<=G5649;
			G330<=G5650;
			G333<=G5651;
			G336<=G11653;
			G339<=G11505;
			G342<=G11513;
			G345<=G11642;
			G348<=G11506;
			G351<=G11507;
			G354<=G11508;
			G357<=G11509;
			G360<=G11510;
			G363<=G11511;
			G366<=G11512;
			G369<=G11439;
			G374<=G11440;
			G378<=G11441;
			G382<=G11442;
			G386<=G11263;
			G391<=G11264;
			G396<=G11265;
			G401<=G11266;
			G406<=G11267;
			G411<=G11268;
			G416<=G11269;
			G421<=G11270;
			G426<=G11256;
			G431<=G11262;
			G435<=G11261;
			G440<=G11260;
			G444<=G11259;
			G448<=G11258;
			G452<=G11257;
			G456<=G11466;
			G461<=G11467;
			G466<=G11468;
			G471<=G11469;
			G476<=G11338;
			G481<=G11324;
			G486<=G11331;
			G491<=G11332;
			G496<=G11333;
			G501<=G11334;
			G506<=G11335;
			G511<=G11336;
			G516<=G11337;
			G521<=G11330;
			G525<=G11329;
			G530<=G11328;
			G534<=G11327;
			G538<=G11326;
			G542<=G11325;
			G546<=G11043;
			G549<=G11044;
			G552<=G11045;
			G553<=G11046;
			G554<=G11047;
			G557<=G11048;
			G560<=G11049;
			G563<=G11050;
			G566<=G11051;
			G569<=G10876;
			G572<=G10877;
			G575<=G11052;
			G578<=G6286;
			G579<=G6287;
			G580<=G6288;
			G581<=G6289;
			G582<=G6290;
			G583<=G6291;
			G584<=G6292;
			G585<=G6293;
			G586<=G6294;
			G587<=G6295;
			G588<=G6296;
			G589<=G6297;
			G590<=G5653;
			G591<=G9818;
			G599<=G9819;
			G605<=G9820;
			G611<=G9930;
			G617<=G8780;
			G622<=G9338;
			G627<=G5657;
			G630<=G7287;
			G631<=G5654;
			G632<=G5655;
			G635<=G5656;
			G636<=G8781;
			G639<=G8063;
			G643<=G8064;
			G646<=G8065;
			G650<=G8066;
			G654<=G8067;
			G658<=G9339;
			G664<=G8782;
			G668<=G9340;
			G673<=G8428;
			G677<=G9341;
			G682<=G8429;
			G686<=G9342;
			G691<=G8430;
			G695<=G9343;
			G700<=G8431;
			G704<=G9344;
			G709<=G8432;
			G713<=G9345;
			G718<=G8433;
			G722<=G9346;
			G727<=G8434;
			G731<=G9347;
			G736<=G8435;
			G745<=G2639;
			G746<=G2638;
			G754<=G4895;
			G755<=G6298;
			G756<=G755;
			G757<=G11179;
			G758<=G6797;
			G762<=G6798;
			G766<=G6799;
			G770<=G7288;
			G774<=G7785;
			G778<=G8076;
			G782<=G8273;
			G786<=G8436;
			G790<=G8567;
			G794<=G6800;
			G798<=G6801;
			G802<=G6802;
			G806<=G7289;
			G810<=G7786;
			G814<=G8077;
			G818<=G8274;
			G822<=G8437;
			G826<=G8568;
			G829<=G4182;
			G833<=G4183;
			G837<=G4184;
			G841<=G4185;
			G845<=G4186;
			G849<=G4187;
			G853<=G4188;
			G857<=G4189;
			G861<=G4190;
			G865<=G8275;
			G868<=G874;
			G869<=G875;
			G874<=G9821;
			G875<=G9822;
			G876<=G878;
			G878<=G4896;
			G882<=G883;
			G883<=G4897;
			G928<=G8569;
			G932<=G8570;
			G936<=G8571;
			G940<=G8572;
			G944<=G11398;
			G947<=G11399;
			G950<=G11400;
			G953<=G11401;
			G956<=G11402;
			G959<=G11403;
			G962<=G11404;
			G965<=G11405;
			G968<=G11406;
			G971<=G11470;
			G976<=G11471;
			G981<=G11472;
			G986<=G11473;
			G991<=G7802;
			G995<=G7801;
			G999<=G7804;
			G1003<=G7803;
			G1007<=G7806;
			G1011<=G7805;
			G1015<=G7808;
			G1019<=G7807;
			G1023<=G7799;
			G1027<=G7798;
			G1032<=G7800;
			G1035<=G7787;
			G1038<=G7797;
			G1041<=G7788;
			G1044<=G7789;
			G1047<=G7790;
			G1050<=G7791;
			G1053<=G7792;
			G1056<=G7793;
			G1059<=G7794;
			G1062<=G7795;
			G1065<=G7796;
			G1068<=G6803;
			G1071<=G6804;
			G1074<=G6813;
			G1077<=G6805;
			G1080<=G6806;
			G1083<=G6807;
			G1086<=G6808;
			G1089<=G6809;
			G1092<=G6810;
			G1095<=G6811;
			G1098<=G6812;
			G1101<=G6814;
			G1104<=G6815;
			G1107<=G6816;
			G1110<=G6817;
			G1113<=G6313;
			G1117<=G6299;
			G1121<=G6306;
			G1125<=G6307;
			G1129<=G6308;
			G1133<=G6309;
			G1137<=G6310;
			G1141<=G6311;
			G1145<=G6312;
			G1149<=G6305;
			G1153<=G6304;
			G1157<=G6303;
			G1160<=G6302;
			G1163<=G6301;
			G1166<=G6300;
			G1169<=G6314;
			G1206<=G4898;
			G1209<=G10873;
			G1212<=G1217;
			G1215<=G6315;
			G1216<=G1360;
			G1217<=G9823;
			G1218<=G8276;
			G1223<=G8277;
			G1227<=G8278;
			G1231<=G8279;
			G1235<=G7296;
			G1240<=G7297;
			G1245<=G7298;
			G1250<=G7299;
			G1255<=G7300;
			G1260<=G7301;
			G1265<=G7302;
			G1270<=G7303;
			G1275<=G11443;
			G1280<=G7295;
			G1284<=G7294;
			G1289<=G5660;
			G1292<=G7293;
			G1296<=G7292;
			G1300<=G7291;
			G1304<=G7290;
			G1308<=G11627;
			G1311<=G11628;
			G1314<=G11629;
			G1317<=G1356;
			G1318<=G11630;
			G1321<=G11631;
			G1324<=G11632;
			G1327<=G11633;
			G1330<=G11634;
			G1333<=G11635;
			G1336<=G11654;
			G1341<=G11655;
			G1346<=G11656;
			G1351<=G11657;
			G1356<=G6818;
			G1357<=G6330;
			G1360<=G9824;
			G1361<=G1206;
			G1362<=G7305;
			G1365<=G7307;
			G1368<=G7308;
			G1371<=G7311;
			G1374<=G6825;
			G1377<=G7312;
			G1380<=G7314;
			G1383<=G7316;
			G1386<=G7318;
			G1389<=G6836;
			G1393<=G7320;
			G1394<=G7809;
			G1397<=G7322;
			G1400<=G7324;
			G1403<=G8991;
			G1407<=G8993;
			G1411<=G7331;
			G1415<=G7335;
			G1419<=G7332;
			G1424<=G7330;
			G1428<=G8992;
			G1432<=G8990;
			G1436<=G8989;
			G1440<=G8988;
			G1444<=G8987;
			G1448<=G11594;
			G1453<=G7326;
			G1458<=G7327;
			G1462<=G8438;
			G1466<=G8439;
			G1470<=G8440;
			G1474<=G8441;
			G1478<=G8442;
			G1482<=G8443;
			G1486<=G8444;
			G1490<=G8445;
			G1494<=G8446;
			G1499<=G8447;
			G1504<=G7328;
			G1508<=G7329;
			G1512<=G8449;
			G1515<=G7333;
			G1520<=G7334;
			G1524<=G7338;
			G1527<=G4899;
			G1528<=G7339;
			G1531<=G7340;
			G1534<=G7341;
			G1537<=G7342;
			G1540<=G7343;
			G1543<=G7344;
			G1546<=G7345;
			G1549<=G7346;
			G1552<=G7347;
			G1555<=G7348;
			G1558<=G7349;
			G1561<=G7350;
			G1564<=G7351;
			G1567<=G7352;
			G1570<=G4900;
			G1571<=G7353;
			G1574<=G7354;
			G1577<=G7355;
			G1580<=G7356;
			G1583<=G7357;
			G1586<=G7358;
			G1589<=G7359;
			G1592<=G7360;
			G1595<=G7361;
			G1598<=G7362;
			G1601<=G7363;
			G1604<=G7364;
			G1607<=G7365;
			G1610<=G6845;
			G1615<=G8868;
			G1618<=G11611;
			G1621<=G8869;
			G1624<=G8870;
			G1627<=G8871;
			G1630<=G8872;
			G1633<=G8873;
			G1636<=G8874;
			G1639<=G8448;
			G1642<=G11183;
			G1645<=G11184;
			G1648<=G11181;
			G1651<=G11182;
			G1654<=G10874;
			G1657<=G10875;
			G1660<=G11033;
			G1663<=G11034;
			G1666<=G11035;
			G1669<=G11036;
			G1672<=G11037;
			G1675<=G11038;
			G1678<=G11039;
			G1681<=G11040;
			G1684<=G11041;
			G1687<=G11042;
			G1690<=G6844;
			G1703<=G6843;
			G1707<=G4907;
			G1710<=G4901;
			G1711<=G6335;
			G1713<=G6336;
			G1718<=G6337;
			G1721<=G10878;
			G1724<=G10879;
			G1727<=G10880;
			G1730<=G10881;
			G1733<=G10882;
			G1736<=G6846;
			G1737<=G1736;
			G1738<=G5661;
			G1741<=G5662;
			G1744<=G5663;
			G1747<=G5664;
			G1750<=G5665;
			G1753<=G5666;
			G1756<=G5667;
			G1759<=G5668;
			G1762<=G5669;
			G1765<=G3329;
			G1766<=G7810;
			G1771<=G7811;
			G1776<=G7812;
			G1781<=G7813;
			G1786<=G7814;
			G1791<=G8080;
			G1796<=G8280;
			G1801<=G8450;
			G1806<=G8573;
			G1810<=G2044;
			G1811<=G11185;
			G1814<=G9825;
			G1822<=G9826;
			G1828<=G9827;
			G1834<=G9895;
			G1840<=G8694;
			G1845<=G5673;
			G1848<=G7366;
			G1849<=G5670;
			G1850<=G5671;
			G1853<=G5672;
			G1854<=G11408;
			G1857<=G11409;
			G1861<=G7815;
			G1864<=G7816;
			G1868<=G7817;
			G1872<=G9348;
			G1878<=G8695;
			G1882<=G9349;
			G1887<=G8281;
			G1891<=G9350;
			G1896<=G8282;
			G1900<=G9351;
			G1905<=G8283;
			G1909<=G9352;
			G1914<=G8284;
			G1918<=G9353;
			G1923<=G8285;
			G1927<=G9354;
			G1932<=G8286;
			G1936<=G9355;
			G1941<=G8287;
			G1945<=G9356;
			G1950<=G8288;
			G1955<=G6338;
			G1956<=G1955;
			G1957<=G1956;
			G1958<=G6339;
			G1959<=G4217;
		end if;
	end process;
	G22<= not I4777;
	G97<= not I4780;
	G98<= not I4783;
	G110<= not I4786;
	G1962<= not G27;
	G1963<= not G110;
	G1964<= not G114;
	G1965<= not G119;
	G1968<= not G369;
	G1969<= not G456;
	G1972<= not G461;
	G1973<= not G466;
	G1974<= not G627;
	G1975<= not G622;
	G1976<= not G643;
	G1980<= not G646;
	G1981<= not G650;
	G1982<= not G736;
	G1983<= not G750;
	G1984<= not G758;
	G1987<= not G762;
	G1988<= not G766;
	G1989<= not G770;
	G1990<= not G774;
	G1991<= not G778;
	G1992<= not G782;
	G1993<= not G786;
	G1994<= not G794;
	G1997<= not G798;
	G1998<= not G802;
	G1999<= not G806;
	G2000<= not G810;
	G2001<= not G814;
	G2002<= not G818;
	G2003<= not G822;
	G2004<= not I4820;
	G2005<= not G928;
	G2006<= not G932;
	G2007<= not G936;
	G2008<= not G971;
	G2011<= not G976;
	G2012<= not G981;
	G2013<= not G1101;
	G2014<= not G1104;
	G2015<= not G1107;
	G2016<= not G1361;
	G2017<= not G1218;
	G2018<= not G1336;
	G2021<= not G1341;
	G2022<= not G1346;
	G2023<= not G1357;
	G2024<= not G1718;
	G2025<= not G1696;
	G2028<= not G1703;
	G2031<= not G1690;
	G2034<= not G1766;
	G2037<= not G1771;
	G2038<= not G1776;
	G2039<= not G1781;
	G2040<= not G1786;
	G2041<= not G1791;
	G2042<= not G1796;
	G2043<= not G1801;
	G2044<= not I4850;
	G2045<= not G1811;
	G2046<= not G1845;
	G2047<= not G1857;
	G2050<= not G1861;
	G2054<= not G1864;
	G2055<= not G1950;
	G2056<= not I4859;
	G2057<= not G754;
	G2060<= not G1380;
	G2061<= not G1828;
	G2067<= not G108;
	G2068<= not I4866;
	G2069<= not I4869;
	G2070<= not G213;
	G2071<= not I4873;
	G2072<= not I4876;
	G2073<= not I4879;
	G2074<= not G1377;
	G2075<= not I4883;
	G2076<= not I4886;
	G2077<= not G219;
	G2078<= not G135;
	G2079<= not I4891;
	G2080<= not I4894;
	G2082<= not G1371;
	G2083<= not G139;
	G2084<= not I4900;
	G2085<= not I4903;
	G2086<= not I4906;
	G2087<= not G225;
	G2089<= not I4917;
	G2090<= not I4920;
	G2094<= not I4924;
	G2095<= not G143;
	G2097<= not I4935;
	G2098<= not I4938;
	G2100<= not I4948;
	G2101<= not I4951;
	G2103<= not I4961;
	G2108<= not I4992;
	G2110<= not I5002;
	G2112<= not G639;
	G2116<= not I5020;
	G2118<= not G1854;
	G2119<= not I5031;
	G2121<= not I5041;
	G2122<= not I5044;
	G2123<= not I5047;
	G2124<= not I5050;
	G2125<= not I5053;
	G2126<= not G12;
	G2130<= not I5057;
	G2131<= not I5060;
	G2135<= not I5064;
	G2154<= not I5067;
	G2155<= not I5070;
	G2156<= not I5073;
	G2157<= not G1703;
	G2158<= not I5077;
	G2159<= not I5080;
	G2162<= not I5089;
	G2163<= not I5092;
	G2164<= not I5095;
	G2165<= not I5098;
	G2166<= not I5101;
	G2168<= not I5111;
	G2169<= not G42;
	G2170<= not G30;
	G2171<= not I5116;
	G2172<= not G43;
	G2173<= not I5120;
	G2174<= not G31;
	G2175<= not G44;
	G2176<= not G82;
	G2178<= not G45;
	G2179<= not G89;
	G2181<= not I5142;
	G2184<= not G1806;
	G2185<= not G46;
	G2186<= not G90;
	G2187<= not G746;
	G2190<= not I5149;
	G2191<= not G1696;
	G2194<= not G47;
	G2195<= not G83;
	G2196<= not G91;
	G2197<= not G101;
	G2198<= not G668;
	G2199<= not G48;
	G2200<= not G92;
	G2201<= not G102;
	G2202<= not G148;
	G2203<= not G677;
	G2206<= not I5171;
	G2207<= not I5174;
	G2208<= not G84;
	G2209<= not G93;
	G2210<= not G103;
	G2211<= not G153;
	G2212<= not G686;
	G2213<= not G1110;
	G2214<= not G115;
	G2216<= not G41;
	G2217<= not I5192;
	G2218<= not G85;
	G2219<= not G94;
	G2220<= not G104;
	G2221<= not I5198;
	G2222<= not G158;
	G2224<= not G695;
	G2225<= not I5210;
	G2226<= not G86;
	G2227<= not G95;
	G2228<= not G28;
	G2229<= not G162;
	G2230<= not G704;
	G2231<= not I5218;
	G2232<= not I5221;
	G2233<= not I5224;
	G2234<= not G87;
	G2235<= not G96;
	G2237<= not G713;
	G2238<= not I5237;
	G2239<= not I5240;
	G2240<= not G88;
	G2241<= not G722;
	G2242<= not I5245;
	G2243<= not I5248;
	G2244<= not I5251;
	G2245<= not I5254;
	G2246<= not G1810;
	G2247<= not I5258;
	G2248<= not G99;
	G2249<= not G127;
	G2251<= not G731;
	G2252<= not I5271;
	G2253<= not G100;
	G2254<= not G131;
	G2255<= not I5276;
	G2256<= not I5279;
	G2258<= not I5289;
	G2259<= not I5292;
	G2261<= not G1713;
	G2267<= not I5304;
	G2268<= not G654;
	G2269<= not I5308;
	G2270<= not I5311;
	G2271<= not G877;
	G2273<= not G881;
	G2275<= not G757;
	G2296<= not I5332;
	G2297<= not G865;
	G2298<= not I5336;
	G2299<= not G1707;
	G2302<= not G29;
	G2304<= not I5348;
	G2317<= not G622;
	G2320<= not G18;
	G2322<= not I5378;
	G2328<= not G1882;
	G2329<= not I5383;
	G2330<= not G1891;
	G2331<= not G658;
	G2334<= not I5388;
	G2335<= not I5391;
	G2336<= not G1900;
	G2337<= not I5395;
	G2338<= not G1909;
	G2339<= not I5399;
	G2340<= not G1918;
	G2341<= not I5403;
	G2342<= not I5406;
	G2343<= not G1927;
	G2344<= not I5410;
	G2345<= not G1936;
	G2346<= not I5414;
	G2347<= not G1945;
	G2348<= not I5418;
	G2349<= not I5421;
	G2350<= not I5424;
	G2351<= not I5427;
	G2352<= not I5430;
	G2355<= not I5435;
	G2356<= not I5438;
	G2363<= not I5441;
	G2364<= not G611;
	G2368<= not I5445;
	G2369<= not G617;
	G2373<= not G471;
	G2374<= not G591;
	G2381<= not G1368;
	G2382<= not G599;
	G2390<= not I5475;
	G2391<= not I5478;
	G2395<= not G231;
	G2396<= not G1389;
	G2399<= not G605;
	G2406<= not G1365;
	G2407<= not G197;
	G2410<= not G1453;
	G2411<= not I5494;
	G2418<= not I5497;
	G2420<= not G237;
	G2421<= not G1374;
	G2424<= not G1690;
	G2431<= not I5510;
	G2432<= not I5513;
	G2434<= not G1362;
	G2435<= not G201;
	G2436<= not I5525;
	G2438<= not G243;
	G2444<= not G876;
	G2446<= not G1400;
	G2449<= not G790;
	G2450<= not G1351;
	G2451<= not G248;
	G2454<= not I5549;
	G2455<= not G826;
	G2456<= not G1397;
	G2462<= not I5555;
	G2475<= not G192;
	G2479<= not G26;
	G2480<= not I5561;
	G2481<= not G882;
	G2482<= not I5565;
	G2502<= not I5579;
	G2503<= not G1872;
	G2506<= not G636;
	G2507<= not I5584;
	G2508<= not G940;
	G2509<= not I5588;
	G2518<= not G590;
	G2523<= not I5632;
	G2524<= not G986;
	G2529<= not I5638;
	G2530<= not I5641;
	G2537<= not I5646;
	G2539<= not I5652;
	G2540<= not I5655;
	G2541<= not I5658;
	G2542<= not G1868;
	G2543<= not I5662;
	G2547<= not G23;
	G2548<= not I5667;
	G2549<= not G1386;
	G2550<= not G1834;
	G2554<= not I5672;
	G2556<= not G186;
	G2557<= not G1840;
	G2560<= not I5684;
	G2562<= not G1383;
	G2564<= not G1814;
	G2569<= not I5695;
	G2570<= not G207;
	G2571<= not G1822;
	G2578<= not G1962;
	G2579<= not G1969;
	G2586<= not G1972;
	G2593<= not G1973;
	G2601<= not I5704;
	G2602<= not I5707;
	G2603<= not I5710;
	G2604<= not I5713;
	G2605<= not I5716;
	G2606<= not I5719;
	G2607<= not I5722;
	G2608<= not I5725;
	G2609<= not I5728;
	G2610<= not I5731;
	G2611<= not I5734;
	G2612<= not I5737;
	G2613<= not I5740;
	G2614<= not G1994;
	G2617<= not G1997;
	G2620<= not G1998;
	G2623<= not G1999;
	G2626<= not G2000;
	G2629<= not G2001;
	G2632<= not G2002;
	G2635<= not G2003;
	G2638<= not I5751;
	G2639<= not I5754;
	G2640<= not G1984;
	G2641<= not G1987;
	G2642<= not G1988;
	G2643<= not G1989;
	G2644<= not G1990;
	G2645<= not G1991;
	G2646<= not G1992;
	G2647<= not G1993;
	G2648<= not I5765;
	G2649<= not G2005;
	G2650<= not G2006;
	G2651<= not G2007;
	G2652<= not G2008;
	G2653<= not G2011;
	G2654<= not G2012;
	G2655<= not G2013;
	G2662<= not G2014;
	G2669<= not G2015;
	G2677<= not G2034;
	G2683<= not G2037;
	G2689<= not G2038;
	G2695<= not G2039;
	G2701<= not G2040;
	G2707<= not G2041;
	G2713<= not G2042;
	G2719<= not G2043;
	G2725<= not G2018;
	G2726<= not G2021;
	G2727<= not G2022;
	G2728<= not G2025;
	G2731<= not I5789;
	G2732<= not I5792;
	G2733<= not I5795;
	G2742<= not I5798;
	G2743<= not I5801;
	G2745<= not I5809;
	G2748<= not I5812;
	G2749<= not I5815;
	G2750<= not I5818;
	G2751<= not I5821;
	G2752<= not I5824;
	G2753<= not I5827;
	G2754<= not I5830;
	G2755<= not I5833;
	G2757<= not I5837;
	G2758<= not I5840;
	G2759<= not I5843;
	G2763<= not I5847;
	G2764<= not I5850;
	G2765<= not G2184;
	G2771<= not I5854;
	G2772<= not G2508;
	G2773<= not I5858;
	G2774<= not G2276;
	G2775<= not I5862;
	G2777<= not G2276;
	G2778<= not G2276;
	G2779<= not G1974;
	G2789<= not G2276;
	G2790<= not G2276;
	G2793<= not G2276;
	G2796<= not G2276;
	G2797<= not G2524;
	G2798<= not G2449;
	G2799<= not G2276;
	G2801<= not G2117;
	G2802<= not G2276;
	G2803<= not G2154;
	G2808<= not G2156;
	G2809<= not I5909;
	G2812<= not G2158;
	G2813<= not I5913;
	G2814<= not I5916;
	G2817<= not I5919;
	G2818<= not I5922;
	G2819<= not G2159;
	G2820<= not I5926;
	G2821<= not I5929;
	G2824<= not I5932;
	G2825<= not I5935;
	G2826<= not G2163;
	G2827<= not G2164;
	G2828<= not I5940;
	G2829<= not I5943;
	G2832<= not I5946;
	G2833<= not I5949;
	G2834<= not I5952;
	G2837<= not G2130;
	G2838<= not G2165;
	G2839<= not I5957;
	G2840<= not I5960;
	G2843<= not I5963;
	G2844<= not I5966;
	G2845<= not G2168;
	G2846<= not I5970;
	G2847<= not I5973;
	G2850<= not I5976;
	G2851<= not I5979;
	G2852<= not I5982;
	G2853<= not G2171;
	G2854<= not I5986;
	G2855<= not I5989;
	G2858<= not I5992;
	G2859<= not I5995;
	G2860<= not I5998;
	G2861<= not I6001;
	G2864<= not G2298;
	G2867<= not I6007;
	G2868<= not I6010;
	G2871<= not I6013;
	G2872<= not I6016;
	G2873<= not I6019;
	G2874<= not I6022;
	G2877<= not I6025;
	G2880<= not I6028;
	G2881<= not I6031;
	G2882<= not I6034;
	G2883<= not I6037;
	G2884<= not I6040;
	G2885<= not I6043;
	G2888<= not I6046;
	G2889<= not I6049;
	G2890<= not I6052;
	G2891<= not I6055;
	G2896<= not G2356;
	G2902<= not I6061;
	G2903<= not G2166;
	G2904<= not I6065;
	G2905<= not I6068;
	G2906<= not I6071;
	G2907<= not I6074;
	G2908<= not I6077;
	G2909<= not I6080;
	G2912<= not I6085;
	G2913<= not I6088;
	G2914<= not I6091;
	G2915<= not I6094;
	G2916<= not I6097;
	G2919<= not I6102;
	G2920<= not G2462;
	G2937<= not I6106;
	G2941<= not I6118;
	G2942<= not I6121;
	G2946<= not I6133;
	G2949<= not I6150;
	G2952<= not G2455;
	G2955<= not I6156;
	G2956<= not I6159;
	G2958<= not I6163;
	G2960<= not I6173;
	G2962<= not I6183;
	G2964<= not I6193;
	G2965<= not I6196;
	G2971<= not G2046;
	G2980<= not G1983;
	G2985<= not I6217;
	G2986<= not I6220;
	G2989<= not G2135;
	G2991<= not I6233;
	G2994<= not G2057;
	G2997<= not G2135;
	G2998<= not G2462;
	G3007<= not I6240;
	G3009<= not G2135;
	G3012<= not I6247;
	G3037<= not G2135;
	G3038<= not G1982;
	G3039<= not G2310;
	G3040<= not G2135;
	G3044<= not I6256;
	G3050<= not I6260;
	G3051<= not G2135;
	G3052<= not I6264;
	G3055<= not G2135;
	G3060<= not G2135;
	G3066<= not G2135;
	G3067<= not I6273;
	G3068<= not G2303;
	G3069<= not I6277;
	G3076<= not I6282;
	G3077<= not G2213;
	G3086<= not G2276;
	G3088<= not I6294;
	G3092<= not G2181;
	G3093<= not I6299;
	G3094<= not I6302;
	G3095<= not G2482;
	G3096<= not G2482;
	G3097<= not G2482;
	G3102<= not G2482;
	G3103<= not G2391;
	G3105<= not G2482;
	G3109<= not G2482;
	G3110<= not G2482;
	G3112<= not G2482;
	G3113<= not I6343;
	G3119<= not I6347;
	G3121<= not G2462;
	G3138<= not I6356;
	G3141<= not G2563;
	G3142<= not I6360;
	G3143<= not I6363;
	G3144<= not G2462;
	G3161<= not I6367;
	G3164<= not I6370;
	G3186<= not I6373;
	G3206<= not G2055;
	G3207<= not G2439;
	G3208<= not I6381;
	G3212<= not I6385;
	G3213<= not I6388;
	G3214<= not I6391;
	G3219<= not I6395;
	G3220<= not I6398;
	G3226<= not I6403;
	G3227<= not I6406;
	G3228<= not I6409;
	G3246<= not G2482;
	G3252<= not I6414;
	G3253<= not I6417;
	G3254<= not G2322;
	G3255<= not I6421;
	G3256<= not I6424;
	G3260<= not I6428;
	G3262<= not I6432;
	G3266<= not I6436;
	G3267<= not I6439;
	G3271<= not I6443;
	G3272<= not G2450;
	G3274<= not I6454;
	G3290<= not I6461;
	G3291<= not G2161;
	G3292<= not G2373;
	G3305<= not I6474;
	G3306<= not I6477;
	G3307<= not I6480;
	G3318<= not G2245;
	G3321<= not I6484;
	G3323<= not G2157;
	G3326<= not I6495;
	G3327<= not I6498;
	G3328<= not I6501;
	G3329<= not I6504;
	G3330<= not I6507;
	G3331<= not I6510;
	G3332<= not I6513;
	G3333<= not G2779;
	G3334<= not I6517;
	G3335<= not I6520;
	G3336<= not I6523;
	G3337<= not G2745;
	G3343<= not G2779;
	G3344<= not I6528;
	G3345<= not I6531;
	G3348<= not G2733;
	G3351<= not I6535;
	G3352<= not I6538;
	G3353<= not G3121;
	G3359<= not I6543;
	G3362<= not I6546;
	G3363<= not I6549;
	G3364<= not G3121;
	G3365<= not I6553;
	G3368<= not G3138;
	G3369<= not I6557;
	G3370<= not I6560;
	G3371<= not G2837;
	G3372<= not G3121;
	G3373<= not I6565;
	G3375<= not I6569;
	G3378<= not I6572;
	G3379<= not G3121;
	G3380<= not I6576;
	G3382<= not I6580;
	G3384<= not G3143;
	G3385<= not G3121;
	G3386<= not G3144;
	G3387<= not I6587;
	G3388<= not I6590;
	G3390<= not G3161;
	G3391<= not G2896;
	G3392<= not G3121;
	G3393<= not G3144;
	G3394<= not I6598;
	G3395<= not I6601;
	G3397<= not G2896;
	G3398<= not G2896;
	G3404<= not G3121;
	G3405<= not G3144;
	G3406<= not I6611;
	G3408<= not G3108;
	G3411<= not I6616;
	G3413<= not G2896;
	G3415<= not G3121;
	G3416<= not G3144;
	G3417<= not I6624;
	G3419<= not G3104;
	G3424<= not G2896;
	G3426<= not G3121;
	G3427<= not G3144;
	G3428<= not I6639;
	G3430<= not I6643;
	G3432<= not G3144;
	G3433<= not I6648;
	G3436<= not G3144;
	G3437<= not I6654;
	G3439<= not G3144;
	G3440<= not G3041;
	G3458<= not G3144;
	G3459<= not I6661;
	G3461<= not I6671;
	G3463<= not G3256;
	G3473<= not I6676;
	G3474<= not I6679;
	G3475<= not G3056;
	G3479<= not G2655;
	G3485<= not G2662;
	G3491<= not G2669;
	G3496<= not I6686;
	G3500<= not I6690;
	G3501<= not G3077;
	G3505<= not I6694;
	G3507<= not G3307;
	G3517<= not I6702;
	G3518<= not G3164;
	G3519<= not G3164;
	G3520<= not G2779;
	G3521<= not G3164;
	G3522<= not G3164;
	G3523<= not G2971;
	G3528<= not G3164;
	G3531<= not G2971;
	G3532<= not G3164;
	G3537<= not G3164;
	G3538<= not I6726;
	G3539<= not G3015;
	G3540<= not G3307;
	G3543<= not G3101;
	G3544<= not G3164;
	G3545<= not I6733;
	G3546<= not G3307;
	G3566<= not I6738;
	G3582<= not G3164;
	G3583<= not I6742;
	G3621<= not I6754;
	G3622<= not I6757;
	G3624<= not I6767;
	G3627<= not I6784;
	G3628<= not G3111;
	G3629<= not G3228;
	G3630<= not I6789;
	G3632<= not I6799;
	G3633<= not I6802;
	G3635<= not I6812;
	G3636<= not I6815;
	G3637<= not I6818;
	G3638<= not I6821;
	G3663<= not I6832;
	G3664<= not G3209;
	G3682<= not G2920;
	G3683<= not I6844;
	G3693<= not G2920;
	G3694<= not I6851;
	G3697<= not I6856;
	G3703<= not G2920;
	G3704<= not I6861;
	G3705<= not G3113;
	G3707<= not G2920;
	G3708<= not I6867;
	G3709<= not I6870;
	G3710<= not G3215;
	G3715<= not G2920;
	G3716<= not I6876;
	G3719<= not G2920;
	G3720<= not I6888;
	G3721<= not I6891;
	G3722<= not I6894;
	G3723<= not G3071;
	G3726<= not I6898;
	G3727<= not I6901;
	G3728<= not I6904;
	G3729<= not I6907;
	G3730<= not G3015;
	G3731<= not I6911;
	G3732<= not I6914;
	G3733<= not I6917;
	G3735<= not I6921;
	G3736<= not I6924;
	G3737<= not G2834;
	G3738<= not G3062;
	G3742<= not I6929;
	G3743<= not I6932;
	G3744<= not G3307;
	G3747<= not G3015;
	G3748<= not G2971;
	G3749<= not I6938;
	G3750<= not I6941;
	G3751<= not I6944;
	G3752<= not I6947;
	G3756<= not G3015;
	G3757<= not I6952;
	G3758<= not I6955;
	G3759<= not I6958;
	G3760<= not G3003;
	G3761<= not I6962;
	G3762<= not I6965;
	G3763<= not I6968;
	G3764<= not I6971;
	G3765<= not G3120;
	G3767<= not I6976;
	G3768<= not I6979;
	G3769<= not I6982;
	G3770<= not I6985;
	G3773<= not I6996;
	G3774<= not I6999;
	G3775<= not I7002;
	G3776<= not G2579;
	G3782<= not I7006;
	G3783<= not I7009;
	G3784<= not G2586;
	G3790<= not G3228;
	G3791<= not I7014;
	G3792<= not I7017;
	G3793<= not G2593;
	G3798<= not G3228;
	G3799<= not I7022;
	G3800<= not G3292;
	G3810<= not G3228;
	G3811<= not I7029;
	G3812<= not G3228;
	G3814<= not G3228;
	G3815<= not G3228;
	G3816<= not G3228;
	G3817<= not I7043;
	G3820<= not I7048;
	G3828<= not G2920;
	G3861<= not I7054;
	G3862<= not G2920;
	G3874<= not G2920;
	G3876<= not I7061;
	G3877<= not I7064;
	G3878<= not G2920;
	G3903<= not I7070;
	G3905<= not G2920;
	G3906<= not G3015;
	G3907<= not I7076;
	G3909<= not G2920;
	G3910<= not G3015;
	G3911<= not G3015;
	G3913<= not G2920;
	G3914<= not G3015;
	G3937<= not I7086;
	G3938<= not G2991;
	G3940<= not G2920;
	G3941<= not G3015;
	G3943<= not G2779;
	G3944<= not G2920;
	G3945<= not I7096;
	G3946<= not I7099;
	G3967<= not G3247;
	G3971<= not I7104;
	G3975<= not G3121;
	G3976<= not I7109;
	G3977<= not I7112;
	G3980<= not G3121;
	G3981<= not I7118;
	G3982<= not G3052;
	G3983<= not G3222;
	G3988<= not G3121;
	G3990<= not G3121;
	G3995<= not G3121;
	G3996<= not G3144;
	G3997<= not I7131;
	G4001<= not G3200;
	G4002<= not G3121;
	G4003<= not G3144;
	G4004<= not I7140;
	G4005<= not I7143;
	G4010<= not G3144;
	G4011<= not I7151;
	G4012<= not I7154;
	G4013<= not I7157;
	G4049<= not G3144;
	G4050<= not I7163;
	G4051<= not I7166;
	G4055<= not G3144;
	G4056<= not I7173;
	G4057<= not I7176;
	G4060<= not G3144;
	G4061<= not I7182;
	G4062<= not I7185;
	G4065<= not G2794;
	G4066<= not I7191;
	G4067<= not I7194;
	G4077<= not I7202;
	G4078<= not I7205;
	G4080<= not G2903;
	G4081<= not I7210;
	G4082<= not I7213;
	G4083<= not I7216;
	G4084<= not G3119;
	G4087<= not I7220;
	G4093<= not G2965;
	G4094<= not G2744;
	G4095<= not I7233;
	G4096<= not I7236;
	G4098<= not I7240;
	G4102<= not I7244;
	G4105<= not I7249;
	G4112<= not G2994;
	G4113<= not I7255;
	G4116<= not I7260;
	G4121<= not I7264;
	G4124<= not I7269;
	G4125<= not I7272;
	G4127<= not I7276;
	G4129<= not I7280;
	G4140<= not I7284;
	G4142<= not I7288;
	G4143<= not I7291;
	G4156<= not I7295;
	G4158<= not G3304;
	G4159<= not I7300;
	G4160<= not I7303;
	G4163<= not I7308;
	G4164<= not I7311;
	G4165<= not G3164;
	G4166<= not I7315;
	G4167<= not I7318;
	G4170<= not G3328;
	G4171<= not I7330;
	G4172<= not I7333;
	G4173<= not I7336;
	G4174<= not I7339;
	G4175<= not I7342;
	G4176<= not I7345;
	G4177<= not I7348;
	G4178<= not I7351;
	G4179<= not I7354;
	G4180<= not I7357;
	G4181<= not I7360;
	G4182<= not I7363;
	G4183<= not I7366;
	G4184<= not I7369;
	G4185<= not I7372;
	G4186<= not I7375;
	G4187<= not I7378;
	G4188<= not I7381;
	G4189<= not I7384;
	G4190<= not I7387;
	G4191<= not I7390;
	G4192<= not I7393;
	G4193<= not I7396;
	G4194<= not I7399;
	G4195<= not I7402;
	G4196<= not I7405;
	G4197<= not I7408;
	G4198<= not I7411;
	G4199<= not I7414;
	G4200<= not I7417;
	G4201<= not I7420;
	G4202<= not I7423;
	G4203<= not I7426;
	G4204<= not I7429;
	G4205<= not I7432;
	G4206<= not I7435;
	G4207<= not I7438;
	G4208<= not I7441;
	G4209<= not I7444;
	G4210<= not I7447;
	G4211<= not I7450;
	G4212<= not I7453;
	G4213<= not I7456;
	G4214<= not I7459;
	G4215<= not I7462;
	G4216<= not I7465;
	G4217<= not I7468;
	G4219<= not G3635;
	G4221<= not G3914;
	G4222<= not G3638;
	G4225<= not I7478;
	G4226<= not G3698;
	G4228<= not G3914;
	G4232<= not I7487;
	G4233<= not G3698;
	G4237<= not G4013;
	G4240<= not G3664;
	G4241<= not G3664;
	G4242<= not G3664;
	G4243<= not G3524;
	G4250<= not G3698;
	G4254<= not G4013;
	G4256<= not G3664;
	G4257<= not G3664;
	G4258<= not I7509;
	G4260<= not I7513;
	G4262<= not G4013;
	G4263<= not G3586;
	G4265<= not G3664;
	G4266<= not G3688;
	G4268<= not I7523;
	G4270<= not G4013;
	G4271<= not G3971;
	G4272<= not G3586;
	G4273<= not G4013;
	G4275<= not G3664;
	G4277<= not G3688;
	G4279<= not I7536;
	G4280<= not G4013;
	G4281<= not G3586;
	G4282<= not G4013;
	G4284<= not G3664;
	G4285<= not G3688;
	G4287<= not I7546;
	G4288<= not G4130;
	G4289<= not G4013;
	G4290<= not G3586;
	G4291<= not G4013;
	G4292<= not G3863;
	G4294<= not G3664;
	G4295<= not I7556;
	G4296<= not I7559;
	G4298<= not G4130;
	G4299<= not G4144;
	G4305<= not G4013;
	G4306<= not G3586;
	G4307<= not G4013;
	G4308<= not G3863;
	G4310<= not I7577;
	G4311<= not G4130;
	G4312<= not G4144;
	G4313<= not G3586;
	G4314<= not G4013;
	G4315<= not G3863;
	G4317<= not I7586;
	G4318<= not G4130;
	G4319<= not G4144;
	G4320<= not G4013;
	G4321<= not G3863;
	G4322<= not I7593;
	G4323<= not G4130;
	G4324<= not G4144;
	G4326<= not G3863;
	G4327<= not I7600;
	G4328<= not G4130;
	G4329<= not G4144;
	G4331<= not I7606;
	G4332<= not G4130;
	G4333<= not G4144;
	G4335<= not I7612;
	G4336<= not G4130;
	G4337<= not G4144;
	G4339<= not G4144;
	G4344<= not G3946;
	G4346<= not I7625;
	G4347<= not G3880;
	G4351<= not I7630;
	G4352<= not I7633;
	G4353<= not I7636;
	G4354<= not I7639;
	G4355<= not I7642;
	G4359<= not G3880;
	G4361<= not I7648;
	G4362<= not I7651;
	G4363<= not I7654;
	G4365<= not G3880;
	G4366<= not I7659;
	G4367<= not I7662;
	G4368<= not I7665;
	G4369<= not I7668;
	G4370<= not I7671;
	G4371<= not I7674;
	G4372<= not I7677;
	G4373<= not I7680;
	G4375<= not G3638;
	G4376<= not I7691;
	G4377<= not I7694;
	G4378<= not I7697;
	G4379<= not G3698;
	G4380<= not I7701;
	G4381<= not G3914;
	G4382<= not G3638;
	G4384<= not I7707;
	G4385<= not I7710;
	G4386<= not I7713;
	G4387<= not I7716;
	G4388<= not I7719;
	G4390<= not G3914;
	G4391<= not G3638;
	G4393<= not I7726;
	G4394<= not I7729;
	G4395<= not I7732;
	G4396<= not I7735;
	G4398<= not G3914;
	G4399<= not G3638;
	G4411<= not I7743;
	G4412<= not I7746;
	G4413<= not I7749;
	G4414<= not I7752;
	G4415<= not G3914;
	G4416<= not G3638;
	G4417<= not I7757;
	G4418<= not I7760;
	G4419<= not I7763;
	G4420<= not I7766;
	G4424<= not G3688;
	G4425<= not I7771;
	G4426<= not G3914;
	G4427<= not G3638;
	G4428<= not I7776;
	G4429<= not I7779;
	G4430<= not I7782;
	G4435<= not G3914;
	G4436<= not G3638;
	G4437<= not G3345;
	G4438<= not I7790;
	G4439<= not I7793;
	G4440<= not G4130;
	G4441<= not G3914;
	G4442<= not G3638;
	G4443<= not G3359;
	G4444<= not I7800;
	G4445<= not I7803;
	G4449<= not G4144;
	G4450<= not G3914;
	G4451<= not G3638;
	G4452<= not G3365;
	G4453<= not I7810;
	G4454<= not G3914;
	G4456<= not G3375;
	G4457<= not G3829;
	G4458<= not I7817;
	G4459<= not I7820;
	G4460<= not G3820;
	G4461<= not G3829;
	G4462<= not I7825;
	G4463<= not G3829;
	G4464<= not I7829;
	G4466<= not I7833;
	G4467<= not G3829;
	G4468<= not I7837;
	G4469<= not I7840;
	G4470<= not I7843;
	G4472<= not I7847;
	G4474<= not G3820;
	G4475<= not I7852;
	G4478<= not G3820;
	G4479<= not I7858;
	G4485<= not G3546;
	G4491<= not G3546;
	G4495<= not I7886;
	G4496<= not I7889;
	G4499<= not G3546;
	G4501<= not G3946;
	G4504<= not I7899;
	G4507<= not G3546;
	G4508<= not G3946;
	G4509<= not I7906;
	G4510<= not I7909;
	G4511<= not G3586;
	G4513<= not G3546;
	G4514<= not G3946;
	G4515<= not I7916;
	G4519<= not I7920;
	G4520<= not I7923;
	G4521<= not G3586;
	G4523<= not G3546;
	G4524<= not G3946;
	G4525<= not G3880;
	G4526<= not I7931;
	G4530<= not I7935;
	G4533<= not I7938;
	G4535<= not G3946;
	G4536<= not G3880;
	G4541<= not I7946;
	G4543<= not G3946;
	G4544<= not G3880;
	G4545<= not I7952;
	G4549<= not I7956;
	G4551<= not G3946;
	G4552<= not G3880;
	G4555<= not I7964;
	G4557<= not G3946;
	G4558<= not G3880;
	G4562<= not I7973;
	G4563<= not G3946;
	G4564<= not G3880;
	G4566<= not G3753;
	G4567<= not G3374;
	G4575<= not G3880;
	G4577<= not I7984;
	G4580<= not G3880;
	G4583<= not G3880;
	G4586<= not G4089;
	G4587<= not G3829;
	G4589<= not I7996;
	G4590<= not I7999;
	G4591<= not G3829;
	G4592<= not G3829;
	G4593<= not I8004;
	G4596<= not I8007;
	G4602<= not I8011;
	G4603<= not G3829;
	G4606<= not G3829;
	G4608<= not G3829;
	G4614<= not G3829;
	G4615<= not I8024;
	G4618<= not G3829;
	G4620<= not I8031;
	G4631<= not G3820;
	G4636<= not I8036;
	G4637<= not I8039;
	G4638<= not G3354;
	G4669<= not G4013;
	G4671<= not G3354;
	G4673<= not G4013;
	G4674<= not I8050;
	G4676<= not G3354;
	G4678<= not G3546;
	G4679<= not G4013;
	G4680<= not G3829;
	G4681<= not G3546;
	G4711<= not I8061;
	G4713<= not G3546;
	G4716<= not G3546;
	G4717<= not G3829;
	G4719<= not G3586;
	G4721<= not G3546;
	G4724<= not G3586;
	G4726<= not G3546;
	G4728<= not I8080;
	G4729<= not G3586;
	G4730<= not G3546;
	G4731<= not I8085;
	G4733<= not I8089;
	G4734<= not G3586;
	G4735<= not G3546;
	G4737<= not G3440;
	G4738<= not G3440;
	G4739<= not G4117;
	G4746<= not I8098;
	G4747<= not G3586;
	G4748<= not G3546;
	G4754<= not G3440;
	G4755<= not G3440;
	G4756<= not G3440;
	G4757<= not I8109;
	G4758<= not G3586;
	G4761<= not G3440;
	G4762<= not I8116;
	G4763<= not G3586;
	G4766<= not G3440;
	G4767<= not I8123;
	G4768<= not I8126;
	G4769<= not G3586;
	G4772<= not G3440;
	G4773<= not I8133;
	G4774<= not I8136;
	G4775<= not I8139;
	G4776<= not G3586;
	G4777<= not G3992;
	G4780<= not G3440;
	G4781<= not I8147;
	G4782<= not G4089;
	G4783<= not G3829;
	G4785<= not G3337;
	G4786<= not I8154;
	G4787<= not G3423;
	G4789<= not G3337;
	G4790<= not G3337;
	G4791<= not I8161;
	G4794<= not I8164;
	G4802<= not G3337;
	G4805<= not G3337;
	G4811<= not G3661;
	G4819<= not G3354;
	G4822<= not G3706;
	G4835<= not I8192;
	G4840<= not I8199;
	G4867<= not I8204;
	G4872<= not I8211;
	G4874<= not I8215;
	G4880<= not G3638;
	G4885<= not I8228;
	G4886<= not I8231;
	G4887<= not I8234;
	G4888<= not I8237;
	G4889<= not I8240;
	G4894<= not I8247;
	G4895<= not I8250;
	G4896<= not I8253;
	G4897<= not I8256;
	G4898<= not I8259;
	G4899<= not I8262;
	G4900<= not I8265;
	G4901<= not I8268;
	G4906<= not I8275;
	G4907<= not I8278;
	G4908<= not G4396;
	G4912<= not I8282;
	G4913<= not I8285;
	G4915<= not G4413;
	G4919<= not I8290;
	G4920<= not I8293;
	G4933<= not I8298;
	G4934<= not G4243;
	G4935<= not G4420;
	G4939<= not I8303;
	G4942<= not I8308;
	G4943<= not I8311;
	G4944<= not G4430;
	G4948<= not I8315;
	G4951<= not I8320;
	G4953<= not I8324;
	G4954<= not G4509;
	G4958<= not I8328;
	G4961<= not I8333;
	G4963<= not I8337;
	G4966<= not I8340;
	G4970<= not G4411;
	G4975<= not I8351;
	G4988<= not I8358;
	G5007<= not I8379;
	G5011<= not I8385;
	G5012<= not I8388;
	G5027<= not I8396;
	G5032<= not I8403;
	G5033<= not I8406;
	G5035<= not I8410;
	G5037<= not I8414;
	G5039<= not I8418;
	G5040<= not I8421;
	G5042<= not G4840;
	G5043<= not G4840;
	G5047<= not G4354;
	G5050<= not I8429;
	G5052<= not G4394;
	G5062<= not G4840;
	G5063<= not G4363;
	G5066<= not I8436;
	G5068<= not G4840;
	G5069<= not G4368;
	G5072<= not I8442;
	G5073<= not G4840;
	G5075<= not G4439;
	G5078<= not G4372;
	G5081<= not I8449;
	G5082<= not G4840;
	G5085<= not G4377;
	G5088<= not I8456;
	G5089<= not G4840;
	G5091<= not G4385;
	G5094<= not I8462;
	G5095<= not I8465;
	G5096<= not G4840;
	G5098<= not G4840;
	G5101<= not I8473;
	G5102<= not I8476;
	G5105<= not I8487;
	G5106<= not I8490;
	G5107<= not G4459;
	G5109<= not I8495;
	G5111<= not I8499;
	G5112<= not G4682;
	G5113<= not I8503;
	G5114<= not I8506;
	G5116<= not G4682;
	G5117<= not G4682;
	G5120<= not I8520;
	G5121<= not G4682;
	G5122<= not G4682;
	G5124<= not G4596;
	G5127<= not I8535;
	G5143<= not G4682;
	G5144<= not G4682;
	G5146<= not G4596;
	G5149<= not I8551;
	G5166<= not G4682;
	G5167<= not G4682;
	G5169<= not G4596;
	G5175<= not G4682;
	G5176<= not G4682;
	G5177<= not G4596;
	G5183<= not G4640;
	G5184<= not G4682;
	G5185<= not G4682;
	G5191<= not G4640;
	G5192<= not G4640;
	G5193<= not G4682;
	G5195<= not G4453;
	G5197<= not I8611;
	G5198<= not I8614;
	G5200<= not G4567;
	G5202<= not G4640;
	G5203<= not G4640;
	G5205<= not G4366;
	G5210<= not I8631;
	G5213<= not G4640;
	G5214<= not G4640;
	G5216<= not G4445;
	G5218<= not I8647;
	G5222<= not G4640;
	G5223<= not G4640;
	G5231<= not G4640;
	G5232<= not G4640;
	G5236<= not G4361;
	G5241<= not G4386;
	G5245<= not G4369;
	G5251<= not G4640;
	G5252<= not G4640;
	G5253<= not G4346;
	G5261<= not G4640;
	G5262<= not G4353;
	G5265<= not G4362;
	G5267<= not I8711;
	G5270<= not G4367;
	G5272<= not I8724;
	G5275<= not G4371;
	G5281<= not G4428;
	G5284<= not G4376;
	G5285<= not G4355;
	G5288<= not G4438;
	G5291<= not G4384;
	G5292<= not G4445;
	G5296<= not G4444;
	G5299<= not G4393;
	G5301<= not G4373;
	G5305<= not G4378;
	G5314<= not G4387;
	G5320<= not G4418;
	G5344<= not I8811;
	G5348<= not I8815;
	G5353<= not I8820;
	G5391<= not I8827;
	G5395<= not I8831;
	G5397<= not I8835;
	G5401<= not I8839;
	G5402<= not I8842;
	G5415<= not I8848;
	G5416<= not I8851;
	G5417<= not I8854;
	G5419<= not I8858;
	G5420<= not G4300;
	G5422<= not G4470;
	G5423<= not G4300;
	G5424<= not I8865;
	G5425<= not G4300;
	G5426<= not I8869;
	G5443<= not I8872;
	G5446<= not I8877;
	G5469<= not I8880;
	G5471<= not G4370;
	G5472<= not I8885;
	G5474<= not I8889;
	G5475<= not I8892;
	G5481<= not I8900;
	G5482<= not I8903;
	G5486<= not G4395;
	G5490<= not I8911;
	G5494<= not G4412;
	G5498<= not I8919;
	G5503<= not G4515;
	G5504<= not G4419;
	G5508<= not I8929;
	G5509<= not G4739;
	G5511<= not I8934;
	G5515<= not G4429;
	G5519<= not G4811;
	G5520<= not I8943;
	G5521<= not G4530;
	G5534<= not G4545;
	G5542<= not I8967;
	G5546<= not I8973;
	G5567<= not I8982;
	G5568<= not I8985;
	G5572<= not I8989;
	G5574<= not G4300;
	G5586<= not I8996;
	G5589<= not I9001;
	G5593<= not I9013;
	G5594<= not I9016;
	G5596<= not I9020;
	G5597<= not I9023;
	G5603<= not I9029;
	G5604<= not I9032;
	G5613<= not G4840;
	G5614<= not I9040;
	G5615<= not I9043;
	G5616<= not I9046;
	G5619<= not G4840;
	G5620<= not G4417;
	G5623<= not I9053;
	G5624<= not I9056;
	G5627<= not G4840;
	G5628<= not I9062;
	G5629<= not I9065;
	G5630<= not I9068;
	G5633<= not G4388;
	G5637<= not I9074;
	G5638<= not I9077;
	G5639<= not I9080;
	G5641<= not I9084;
	G5642<= not I9087;
	G5643<= not I9090;
	G5644<= not I9093;
	G5645<= not I9096;
	G5646<= not I9099;
	G5647<= not I9102;
	G5648<= not I9105;
	G5649<= not I9108;
	G5650<= not I9111;
	G5651<= not I9114;
	G5652<= not I9117;
	G5653<= not I9120;
	G5654<= not I9123;
	G5655<= not I9126;
	G5656<= not I9129;
	G5657<= not I9132;
	G5658<= not I9135;
	G5659<= not I9138;
	G5660<= not I9141;
	G5661<= not I9144;
	G5662<= not I9147;
	G5663<= not I9150;
	G5664<= not I9153;
	G5665<= not I9156;
	G5666<= not I9159;
	G5667<= not I9162;
	G5668<= not I9165;
	G5669<= not I9168;
	G5670<= not I9171;
	G5671<= not I9174;
	G5672<= not I9177;
	G5673<= not I9180;
	G5676<= not I9185;
	G5677<= not I9188;
	G5678<= not I9191;
	G5679<= not I9194;
	G5682<= not I9199;
	G5683<= not I9202;
	G5684<= not I9205;
	G5685<= not I9208;
	G5688<= not I9213;
	G5689<= not I9216;
	G5691<= not G5236;
	G5692<= not I9221;
	G5693<= not I9224;
	G5696<= not I9229;
	G5697<= not I9232;
	G5700<= not I9237;
	G5701<= not I9240;
	G5702<= not I9243;
	G5705<= not I9248;
	G5708<= not I9253;
	G5718<= not I9256;
	G5719<= not I9259;
	G5723<= not I9265;
	G5724<= not I9268;
	G5727<= not I9273;
	G5728<= not I9276;
	G5729<= not I9279;
	G5730<= not I9282;
	G5733<= not I9287;
	G5734<= not I9290;
	G5735<= not I9293;
	G5736<= not I9296;
	G5740<= not I9302;
	G5741<= not I9305;
	G5742<= not I9308;
	G5743<= not I9311;
	G5747<= not I9317;
	G5748<= not I9320;
	G5751<= not I9323;
	G5752<= not I9326;
	G5753<= not I9329;
	G5754<= not I9332;
	G5758<= not I9338;
	G5759<= not I9341;
	G5766<= not I9346;
	G5767<= not I9349;
	G5768<= not I9352;
	G5773<= not I9359;
	G5774<= not I9362;
	G5777<= not I9365;
	G5778<= not I9368;
	G5779<= not I9371;
	G5783<= not I9377;
	G5784<= not I9380;
	G5787<= not I9383;
	G5790<= not I9388;
	G5791<= not I9391;
	G5794<= not I9394;
	G5797<= not I9399;
	G5800<= not I9402;
	G5801<= not G5320;
	G5805<= not I9409;
	G5808<= not G5320;
	G5811<= not I9415;
	G5812<= not G5320;
	G5815<= not I9421;
	G5816<= not I9424;
	G5817<= not I9427;
	G5818<= not G5320;
	G5821<= not I9433;
	G5822<= not G5320;
	G5826<= not I9440;
	G5827<= not I9443;
	G5830<= not I9446;
	G5836<= not G5320;
	G5839<= not I9452;
	G5840<= not G5320;
	G5843<= not I9458;
	G5844<= not I9461;
	G5845<= not G5320;
	G5850<= not G5320;
	G5856<= not G5245;
	G5858<= not I9475;
	G5862<= not I9479;
	G5864<= not I9483;
	G5865<= not I9486;
	G5866<= not G5361;
	G5874<= not I9491;
	G5875<= not G5361;
	G5876<= not G5361;
	G5878<= not G5309;
	G5879<= not I9498;
	G5880<= not G5361;
	G5881<= not G5361;
	G5883<= not G5309;
	G5884<= not I9505;
	G5885<= not G5361;
	G5886<= not G5361;
	G5887<= not I9510;
	G5888<= not G5102;
	G5889<= not I9514;
	G5890<= not G5361;
	G5891<= not G5361;
	G5892<= not I9519;
	G5893<= not G5106;
	G5894<= not G5361;
	G5895<= not G5361;
	G5896<= not I9525;
	G5898<= not G5361;
	G5899<= not G5361;
	G5900<= not I9531;
	G5901<= not G5361;
	G5903<= not I9536;
	G5904<= not I9539;
	G5912<= not I9544;
	G5916<= not I9550;
	G5936<= not I9564;
	G5937<= not I9567;
	G5941<= not I9571;
	G5943<= not I9581;
	G5947<= not I9585;
	G5948<= not I9588;
	G5949<= not I9591;
	G5980<= not I9594;
	G5982<= not I9598;
	G5984<= not I9602;
	G5987<= not I9605;
	G5992<= not I9608;
	G5994<= not I9612;
	G5997<= not I9617;
	G5998<= not I9620;
	G6001<= not I9625;
	G6014<= not G5309;
	G6016<= not I9632;
	G6030<= not I9639;
	G6031<= not I9642;
	G6036<= not I9647;
	G6039<= not I9652;
	G6040<= not I9655;
	G6041<= not I9658;
	G6043<= not I9662;
	G6044<= not I9665;
	G6046<= not I9669;
	G6048<= not I9673;
	G6050<= not I9677;
	G6051<= not I9680;
	G6052<= not G5426;
	G6053<= not I9684;
	G6055<= not I9688;
	G6056<= not G5426;
	G6057<= not G5446;
	G6060<= not I9695;
	G6062<= not I9699;
	G6063<= not G5446;
	G6069<= not I9706;
	G6072<= not G4977;
	G6073<= not I9712;
	G6076<= not I9717;
	G6077<= not I9720;
	G6081<= not G4977;
	G6082<= not I9727;
	G6084<= not I9731;
	G6085<= not I9734;
	G6086<= not I9737;
	G6089<= not G4977;
	G6091<= not I9744;
	G6094<= not I9749;
	G6097<= not I9754;
	G6100<= not I9759;
	G6101<= not I9762;
	G6103<= not I9766;
	G6104<= not I9769;
	G6106<= not I9773;
	G6107<= not I9776;
	G6108<= not I9779;
	G6109<= not G5052;
	G6110<= not I9783;
	G6111<= not I9786;
	G6112<= not I9789;
	G6113<= not I9792;
	G6114<= not I9795;
	G6115<= not I9798;
	G6116<= not I9801;
	G6117<= not I9804;
	G6118<= not I9807;
	G6119<= not I9810;
	G6120<= not I9813;
	G6121<= not I9816;
	G6125<= not I9822;
	G6127<= not I9826;
	G6128<= not I9829;
	G6131<= not G5548;
	G6132<= not I9833;
	G6133<= not I9836;
	G6134<= not I9839;
	G6135<= not I9842;
	G6136<= not I9845;
	G6137<= not I9848;
	G6140<= not I9851;
	G6141<= not I9854;
	G6144<= not I9857;
	G6145<= not I9860;
	G6146<= not I9863;
	G6149<= not I9866;
	G6150<= not I9869;
	G6151<= not I9872;
	G6154<= not I9875;
	G6156<= not G5426;
	G6157<= not I9880;
	G6158<= not I9883;
	G6161<= not I9886;
	G6164<= not G5426;
	G6165<= not G5446;
	G6166<= not I9893;
	G6169<= not I9896;
	G6170<= not G5426;
	G6171<= not G5446;
	G6172<= not I9901;
	G6175<= not G5320;
	G6176<= not I9905;
	G6178<= not G4977;
	G6181<= not G5426;
	G6182<= not G5446;
	G6183<= not G5320;
	G6184<= not I9915;
	G6190<= not G5426;
	G6191<= not G5446;
	G6192<= not I9923;
	G6195<= not G5426;
	G6196<= not G5446;
	G6197<= not I9930;
	G6200<= not I9935;
	G6201<= not I9938;
	G6202<= not G5426;
	G6203<= not G5446;
	G6208<= not I9953;
	G6209<= not I9956;
	G6210<= not G5205;
	G6213<= not G5426;
	G6214<= not G5446;
	G6218<= not I9965;
	G6219<= not G5426;
	G6220<= not G5446;
	G6226<= not I9973;
	G6227<= not G5446;
	G6236<= not I9981;
	G6237<= not I9984;
	G6239<= not I9988;
	G6241<= not I9992;
	G6242<= not I9995;
	G6248<= not I10003;
	G6249<= not I10006;
	G6250<= not I10009;
	G6251<= not I10012;
	G6252<= not I10015;
	G6253<= not I10018;
	G6254<= not I10021;
	G6255<= not I10024;
	G6256<= not I10027;
	G6257<= not I10030;
	G6258<= not I10033;
	G6259<= not I10036;
	G6260<= not I10039;
	G6261<= not I10042;
	G6262<= not I10045;
	G6263<= not I10048;
	G6264<= not I10051;
	G6265<= not I10054;
	G6266<= not I10057;
	G6267<= not I10060;
	G6268<= not I10063;
	G6269<= not I10066;
	G6270<= not I10069;
	G6271<= not I10072;
	G6272<= not I10075;
	G6273<= not I10078;
	G6274<= not I10081;
	G6275<= not I10084;
	G6276<= not I10087;
	G6277<= not I10090;
	G6278<= not I10093;
	G6279<= not I10096;
	G6280<= not I10099;
	G6281<= not I10102;
	G6282<= not I10105;
	G6283<= not I10108;
	G6284<= not I10111;
	G6285<= not I10114;
	G6286<= not I10117;
	G6287<= not I10120;
	G6288<= not I10123;
	G6289<= not I10126;
	G6290<= not I10129;
	G6291<= not I10132;
	G6292<= not I10135;
	G6293<= not I10138;
	G6294<= not I10141;
	G6295<= not I10144;
	G6296<= not I10147;
	G6297<= not I10150;
	G6298<= not I10153;
	G6299<= not I10156;
	G6300<= not I10159;
	G6301<= not I10162;
	G6302<= not I10165;
	G6303<= not I10168;
	G6304<= not I10171;
	G6305<= not I10174;
	G6306<= not I10177;
	G6307<= not I10180;
	G6308<= not I10183;
	G6309<= not I10186;
	G6310<= not I10189;
	G6311<= not I10192;
	G6312<= not I10195;
	G6313<= not I10198;
	G6314<= not I10201;
	G6315<= not I10204;
	G6330<= not I10221;
	G6335<= not I10228;
	G6336<= not I10231;
	G6337<= not I10234;
	G6338<= not I10237;
	G6339<= not I10240;
	G6340<= not I10243;
	G6343<= not I10248;
	G6344<= not I10251;
	G6349<= not I10258;
	G6354<= not G5867;
	G6361<= not G5867;
	G6365<= not I10274;
	G6368<= not G5987;
	G6382<= not I10278;
	G6385<= not G6119;
	G6386<= not I10282;
	G6387<= not G6121;
	G6388<= not I10286;
	G6389<= not I10289;
	G6395<= not I10293;
	G6396<= not I10296;
	G6397<= not I10299;
	G6398<= not I10302;
	G6399<= not I10305;
	G6400<= not I10308;
	G6403<= not G6128;
	G6405<= not G6133;
	G6406<= not I10314;
	G6407<= not I10317;
	G6411<= not G6135;
	G6412<= not I10322;
	G6413<= not I10325;
	G6417<= not G6136;
	G6418<= not G6137;
	G6419<= not I10331;
	G6420<= not I10334;
	G6424<= not G6140;
	G6425<= not G6141;
	G6426<= not I10340;
	G6427<= not I10343;
	G6431<= not G6145;
	G6432<= not G6146;
	G6433<= not I10349;
	G6434<= not I10352;
	G6435<= not I10355;
	G6440<= not G6150;
	G6441<= not G6151;
	G6442<= not I10362;
	G6443<= not G6157;
	G6444<= not G6158;
	G6445<= not I10367;
	G6446<= not I10370;
	G6447<= not G6166;
	G6448<= not I10374;
	G6449<= not G6172;
	G6450<= not I10378;
	G6451<= not I10381;
	G6452<= not I10384;
	G6453<= not G5817;
	G6454<= not I10388;
	G6461<= not I10391;
	G6462<= not I10394;
	G6464<= not I10398;
	G6475<= not G5987;
	G6482<= not I10412;
	G6499<= not G5867;
	G6503<= not I10421;
	G6509<= not I10427;
	G6517<= not I10434;
	G6521<= not I10437;
	G6527<= not I10445;
	G6536<= not I10456;
	G6539<= not I10461;
	G6543<= not G5888;
	G6547<= not G5893;
	G6552<= not G5733;
	G6553<= not I10477;
	G6555<= not G5740;
	G6556<= not G5747;
	G6557<= not G5748;
	G6558<= not I10484;
	G6559<= not G5758;
	G6560<= not G5759;
	G6561<= not G5773;
	G6562<= not G5774;
	G6563<= not G5783;
	G6564<= not G5784;
	G6565<= not G5790;
	G6566<= not G5791;
	G6567<= not I10495;
	G6568<= not G5797;
	G6569<= not I10499;
	G6570<= not G5949;
	G6571<= not I10503;
	G6572<= not G5805;
	G6574<= not I10514;
	G6575<= not G5949;
	G6578<= not I10526;
	G6579<= not G5949;
	G6581<= not I10531;
	G6582<= not G5949;
	G6583<= not I10535;
	G6584<= not I10538;
	G6585<= not I10541;
	G6586<= not G5949;
	G6587<= not G5827;
	G6588<= not I10546;
	G6589<= not I10549;
	G6590<= not G5949;
	G6591<= not I10553;
	G6593<= not I10557;
	G6594<= not I10560;
	G6595<= not I10563;
	G6596<= not I10566;
	G6617<= not G6019;
	G6620<= not I10573;
	G6629<= not I10584;
	G6634<= not I10589;
	G6635<= not I10592;
	G6641<= not I10598;
	G6644<= not I10601;
	G6648<= not I10607;
	G6649<= not I10610;
	G6652<= not I10613;
	G6657<= not I10620;
	G6660<= not I10623;
	G6667<= not I10630;
	G6670<= not I10633;
	G6674<= not I10639;
	G6680<= not I10643;
	G6681<= not G5830;
	G6685<= not I10648;
	G6686<= not I10651;
	G6688<= not I10655;
	G6689<= not G5830;
	G6692<= not I10659;
	G6694<= not I10663;
	G6695<= not I10666;
	G6697<= not G5949;
	G6698<= not I10671;
	G6700<= not G5949;
	G6702<= not G5949;
	G6703<= not I10678;
	G6704<= not G5949;
	G6705<= not I10682;
	G6706<= not I10685;
	G6707<= not G5949;
	G6708<= not I10689;
	G6709<= not G5949;
	G6710<= not I10693;
	G6711<= not G5949;
	G6712<= not G5984;
	G6713<= not I10698;
	G6714<= not G5867;
	G6715<= not I10702;
	G6716<= not G5949;
	G6717<= not I10706;
	G6718<= not G5949;
	G6719<= not I10710;
	G6720<= not I10713;
	G6723<= not I10716;
	G6724<= not I10719;
	G6727<= not G5997;
	G6729<= not I10724;
	G6731<= not G6001;
	G6732<= not I10729;
	G6734<= not I10733;
	G6735<= not I10736;
	G6736<= not I10739;
	G6737<= not G6016;
	G6742<= not G5830;
	G6748<= not I10753;
	G6749<= not I10756;
	G6750<= not I10759;
	G6751<= not I10762;
	G6764<= not G5987;
	G6778<= not G5987;
	G6789<= not I10789;
	G6793<= not I10795;
	G6796<= not G6252;
	G6797<= not I10801;
	G6798<= not I10804;
	G6799<= not I10807;
	G6800<= not I10810;
	G6801<= not I10813;
	G6802<= not I10816;
	G6803<= not I10819;
	G6804<= not I10822;
	G6805<= not I10825;
	G6806<= not I10828;
	G6807<= not I10831;
	G6808<= not I10834;
	G6809<= not I10837;
	G6810<= not I10840;
	G6811<= not I10843;
	G6812<= not I10846;
	G6813<= not I10849;
	G6814<= not I10852;
	G6815<= not I10855;
	G6816<= not I10858;
	G6817<= not I10861;
	G6818<= not I10864;
	G6825<= not I10873;
	G6835<= not I10885;
	G6836<= not I10888;
	G6837<= not I10891;
	G6842<= not I10898;
	G6843<= not I10901;
	G6844<= not I10904;
	G6845<= not I10907;
	G6846<= not I10910;
	G6847<= not G6482;
	G6852<= not I10914;
	G6853<= not I10917;
	G6854<= not I10920;
	G6856<= not I10924;
	G6857<= not I10927;
	G6859<= not I10937;
	G6860<= not G6475;
	G6861<= not I10941;
	G6862<= not G6720;
	G6863<= not G6740;
	G6868<= not I10946;
	G6869<= not I10949;
	G6870<= not I10952;
	G6871<= not G6724;
	G6874<= not I10958;
	G6877<= not I10963;
	G6878<= not I10966;
	G6881<= not I10971;
	G6882<= not I10974;
	G6885<= not I10979;
	G6888<= not I10984;
	G6893<= not I10991;
	G6896<= not I10996;
	G6903<= not I11005;
	G6904<= not I11008;
	G6905<= not I11011;
	G6913<= not I11021;
	G6914<= not I11024;
	G6917<= not I11029;
	G6919<= not G6453;
	G6920<= not I11034;
	G6921<= not I11037;
	G6925<= not I11043;
	G6926<= not I11046;
	G6927<= not I11049;
	G6931<= not I11055;
	G6932<= not I11058;
	G6933<= not I11061;
	G6935<= not I11065;
	G6938<= not I11068;
	G6939<= not I11071;
	G6941<= not G6503;
	G6942<= not I11076;
	G6943<= not I11079;
	G6944<= not I11082;
	G6947<= not I11085;
	G6948<= not I11088;
	G6949<= not I11091;
	G6950<= not I11094;
	G6951<= not I11097;
	G6954<= not I11100;
	G6955<= not I11103;
	G6956<= not I11106;
	G6957<= not I11109;
	G6960<= not I11112;
	G6961<= not I11115;
	G6964<= not G6509;
	G6967<= not I11119;
	G6970<= not I11122;
	G6971<= not G6517;
	G6974<= not G6365;
	G6980<= not I11127;
	G6984<= not G6382;
	G6990<= not I11132;
	G6993<= not I11135;
	G6995<= not G6482;
	G7001<= not I11140;
	G7004<= not I11143;
	G7007<= not I11146;
	G7008<= not I11149;
	G7009<= not I11152;
	G7010<= not I11155;
	G7011<= not G6503;
	G7020<= not I11159;
	G7021<= not I11162;
	G7022<= not G6389;
	G7023<= not I11166;
	G7024<= not I11169;
	G7025<= not G6400;
	G7026<= not I11173;
	G7027<= not I11176;
	G7028<= not G6407;
	G7029<= not I11180;
	G7030<= not I11183;
	G7031<= not G6413;
	G7033<= not I11188;
	G7034<= not I11191;
	G7035<= not I11194;
	G7036<= not G6420;
	G7037<= not I11198;
	G7038<= not I11201;
	G7039<= not I11204;
	G7040<= not I11207;
	G7041<= not G6427;
	G7042<= not I11211;
	G7043<= not I11214;
	G7044<= not I11217;
	G7045<= not G6435;
	G7047<= not I11222;
	G7048<= not I11225;
	G7049<= not I11228;
	G7051<= not I11232;
	G7052<= not I11235;
	G7053<= not I11238;
	G7056<= not I11249;
	G7057<= not I11252;
	G7058<= not I11255;
	G7064<= not I11269;
	G7065<= not I11272;
	G7066<= not I11275;
	G7069<= not I11286;
	G7070<= not I11289;
	G7072<= not I11293;
	G7073<= not I11296;
	G7074<= not I11299;
	G7076<= not I11303;
	G7077<= not I11306;
	G7078<= not I11309;
	G7079<= not I11312;
	G7082<= not I11315;
	G7085<= not I11318;
	G7089<= not I11322;
	G7093<= not I11326;
	G7097<= not I11330;
	G7098<= not I11333;
	G7103<= not I11338;
	G7107<= not I11342;
	G7110<= not I11345;
	G7113<= not I11348;
	G7116<= not I11351;
	G7119<= not I11354;
	G7122<= not I11357;
	G7123<= not I11360;
	G7124<= not I11363;
	G7126<= not I11367;
	G7142<= not I11383;
	G7144<= not I11387;
	G7146<= not I11391;
	G7147<= not I11394;
	G7148<= not I11397;
	G7187<= not I11405;
	G7188<= not I11408;
	G7190<= not I11412;
	G7192<= not G6742;
	G7195<= not I11417;
	G7196<= not I11420;
	G7197<= not I11423;
	G7201<= not I11427;
	G7205<= not I11433;
	G7206<= not I11436;
	G7210<= not I11440;
	G7212<= not I11444;
	G7213<= not I11447;
	G7214<= not I11450;
	G7220<= not I11456;
	G7221<= not I11459;
	G7226<= not I11464;
	G7227<= not I11467;
	G7232<= not I11472;
	G7237<= not I11477;
	G7243<= not I11483;
	G7256<= not I11489;
	G7259<= not I11494;
	G7263<= not I11498;
	G7264<= not I11501;
	G7268<= not I11505;
	G7270<= not I11515;
	G7272<= not I11519;
	G7273<= not G6365;
	G7278<= not I11524;
	G7279<= not G6382;
	G7284<= not I11528;
	G7285<= not I11531;
	G7286<= not I11534;
	G7287<= not I11537;
	G7288<= not I11540;
	G7289<= not I11543;
	G7304<= not I11560;
	G7305<= not I11563;
	G7306<= not I11566;
	G7307<= not I11569;
	G7308<= not I11572;
	G7309<= not I11575;
	G7310<= not I11578;
	G7311<= not I11581;
	G7312<= not I11584;
	G7313<= not I11587;
	G7314<= not I11590;
	G7315<= not I11593;
	G7316<= not I11596;
	G7317<= not I11599;
	G7318<= not I11602;
	G7319<= not I11605;
	G7320<= not I11608;
	G7321<= not I11611;
	G7322<= not I11614;
	G7323<= not I11617;
	G7324<= not I11620;
	G7325<= not I11623;
	G7326<= not I11626;
	G7327<= not I11629;
	G7328<= not I11632;
	G7329<= not I11635;
	G7330<= not I11638;
	G7331<= not I11641;
	G7332<= not I11644;
	G7333<= not I11647;
	G7334<= not I11650;
	G7335<= not I11653;
	G7336<= not I11656;
	G7337<= not I11659;
	G7338<= not I11662;
	G7339<= not I11665;
	G7340<= not I11668;
	G7341<= not I11671;
	G7342<= not I11674;
	G7343<= not I11677;
	G7344<= not I11680;
	G7345<= not I11683;
	G7346<= not I11686;
	G7347<= not I11689;
	G7348<= not I11692;
	G7349<= not I11695;
	G7350<= not I11698;
	G7351<= not I11701;
	G7352<= not I11704;
	G7353<= not I11707;
	G7354<= not I11710;
	G7355<= not I11713;
	G7356<= not I11716;
	G7357<= not I11719;
	G7358<= not I11722;
	G7359<= not I11725;
	G7360<= not I11728;
	G7361<= not I11731;
	G7362<= not I11734;
	G7363<= not I11737;
	G7364<= not I11740;
	G7365<= not I11743;
	G7366<= not I11746;
	G7369<= not G7273;
	G7374<= not I11752;
	G7376<= not I11756;
	G7377<= not I11759;
	G7379<= not G6863;
	G7380<= not G7279;
	G7386<= not I11767;
	G7387<= not I11770;
	G7388<= not I11773;
	G7390<= not G6847;
	G7394<= not I11778;
	G7395<= not G6941;
	G7402<= not G6860;
	G7403<= not I11783;
	G7406<= not I11786;
	G7410<= not I11790;
	G7413<= not G7197;
	G7414<= not I11794;
	G7415<= not I11797;
	G7416<= not I11800;
	G7419<= not G7206;
	G7420<= not I11804;
	G7421<= not I11807;
	G7422<= not I11810;
	G7425<= not G7214;
	G7426<= not I11814;
	G7427<= not I11817;
	G7430<= not G7221;
	G7431<= not I11821;
	G7432<= not I11824;
	G7436<= not G7227;
	G7437<= not I11829;
	G7438<= not G7232;
	G7439<= not I11833;
	G7440<= not I11836;
	G7442<= not G7237;
	G7443<= not I11841;
	G7445<= not I11845;
	G7446<= not G7148;
	G7450<= not G7148;
	G7454<= not G7148;
	G7458<= not G7123;
	G7460<= not G7148;
	G7463<= not G6921;
	G7464<= not I11858;
	G7467<= not G7148;
	G7470<= not G6927;
	G7473<= not G7148;
	G7476<= not G6933;
	G7477<= not I11869;
	G7479<= not I11873;
	G7497<= not G7148;
	G7500<= not G6943;
	G7501<= not I11879;
	G7502<= not I11882;
	G7505<= not G7148;
	G7508<= not G6950;
	G7509<= not I11889;
	G7512<= not G7148;
	G7516<= not G7148;
	G7519<= not G6956;
	G7520<= not I11898;
	G7521<= not I11901;
	G7522<= not I11904;
	G7525<= not I11921;
	G7527<= not G7148;
	G7530<= not I11926;
	G7531<= not I11929;
	G7532<= not I11932;
	G7534<= not I11942;
	G7537<= not I11947;
	G7538<= not I11950;
	G7539<= not I11953;
	G7540<= not I11956;
	G7543<= not I11961;
	G7544<= not I11964;
	G7545<= not I11967;
	G7546<= not I11970;
	G7550<= not G6974;
	G7555<= not I11989;
	G7556<= not I11992;
	G7559<= not I12009;
	G7560<= not I12012;
	G7561<= not I12015;
	G7562<= not G6984;
	G7568<= not I12026;
	G7569<= not I12029;
	G7570<= not I12032;
	G7571<= not I12035;
	G7574<= not G6995;
	G7579<= not I12053;
	G7580<= not I12056;
	G7585<= not I12081;
	G7589<= not I12099;
	G7591<= not I12103;
	G7594<= not I12120;
	G7595<= not I12123;
	G7597<= not I12133;
	G7600<= not I12150;
	G7601<= not I12153;
	G7602<= not I12156;
	G7603<= not I12159;
	G7604<= not I12162;
	G7605<= not I12165;
	G7606<= not I12168;
	G7607<= not I12171;
	G7608<= not I12174;
	G7609<= not I12177;
	G7610<= not I12180;
	G7611<= not I12183;
	G7612<= not I12186;
	G7614<= not I12190;
	G7615<= not I12193;
	G7616<= not I12196;
	G7617<= not I12199;
	G7618<= not I12202;
	G7619<= not I12205;
	G7620<= not I12208;
	G7622<= not G7067;
	G7627<= not I12223;
	G7628<= not I12226;
	G7629<= not I12229;
	G7630<= not I12232;
	G7631<= not I12235;
	G7633<= not I12239;
	G7634<= not I12242;
	G7635<= not I12245;
	G7636<= not I12248;
	G7637<= not I12251;
	G7648<= not I12255;
	G7649<= not I12258;
	G7650<= not I12261;
	G7656<= not I12265;
	G7657<= not I12268;
	G7658<= not I12271;
	G7659<= not I12274;
	G7662<= not I12279;
	G7663<= not I12282;
	G7669<= not I12286;
	G7670<= not I12289;
	G7672<= not I12293;
	G7673<= not I12296;
	G7675<= not I12300;
	G7676<= not I12303;
	G7677<= not G7148;
	G7678<= not I12307;
	G7680<= not G7148;
	G7681<= not G7148;
	G7682<= not G7148;
	G7683<= not G7148;
	G7684<= not G7148;
	G7685<= not G7148;
	G7686<= not G7148;
	G7687<= not I12318;
	G7688<= not G7148;
	G7689<= not I12322;
	G7692<= not G7148;
	G7693<= not I12326;
	G7696<= not G7148;
	G7697<= not G7101;
	G7702<= not G7079;
	G7703<= not G7085;
	G7706<= not I12335;
	G7708<= not I12339;
	G7711<= not I12344;
	G7723<= not I12354;
	G7724<= not I12357;
	G7725<= not I12360;
	G7726<= not I12363;
	G7727<= not I12366;
	G7728<= not I12369;
	G7729<= not I12372;
	G7731<= not I12376;
	G7733<= not I12380;
	G7735<= not I12384;
	G7737<= not I12388;
	G7744<= not I12397;
	G7745<= not I12400;
	G7746<= not I12403;
	G7747<= not I12406;
	G7748<= not I12409;
	G7749<= not I12412;
	G7750<= not I12415;
	G7751<= not I12418;
	G7752<= not I12421;
	G7753<= not I12424;
	G7754<= not I12427;
	G7755<= not I12430;
	G7756<= not I12433;
	G7757<= not I12436;
	G7758<= not I12439;
	G7759<= not I12442;
	G7760<= not I12445;
	G7761<= not I12448;
	G7762<= not I12451;
	G7763<= not I12454;
	G7764<= not I12457;
	G7765<= not I12460;
	G7766<= not I12463;
	G7767<= not I12466;
	G7768<= not I12469;
	G7769<= not I12472;
	G7770<= not I12475;
	G7771<= not I12478;
	G7772<= not I12481;
	G7773<= not I12484;
	G7774<= not I12487;
	G7775<= not I12490;
	G7776<= not I12493;
	G7777<= not I12496;
	G7778<= not I12499;
	G7779<= not I12502;
	G7780<= not I12505;
	G7781<= not I12508;
	G7782<= not I12511;
	G7783<= not I12514;
	G7784<= not I12517;
	G7785<= not I12520;
	G7786<= not I12523;
	G7787<= not I12526;
	G7788<= not I12529;
	G7789<= not I12532;
	G7790<= not I12535;
	G7791<= not I12538;
	G7792<= not I12541;
	G7793<= not I12544;
	G7794<= not I12547;
	G7795<= not I12550;
	G7796<= not I12553;
	G7797<= not I12556;
	G7798<= not I12559;
	G7799<= not I12562;
	G7800<= not I12565;
	G7801<= not I12568;
	G7802<= not I12571;
	G7803<= not I12574;
	G7804<= not I12577;
	G7805<= not I12580;
	G7806<= not I12583;
	G7807<= not I12586;
	G7808<= not I12589;
	G7809<= not I12592;
	G7810<= not I12595;
	G7811<= not I12598;
	G7812<= not I12601;
	G7813<= not I12604;
	G7814<= not I12607;
	G7815<= not I12610;
	G7816<= not I12613;
	G7817<= not I12616;
	G7826<= not I12627;
	G7844<= not I12631;
	G7845<= not I12634;
	G7847<= not I12638;
	G7848<= not I12641;
	G7849<= not I12644;
	G7850<= not I12647;
	G7851<= not G7479;
	G7852<= not G7479;
	G7853<= not I12652;
	G7872<= not I12655;
	G7877<= not G7479;
	G7878<= not G7479;
	G7880<= not G7479;
	G7882<= not G7479;
	G7883<= not G7689;
	G7886<= not G7479;
	G7887<= not G7693;
	G7890<= not G7479;
	G7896<= not I12678;
	G7897<= not G7712;
	G7899<= not I12683;
	G7900<= not G7712;
	G7901<= not G7712;
	G7903<= not G7446;
	G7904<= not I12690;
	G7905<= not G7450;
	G7906<= not I12694;
	G7907<= not G7664;
	G7908<= not G7454;
	G7909<= not G7664;
	G7910<= not G7460;
	G7911<= not G7664;
	G7912<= not G7651;
	G7913<= not G7467;
	G7914<= not G7651;
	G7915<= not G7473;
	G7916<= not G7651;
	G7917<= not G7497;
	G7918<= not G7505;
	G7919<= not G7512;
	G7920<= not G7516;
	G7921<= not G7463;
	G7922<= not I12712;
	G7923<= not G7527;
	G7924<= not G7470;
	G7925<= not G7476;
	G7927<= not G7500;
	G7928<= not G7508;
	G7929<= not G7519;
	G7936<= not G7712;
	G7938<= not G7403;
	G7941<= not G7406;
	G7944<= not G7410;
	G7946<= not G7416;
	G7949<= not G7422;
	G7952<= not G7427;
	G7956<= not G7432;
	G7959<= not I12751;
	G7961<= not G7664;
	G7964<= not G7651;
	G7965<= not I12759;
	G7966<= not I12762;
	G7967<= not I12765;
	G7972<= not I12770;
	G7975<= not I12773;
	G7976<= not I12776;
	G7977<= not I12779;
	G7979<= not I12783;
	G7980<= not I12786;
	G7981<= not G7624;
	G7982<= not I12790;
	G7983<= not I12793;
	G7984<= not I12796;
	G7985<= not I12799;
	G7989<= not I12805;
	G7991<= not I12809;
	G7993<= not I12813;
	G7995<= not I12817;
	G7997<= not G7697;
	G7998<= not I12822;
	G7999<= not I12825;
	G8001<= not I12829;
	G8002<= not I12832;
	G8003<= not I12835;
	G8004<= not I12838;
	G8007<= not I12843;
	G8008<= not I12846;
	G8009<= not I12849;
	G8011<= not I12853;
	G8015<= not I12857;
	G8020<= not I12862;
	G8025<= not I12867;
	G8029<= not I12871;
	G8033<= not I12875;
	G8036<= not I12878;
	G8056<= not G7671;
	G8061<= not I12901;
	G8062<= not I12904;
	G8063<= not I12907;
	G8064<= not I12910;
	G8065<= not I12913;
	G8066<= not I12916;
	G8067<= not I12919;
	G8076<= not I12930;
	G8077<= not I12933;
	G8078<= not I12936;
	G8079<= not I12939;
	G8080<= not I12942;
	G8081<= not G8000;
	G8085<= not G7932;
	G8089<= not G7934;
	G8093<= not I12948;
	G8094<= not G7987;
	G8095<= not G7942;
	G8096<= not I12953;
	G8099<= not G7990;
	G8100<= not G7947;
	G8103<= not G7994;
	G8105<= not G7992;
	G8106<= not G7950;
	G8110<= not G7996;
	G8115<= not G7953;
	G8116<= not I12971;
	G8121<= not I12978;
	G8122<= not I12981;
	G8124<= not G8011;
	G8125<= not I12986;
	G8126<= not I12989;
	G8128<= not I12993;
	G8129<= not G8015;
	G8131<= not G8020;
	G8132<= not I12999;
	G8133<= not I13002;
	G8134<= not I13005;
	G8137<= not I13010;
	G8138<= not I13013;
	G8139<= not G8025;
	G8140<= not I13017;
	G8141<= not I13020;
	G8142<= not I13023;
	G8143<= not G8029;
	G8144<= not I13027;
	G8145<= not I13030;
	G8146<= not G8033;
	G8149<= not I13036;
	G8150<= not I13039;
	G8151<= not G8036;
	G8152<= not I13043;
	G8155<= not I13048;
	G8156<= not I13051;
	G8160<= not I13057;
	G8164<= not G7872;
	G8171<= not I13068;
	G8178<= not I13083;
	G8179<= not I13086;
	G8181<= not I13096;
	G8182<= not I13099;
	G8183<= not I13102;
	G8184<= not I13105;
	G8186<= not I13109;
	G8191<= not I13114;
	G8192<= not I13117;
	G8195<= not I13122;
	G8196<= not I13125;
	G8197<= not I13128;
	G8198<= not I13131;
	G8213<= not G7826;
	G8218<= not G7826;
	G8219<= not G7826;
	G8220<= not G7826;
	G8225<= not G7826;
	G8229<= not G7826;
	G8233<= not G7872;
	G8234<= not G7826;
	G8235<= not G7967;
	G8239<= not G7826;
	G8240<= not G7972;
	G8251<= not I13166;
	G8255<= not G7986;
	G8271<= not I13185;
	G8272<= not I13188;
	G8273<= not I13191;
	G8274<= not I13194;
	G8275<= not I13197;
	G8276<= not I13200;
	G8277<= not I13203;
	G8278<= not I13206;
	G8279<= not I13209;
	G8280<= not I13212;
	G8290<= not I13224;
	G8291<= not I13227;
	G8292<= not I13230;
	G8293<= not I13233;
	G8294<= not I13236;
	G8295<= not I13239;
	G8296<= not I13242;
	G8297<= not I13245;
	G8299<= not I13255;
	G8304<= not I13280;
	G8306<= not I13290;
	G8310<= not I13314;
	G8311<= not I13317;
	G8312<= not I13320;
	G8313<= not I13323;
	G8314<= not I13326;
	G8315<= not I13329;
	G8316<= not I13332;
	G8317<= not I13335;
	G8318<= not I13338;
	G8319<= not I13341;
	G8320<= not I13344;
	G8321<= not I13347;
	G8323<= not I13351;
	G8324<= not I13354;
	G8325<= not I13357;
	G8326<= not I13360;
	G8327<= not G8164;
	G8328<= not I13364;
	G8329<= not I13367;
	G8330<= not I13370;
	G8331<= not I13373;
	G8332<= not I13376;
	G8333<= not I13379;
	G8334<= not I13382;
	G8335<= not I13385;
	G8336<= not I13388;
	G8337<= not I13391;
	G8338<= not I13394;
	G8339<= not I13397;
	G8340<= not I13400;
	G8341<= not I13403;
	G8342<= not I13406;
	G8343<= not I13409;
	G8344<= not I13412;
	G8345<= not I13415;
	G8346<= not I13418;
	G8347<= not I13421;
	G8348<= not I13424;
	G8349<= not I13427;
	G8350<= not I13430;
	G8351<= not I13433;
	G8352<= not I13436;
	G8353<= not I13439;
	G8354<= not I13442;
	G8355<= not I13445;
	G8356<= not I13448;
	G8357<= not I13451;
	G8358<= not I13454;
	G8359<= not I13457;
	G8360<= not I13460;
	G8361<= not I13463;
	G8362<= not I13466;
	G8363<= not I13469;
	G8375<= not I13475;
	G8376<= not I13478;
	G8378<= not I13482;
	G8379<= not I13485;
	G8381<= not I13489;
	G8418<= not I13568;
	G8419<= not I13571;
	G8420<= not I13574;
	G8421<= not I13577;
	G8422<= not I13580;
	G8423<= not I13583;
	G8424<= not I13586;
	G8425<= not I13589;
	G8426<= not I13592;
	G8427<= not I13595;
	G8436<= not I13606;
	G8437<= not I13609;
	G8438<= not I13612;
	G8439<= not I13615;
	G8440<= not I13618;
	G8441<= not I13621;
	G8442<= not I13624;
	G8443<= not I13627;
	G8444<= not I13630;
	G8445<= not I13633;
	G8446<= not I13636;
	G8447<= not I13639;
	G8448<= not I13642;
	G8449<= not I13645;
	G8450<= not I13648;
	G8465<= not G8289;
	G8472<= not I13666;
	G8473<= not I13669;
	G8475<= not G8314;
	G8476<= not I13674;
	G8477<= not G8317;
	G8478<= not I13678;
	G8479<= not G8319;
	G8480<= not I13682;
	G8481<= not G8324;
	G8482<= not G8329;
	G8483<= not G8332;
	G8484<= not G8336;
	G8485<= not G8341;
	G8486<= not G8348;
	G8487<= not G8350;
	G8498<= not G8353;
	G8500<= not I13695;
	G8509<= not G8366;
	G8513<= not I13708;
	G8514<= not I13711;
	G8515<= not I13714;
	G8516<= not I13717;
	G8517<= not I13720;
	G8518<= not I13723;
	G8519<= not I13726;
	G8520<= not I13729;
	G8523<= not I13732;
	G8526<= not I13735;
	G8529<= not I13738;
	G8532<= not I13741;
	G8535<= not I13744;
	G8538<= not I13747;
	G8548<= not G8390;
	G8560<= not I13773;
	G8561<= not I13776;
	G8562<= not I13779;
	G8563<= not I13782;
	G8564<= not I13785;
	G8565<= not I13788;
	G8566<= not I13791;
	G8567<= not I13794;
	G8568<= not I13797;
	G8569<= not I13800;
	G8570<= not I13803;
	G8571<= not I13806;
	G8572<= not I13809;
	G8573<= not I13812;
	G8575<= not I13816;
	G8576<= not I13819;
	G8579<= not I13822;
	G8582<= not I13825;
	G8585<= not I13828;
	G8588<= not I13831;
	G8589<= not I13834;
	G8592<= not I13837;
	G8595<= not I13840;
	G8599<= not G8546;
	G8600<= not G8475;
	G8601<= not G8477;
	G8604<= not G8479;
	G8606<= not G8481;
	G8608<= not G8482;
	G8610<= not G8483;
	G8613<= not G8484;
	G8617<= not G8465;
	G8622<= not G8485;
	G8624<= not G8486;
	G8625<= not G8487;
	G8626<= not G8498;
	G8632<= not I13915;
	G8635<= not I13918;
	G8640<= not G8512;
	G8650<= not I13933;
	G8656<= not I13941;
	G8660<= not I13945;
	G8664<= not I13949;
	G8667<= not I13952;
	G8670<= not G8551;
	G8671<= not I13956;
	G8674<= not I13959;
	G8677<= not I13962;
	G8680<= not I13965;
	G8684<= not I13969;
	G8688<= not G8507;
	G8694<= not I13975;
	G8695<= not I13978;
	G8696<= not G8656;
	G8697<= not G8660;
	G8700<= not G8574;
	G8702<= not G8664;
	G8704<= not G8667;
	G8707<= not G8671;
	G8709<= not G8674;
	G8711<= not G8677;
	G8712<= not G8680;
	G8713<= not G8684;
	G8714<= not I14005;
	G8716<= not G8576;
	G8717<= not I14010;
	G8719<= not G8579;
	G8721<= not G8582;
	G8723<= not G8585;
	G8725<= not G8589;
	G8727<= not G8592;
	G8729<= not G8595;
	G8739<= not G8640;
	G8747<= not I14040;
	G8750<= not I14045;
	G8751<= not G8632;
	G8752<= not G8635;
	G8758<= not I14055;
	G8760<= not G8670;
	G8780<= not I14077;
	G8781<= not I14080;
	G8782<= not I14083;
	G8783<= not G8746;
	G8784<= not I14087;
	G8785<= not I14090;
	G8787<= not I14094;
	G8788<= not I14097;
	G8790<= not I14101;
	G8792<= not I14105;
	G8794<= not I14109;
	G8795<= not I14112;
	G8797<= not I14116;
	G8798<= not I14119;
	G8800<= not I14123;
	G8802<= not I14127;
	G8803<= not I14130;
	G8804<= not I14133;
	G8805<= not I14136;
	G8807<= not I14140;
	G8828<= not G8744;
	G8849<= not G8745;
	G8858<= not G8743;
	G8868<= not I14176;
	G8869<= not I14179;
	G8870<= not I14182;
	G8871<= not I14185;
	G8872<= not I14188;
	G8873<= not I14191;
	G8874<= not I14194;
	G8884<= not I14224;
	G8886<= not I14228;
	G8888<= not I14232;
	G8890<= not I14236;
	G8891<= not I14239;
	G8892<= not I14242;
	G8924<= not I14249;
	G8925<= not I14252;
	G8928<= not I14257;
	G8946<= not I14295;
	G8948<= not I14299;
	G8950<= not I14303;
	G8951<= not I14306;
	G8952<= not I14309;
	G8953<= not I14312;
	G8954<= not I14315;
	G8956<= not I14319;
	G8958<= not I14323;
	G8959<= not I14326;
	G8961<= not I14330;
	G8969<= not I14340;
	G8976<= not I14349;
	G8977<= not I14352;
	G8978<= not I14355;
	G8979<= not I14358;
	G8980<= not I14361;
	G8981<= not I14364;
	G8982<= not I14367;
	G8983<= not I14370;
	G8984<= not I14373;
	G8985<= not I14376;
	G8986<= not I14379;
	G8987<= not I14382;
	G8988<= not I14385;
	G8989<= not I14388;
	G8990<= not I14391;
	G8991<= not I14394;
	G8992<= not I14397;
	G8993<= not I14400;
	G9009<= not I14405;
	G9024<= not I14409;
	G9025<= not I14412;
	G9026<= not I14415;
	G9027<= not I14418;
	G9028<= not I14421;
	G9029<= not I14424;
	G9076<= not G8892;
	G9079<= not G8892;
	G9082<= not G8892;
	G9085<= not G8892;
	G9091<= not G8892;
	G9094<= not G8892;
	G9097<= not G8892;
	G9100<= not G8892;
	G9103<= not G8892;
	G9106<= not I14439;
	G9108<= not I14449;
	G9109<= not I14452;
	G9258<= not G8892;
	G9259<= not G8892;
	G9260<= not G8892;
	G9261<= not G8892;
	G9262<= not I14473;
	G9263<= not G8892;
	G9264<= not I14477;
	G9265<= not G8892;
	G9267<= not G8892;
	G9270<= not I14485;
	G9273<= not I14490;
	G9290<= not I14494;
	G9291<= not G8892;
	G9308<= not I14499;
	G9309<= not G8892;
	G9310<= not I14503;
	G9311<= not I14506;
	G9312<= not I14509;
	G9338<= not I14519;
	G9339<= not I14522;
	G9340<= not I14525;
	G9341<= not I14528;
	G9342<= not I14531;
	G9343<= not I14534;
	G9344<= not I14537;
	G9345<= not I14540;
	G9346<= not I14543;
	G9347<= not I14546;
	G9348<= not I14549;
	G9349<= not I14552;
	G9350<= not I14555;
	G9351<= not I14558;
	G9352<= not I14561;
	G9353<= not I14564;
	G9354<= not I14567;
	G9355<= not I14570;
	G9356<= not I14573;
	G9360<= not I14579;
	G9424<= not G9076;
	G9427<= not G9079;
	G9429<= not G9082;
	G9431<= not G9085;
	G9432<= not G9313;
	G9448<= not G9091;
	G9449<= not G9094;
	G9450<= not G9097;
	G9451<= not I14642;
	G9452<= not I14645;
	G9453<= not G9100;
	G9473<= not G9103;
	G9474<= not G9331;
	G9490<= not G9324;
	G9505<= not G9052;
	G9507<= not G9268;
	G9508<= not G9271;
	G9525<= not G9257;
	G9526<= not G9256;
	G9527<= not I14668;
	G9529<= not I14672;
	G9530<= not I14675;
	G9531<= not I14678;
	G9532<= not I14681;
	G9533<= not I14684;
	G9534<= not I14687;
	G9535<= not I14690;
	G9553<= not I14694;
	G9554<= not I14697;
	G9556<= not I14701;
	G9572<= not I14709;
	G9576<= not I14713;
	G9661<= not I14786;
	G9666<= not I14793;
	G9668<= not G9490;
	G9670<= not I14799;
	G9671<= not I14802;
	G9672<= not I14805;
	G9679<= not G9452;
	G9732<= not I14873;
	G9733<= not I14876;
	G9739<= not I14884;
	G9741<= not I14888;
	G9745<= not G9454;
	G9760<= not G9454;
	G9761<= not G9454;
	G9762<= not I14903;
	G9763<= not I14906;
	G9764<= not G9432;
	G9765<= not I14910;
	G9766<= not G9432;
	G9767<= not I14914;
	G9768<= not G9432;
	G9769<= not I14918;
	G9770<= not G9432;
	G9771<= not G9432;
	G9772<= not G9432;
	G9773<= not G9474;
	G9774<= not G9474;
	G9775<= not G9474;
	G9777<= not G9474;
	G9778<= not G9474;
	G9780<= not G9474;
	G9782<= not I14933;
	G9802<= not G9490;
	G9804<= not I14939;
	G9807<= not G9490;
	G9809<= not I14944;
	G9812<= not G9490;
	G9813<= not I14948;
	G9814<= not G9490;
	G9816<= not G9490;
	G9818<= not I14955;
	G9819<= not I14958;
	G9820<= not I14961;
	G9821<= not I14964;
	G9822<= not I14967;
	G9823<= not I14970;
	G9824<= not I14973;
	G9825<= not I14976;
	G9826<= not I14979;
	G9827<= not I14982;
	G9832<= not I14989;
	G9845<= not G9679;
	G9875<= not I15036;
	G9883<= not I15060;
	G9884<= not I15063;
	G9887<= not I15068;
	G9889<= not I15072;
	G9890<= not I15075;
	G9892<= not I15079;
	G9893<= not I15082;
	G9894<= not I15085;
	G9895<= not I15088;
	G9919<= not I15114;
	G9930<= not I15127;
	G9958<= not I15157;
	G9961<= not I15162;
	G9980<= not I15181;
	G9984<= not I15184;
	G9987<= not I15187;
	G9990<= not I15190;
	G9993<= not I15193;
	G9994<= not I15196;
	G10031<= not I15229;
	G10032<= not I15232;
	G10033<= not I15235;
	G10034<= not I15238;
	G10035<= not I15241;
	G10039<= not I15244;
	G10040<= not I15247;
	G10041<= not I15250;
	G10042<= not I15253;
	G10044<= not I15263;
	G10047<= not I15266;
	G10050<= not I15269;
	G10051<= not I15272;
	G10056<= not I15275;
	G10057<= not I15278;
	G10058<= not I15281;
	G10062<= not I15284;
	G10063<= not I15287;
	G10064<= not I15290;
	G10065<= not I15293;
	G10069<= not I15296;
	G10074<= not I15299;
	G10075<= not I15302;
	G10079<= not I15305;
	G10080<= not I15308;
	G10083<= not I15311;
	G10087<= not I15314;
	G10088<= not I15317;
	G10091<= not I15320;
	G10092<= not I15323;
	G10093<= not I15326;
	G10094<= not I15329;
	G10098<= not I15332;
	G10101<= not I15335;
	G10104<= not I15338;
	G10107<= not I15341;
	G10110<= not I15344;
	G10111<= not I15347;
	G10114<= not I15350;
	G10115<= not I15353;
	G10116<= not I15356;
	G10117<= not I15359;
	G10118<= not I15362;
	G10119<= not I15365;
	G10120<= not I15368;
	G10121<= not I15371;
	G10122<= not I15374;
	G10125<= not I15377;
	G10126<= not I15380;
	G10127<= not I15383;
	G10128<= not I15386;
	G10129<= not I15389;
	G10130<= not I15392;
	G10131<= not I15395;
	G10132<= not G10063;
	G10133<= not G10064;
	G10134<= not I15400;
	G10135<= not I15403;
	G10136<= not I15406;
	G10137<= not I15409;
	G10138<= not I15412;
	G10139<= not I15415;
	G10140<= not I15418;
	G10141<= not I15421;
	G10142<= not I15424;
	G10143<= not I15427;
	G10145<= not I15437;
	G10148<= not G10121;
	G10150<= not I15448;
	G10154<= not I15458;
	G10155<= not I15461;
	G10156<= not I15464;
	G10157<= not I15467;
	G10158<= not I15470;
	G10159<= not I15473;
	G10160<= not I15476;
	G10161<= not I15479;
	G10162<= not I15482;
	G10163<= not I15485;
	G10164<= not I15488;
	G10165<= not I15491;
	G10166<= not I15494;
	G10167<= not I15497;
	G10168<= not I15500;
	G10169<= not I15503;
	G10170<= not G10118;
	G10171<= not I15507;
	G10172<= not I15510;
	G10173<= not G10120;
	G10174<= not I15514;
	G10175<= not I15517;
	G10176<= not I15520;
	G10177<= not I15523;
	G10178<= not I15526;
	G10179<= not G10041;
	G10182<= not I15530;
	G10183<= not G10042;
	G10184<= not G10039;
	G10185<= not G10040;
	G10186<= not I15536;
	G10187<= not I15539;
	G10188<= not I15542;
	G10189<= not I15545;
	G10190<= not I15548;
	G10191<= not I15551;
	G10192<= not I15554;
	G10193<= not G10057;
	G10194<= not G10062;
	G10195<= not I15559;
	G10196<= not I15562;
	G10197<= not I15565;
	G10198<= not I15568;
	G10199<= not G10172;
	G10200<= not G10169;
	G10201<= not G10175;
	G10202<= not G10171;
	G10203<= not G10177;
	G10204<= not G10174;
	G10205<= not G10176;
	G10206<= not G10178;
	G10207<= not G10186;
	G10208<= not I15580;
	G10211<= not I15583;
	G10214<= not I15586;
	G10217<= not I15589;
	G10220<= not I15592;
	G10223<= not I15595;
	G10226<= not I15598;
	G10227<= not I15601;
	G10228<= not I15604;
	G10233<= not G10187;
	G10234<= not G10188;
	G10235<= not G10189;
	G10236<= not G10190;
	G10238<= not G10191;
	G10241<= not G10192;
	G10242<= not I15632;
	G10243<= not I15635;
	G10244<= not G10131;
	G10247<= not I15639;
	G10248<= not G10134;
	G10249<= not G10135;
	G10250<= not G10136;
	G10251<= not G10195;
	G10252<= not G10137;
	G10253<= not G10138;
	G10254<= not G10196;
	G10255<= not G10139;
	G10256<= not G10140;
	G10257<= not G10197;
	G10258<= not G10198;
	G10259<= not G10141;
	G10260<= not G10125;
	G10261<= not G10126;
	G10262<= not G10142;
	G10263<= not G10127;
	G10264<= not G10128;
	G10265<= not G10143;
	G10266<= not G10129;
	G10267<= not G10130;
	G10269<= not G10154;
	G10270<= not G10156;
	G10271<= not I15665;
	G10272<= not G10168;
	G10275<= not I15669;
	G10276<= not I15672;
	G10277<= not I15675;
	G10278<= not G10182;
	G10279<= not G10158;
	G10280<= not G10160;
	G10281<= not G10162;
	G10282<= not G10164;
	G10283<= not G10166;
	G10284<= not G10167;
	G10288<= not I15688;
	G10289<= not I15691;
	G10290<= not I15694;
	G10292<= not I15698;
	G10293<= not I15701;
	G10294<= not I15704;
	G10296<= not I15708;
	G10305<= not I15725;
	G10307<= not I15729;
	G10309<= not I15733;
	G10310<= not I15736;
	G10311<= not G10242;
	G10313<= not I15741;
	G10314<= not I15744;
	G10315<= not G10243;
	G10317<= not I15749;
	G10318<= not I15752;
	G10319<= not G10270;
	G10320<= not I15756;
	G10321<= not I15759;
	G10323<= not I15763;
	G10326<= not I15768;
	G10327<= not I15771;
	G10329<= not I15775;
	G10330<= not I15778;
	G10332<= not I15782;
	G10335<= not I15787;
	G10342<= not I15792;
	G10343<= not I15795;
	G10344<= not I15798;
	G10345<= not I15801;
	G10346<= not I15804;
	G10347<= not I15807;
	G10349<= not I15811;
	G10350<= not I15814;
	G10351<= not I15817;
	G10352<= not I15820;
	G10353<= not I15823;
	G10354<= not I15826;
	G10355<= not I15829;
	G10356<= not I15832;
	G10361<= not G10268;
	G10377<= not I15855;
	G10378<= not I15858;
	G10379<= not I15861;
	G10380<= not I15864;
	G10387<= not G10357;
	G10388<= not G10305;
	G10389<= not G10307;
	G10390<= not G10309;
	G10391<= not G10313;
	G10393<= not G10317;
	G10395<= not G10320;
	G10400<= not G10348;
	G10421<= not G10331;
	G10431<= not G10328;
	G10437<= not G10333;
	G10439<= not G10334;
	G10444<= not G10325;
	G10455<= not I15956;
	G10456<= not I15959;
	G10457<= not I15962;
	G10458<= not I15965;
	G10459<= not I15968;
	G10460<= not I15971;
	G10461<= not I15974;
	G10462<= not I15977;
	G10463<= not I15980;
	G10464<= not I15983;
	G10465<= not I15986;
	G10466<= not I15989;
	G10471<= not G10378;
	G10473<= not G10380;
	G10486<= not I16095;
	G10487<= not I16098;
	G10488<= not I16101;
	G10490<= not I16105;
	G10491<= not I16108;
	G10492<= not I16111;
	G10493<= not I16114;
	G10498<= not I16121;
	G10499<= not I16124;
	G10523<= not G10456;
	G10524<= not G10458;
	G10525<= not G10499;
	G10526<= not G10460;
	G10527<= not G10462;
	G10528<= not G10464;
	G10530<= not G10466;
	G10531<= not G10471;
	G10532<= not G10473;
	G10534<= not I16169;
	G10535<= not I16172;
	G10536<= not I16175;
	G10537<= not I16178;
	G10538<= not I16181;
	G10539<= not I16184;
	G10540<= not I16187;
	G10541<= not I16190;
	G10542<= not I16193;
	G10543<= not I16196;
	G10545<= not I16200;
	G10546<= not I16203;
	G10547<= not I16206;
	G10548<= not I16209;
	G10551<= not I16214;
	G10552<= not I16217;
	G10553<= not I16220;
	G10571<= not I16236;
	G10574<= not I16239;
	G10575<= not G10523;
	G10576<= not G10524;
	G10577<= not G10526;
	G10578<= not G10527;
	G10579<= not G10528;
	G10580<= not G10530;
	G10584<= not G10522;
	G10589<= not I16252;
	G10590<= not I16255;
	G10591<= not I16258;
	G10592<= not I16261;
	G10593<= not I16264;
	G10596<= not I16269;
	G10598<= not I16273;
	G10600<= not I16277;
	G10604<= not I16280;
	G10608<= not I16283;
	G10612<= not I16286;
	G10616<= not I16289;
	G10619<= not I16292;
	G10620<= not I16295;
	G10621<= not I16298;
	G10628<= not I16307;
	G10629<= not G10583;
	G10630<= not I16311;
	G10668<= not G10563;
	G10674<= not G10584;
	G10675<= not G10574;
	G10676<= not G10570;
	G10679<= not G10584;
	G10683<= not G10612;
	G10687<= not I16356;
	G10691<= not I16360;
	G10692<= not I16363;
	G10695<= not I16366;
	G10696<= not G10621;
	G10697<= not I16370;
	G10698<= not I16373;
	G10699<= not I16376;
	G10700<= not I16379;
	G10708<= not I16387;
	G10729<= not G10630;
	G10730<= not I16407;
	G10734<= not I16413;
	G10735<= not I16416;
	G10747<= not I16432;
	G10754<= not I16439;
	G10774<= not I16458;
	G10775<= not I16461;
	G10781<= not I16475;
	G10783<= not I16479;
	G10786<= not I16484;
	G10787<= not I16487;
	G10792<= not I16492;
	G10794<= not I16496;
	G10796<= not I16500;
	G10801<= not I16507;
	G10802<= not I16510;
	G10803<= not G10708;
	G10804<= not I16514;
	G10806<= not I16518;
	G10819<= not I16525;
	G10820<= not I16528;
	G10821<= not I16531;
	G10822<= not I16534;
	G10825<= not I16537;
	G10826<= not I16540;
	G10827<= not I16543;
	G10848<= not I16546;
	G10850<= not I16550;
	G10851<= not I16553;
	G10852<= not G10740;
	G10854<= not G10708;
	G10867<= not I16571;
	G10868<= not I16574;
	G10869<= not I16577;
	G10870<= not I16580;
	G10871<= not I16583;
	G10872<= not I16586;
	G10873<= not I16589;
	G10874<= not I16592;
	G10875<= not I16595;
	G10876<= not I16598;
	G10877<= not I16601;
	G10878<= not I16604;
	G10879<= not I16607;
	G10880<= not I16610;
	G10881<= not I16613;
	G10882<= not I16616;
	G10883<= not G10809;
	G10884<= not G10809;
	G10885<= not G10809;
	G10887<= not I16623;
	G10888<= not I16626;
	G10889<= not I16629;
	G10890<= not I16632;
	G10891<= not I16635;
	G10892<= not I16638;
	G10893<= not I16641;
	G10894<= not I16644;
	G10895<= not I16647;
	G10896<= not I16650;
	G10897<= not G10827;
	G10899<= not G10803;
	G10900<= not I16656;
	G10901<= not G10802;
	G10902<= not I16660;
	G10903<= not G10809;
	G10904<= not I16664;
	G10905<= not I16667;
	G10906<= not I16670;
	G10907<= not I16673;
	G10908<= not I16676;
	G10909<= not I16679;
	G10910<= not I16682;
	G10911<= not I16685;
	G10912<= not I16688;
	G10913<= not I16691;
	G10926<= not G10827;
	G10927<= not G10827;
	G10928<= not G10827;
	G10929<= not G10827;
	G10930<= not G10827;
	G10931<= not G10827;
	G10932<= not G10827;
	G10934<= not G10827;
	G10935<= not G10827;
	G10947<= not I16708;
	G10972<= not I16717;
	G10973<= not I16720;
	G10974<= not I16723;
	G11014<= not I16735;
	G11016<= not I16739;
	G11017<= not I16742;
	G11033<= not I16760;
	G11034<= not I16763;
	G11035<= not I16766;
	G11036<= not I16769;
	G11037<= not I16772;
	G11038<= not I16775;
	G11039<= not I16778;
	G11040<= not I16781;
	G11041<= not I16784;
	G11042<= not I16787;
	G11043<= not I16790;
	G11044<= not I16793;
	G11045<= not I16796;
	G11046<= not I16799;
	G11047<= not I16802;
	G11048<= not I16805;
	G11049<= not I16808;
	G11050<= not I16811;
	G11051<= not I16814;
	G11052<= not I16817;
	G11053<= not G10950;
	G11054<= not G10950;
	G11055<= not G10950;
	G11056<= not G10950;
	G11057<= not G10937;
	G11059<= not G10974;
	G11060<= not G10937;
	G11061<= not G10974;
	G11062<= not G10937;
	G11063<= not G10974;
	G11064<= not G10974;
	G11065<= not G10974;
	G11066<= not G10974;
	G11067<= not G10974;
	G11068<= not G10974;
	G11069<= not G10974;
	G11071<= not G10913;
	G11072<= not G10913;
	G11073<= not G10913;
	G11074<= not G10901;
	G11075<= not G10937;
	G11076<= not I16843;
	G11078<= not I16847;
	G11079<= not I16850;
	G11080<= not I16853;
	G11081<= not I16856;
	G11082<= not I16859;
	G11083<= not G10913;
	G11084<= not I16863;
	G11086<= not I16867;
	G11088<= not I16871;
	G11096<= not I16879;
	G11106<= not G10974;
	G11107<= not G10974;
	G11108<= not G10974;
	G11109<= not G10974;
	G11110<= not G10974;
	G11111<= not G10974;
	G11112<= not I16897;
	G11155<= not G10950;
	G11157<= not G10950;
	G11159<= not G10950;
	G11160<= not G10950;
	G11162<= not G10950;
	G11163<= not I16920;
	G11179<= not I16938;
	G11180<= not I16941;
	G11181<= not I16944;
	G11182<= not I16947;
	G11183<= not I16950;
	G11184<= not I16953;
	G11185<= not I16956;
	G11191<= not G11112;
	G11193<= not G11112;
	G11195<= not G11112;
	G11197<= not G11112;
	G11199<= not G11112;
	G11200<= not G11112;
	G11202<= not G11112;
	G11203<= not G11112;
	G11205<= not G11112;
	G11206<= not I16979;
	G11207<= not I16982;
	G11208<= not G11077;
	G11239<= not G11112;
	G11241<= not G11112;
	G11242<= not G11112;
	G11243<= not G11112;
	G11244<= not G11112;
	G11245<= not G11112;
	G11284<= not G11208;
	G11287<= not G11207;
	G11289<= not I17070;
	G11301<= not I17084;
	G11307<= not I17092;
	G11309<= not I17096;
	G11311<= not I17100;
	G11313<= not I17104;
	G11315<= not I17108;
	G11317<= not I17112;
	G11319<= not I17116;
	G11322<= not I17121;
	G11323<= not I17124;
	G11339<= not I17142;
	G11341<= not I17146;
	G11342<= not I17149;
	G11343<= not I17152;
	G11344<= not I17155;
	G11345<= not I17158;
	G11346<= not I17161;
	G11347<= not I17164;
	G11348<= not G11276;
	G11350<= not G11287;
	G11351<= not I17170;
	G11352<= not I17173;
	G11353<= not I17176;
	G11354<= not I17179;
	G11357<= not I17182;
	G11360<= not I17185;
	G11363<= not I17188;
	G11366<= not I17191;
	G11369<= not I17194;
	G11373<= not I17198;
	G11377<= not I17202;
	G11381<= not I17206;
	G11384<= not I17209;
	G11388<= not I17213;
	G11389<= not I17216;
	G11390<= not I17219;
	G11394<= not I17225;
	G11395<= not I17228;
	G11396<= not I17231;
	G11397<= not I17234;
	G11398<= not I17237;
	G11399<= not I17240;
	G11400<= not I17243;
	G11401<= not I17246;
	G11402<= not I17249;
	G11403<= not I17252;
	G11404<= not I17255;
	G11405<= not I17258;
	G11406<= not I17261;
	G11408<= not I17265;
	G11409<= not I17268;
	G11410<= not I17271;
	G11411<= not I17274;
	G11412<= not I17277;
	G11417<= not I17302;
	G11419<= not I17312;
	G11420<= not I17315;
	G11421<= not I17318;
	G11422<= not I17321;
	G11423<= not I17324;
	G11424<= not I17327;
	G11426<= not I17331;
	G11427<= not I17334;
	G11428<= not I17337;
	G11429<= not I17340;
	G11431<= not I17344;
	G11432<= not I17347;
	G11433<= not I17350;
	G11434<= not I17353;
	G11435<= not I17356;
	G11436<= not I17359;
	G11437<= not I17362;
	G11438<= not I17365;
	G11439<= not I17368;
	G11440<= not I17371;
	G11441<= not I17374;
	G11442<= not I17377;
	G11444<= not I17381;
	G11445<= not I17384;
	G11446<= not I17387;
	G11447<= not I17390;
	G11450<= not I17407;
	G11451<= not I17410;
	G11452<= not I17413;
	G11453<= not I17416;
	G11454<= not I17419;
	G11457<= not I17424;
	G11466<= not I17435;
	G11467<= not I17438;
	G11468<= not I17441;
	G11469<= not I17444;
	G11470<= not I17447;
	G11471<= not I17450;
	G11472<= not I17453;
	G11473<= not I17456;
	G11475<= not I17466;
	G11479<= not I17470;
	G11489<= not I17482;
	G11495<= not I17500;
	G11497<= not I17510;
	G11498<= not I17513;
	G11499<= not I17516;
	G11500<= not I17519;
	G11501<= not I17522;
	G11502<= not I17525;
	G11503<= not I17528;
	G11504<= not I17531;
	G11505<= not I17534;
	G11506<= not I17537;
	G11507<= not I17540;
	G11508<= not I17543;
	G11509<= not I17546;
	G11510<= not I17549;
	G11511<= not I17552;
	G11512<= not I17555;
	G11513<= not I17558;
	G11515<= not G11490;
	G11518<= not I17563;
	G11539<= not G11519;
	G11540<= not G11519;
	G11541<= not G11519;
	G11542<= not G11519;
	G11543<= not G11519;
	G11545<= not G11519;
	G11546<= not G11519;
	G11547<= not G11519;
	G11548<= not G11519;
	G11550<= not I17591;
	G11572<= not G11561;
	G11573<= not G11561;
	G11574<= not G11561;
	G11575<= not G11561;
	G11576<= not I17610;
	G11577<= not I17613;
	G11578<= not I17616;
	G11593<= not I17633;
	G11594<= not I17636;
	G11596<= not G11580;
	G11598<= not I17642;
	G11611<= not I17657;
	G11614<= not I17662;
	G11616<= not I17666;
	G11617<= not I17669;
	G11618<= not I17672;
	G11619<= not I17675;
	G11620<= not I17678;
	G11621<= not I17681;
	G11622<= not I17684;
	G11623<= not I17687;
	G11626<= not I17692;
	G11627<= not I17695;
	G11628<= not I17698;
	G11629<= not I17701;
	G11630<= not I17704;
	G11631<= not I17707;
	G11632<= not I17710;
	G11633<= not I17713;
	G11634<= not I17716;
	G11635<= not I17719;
	G11638<= not I17724;
	G11642<= not I17730;
	G11643<= not I17733;
	G11644<= not I17736;
	G11645<= not I17739;
	G11646<= not I17742;
	G11648<= not I17746;
	G11649<= not I17749;
	G11650<= not I17752;
	G11651<= not I17755;
	G11652<= not I17758;
	G11653<= not I17761;
	G11654<= not I17764;
	G11655<= not I17767;
	G11656<= not I17770;
	G11657<= not I17773;
	I4777<= not G18;
	I4780<= not G872;
	I4783<= not G873;
	I4786<= not G109;
	I4820<= not G865;
	I4850<= not G1958;
	I4859<= not G578;
	I4866<= not G579;
	I4869<= not G253;
	I4873<= not G105;
	I4876<= not G580;
	I4879<= not G256;
	I4883<= not G581;
	I4886<= not G257;
	I4891<= not G582;
	I4894<= not G258;
	I4900<= not G583;
	I4903<= not G259;
	I4906<= not G119;
	I4917<= not G584;
	I4920<= not G260;
	I4924<= not G123;
	I4935<= not G585;
	I4938<= not G261;
	I4948<= not G586;
	I4951<= not G262;
	I4961<= not G254;
	I4992<= not G1170;
	I5002<= not G1173;
	I5020<= not G1176;
	I5031<= not G928;
	I5041<= not G1179;
	I5044<= not G1182;
	I5047<= not G1185;
	I5050<= not G1216;
	I5053<= not G1188;
	I5057<= not G1961;
	I5060<= not G1191;
	I5064<= not G1690;
	I5067<= not G33;
	I5070<= not G1194;
	I5073<= not G34;
	I5077<= not G35;
	I5080<= not G36;
	I5089<= not G1854;
	I5092<= not G32;
	I5095<= not G37;
	I5098<= not G38;
	I5101<= not G1960;
	I5111<= not G39;
	I5116<= not G40;
	I5120<= not G622;
	I5142<= not G639;
	I5149<= not G1453;
	I5171<= not G1419;
	I5174<= not G52;
	I5192<= not G55;
	I5198<= not G143;
	I5210<= not G58;
	I5218<= not G1104;
	I5221<= not G1407;
	I5224<= not G61;
	I5237<= not G1107;
	I5240<= not G64;
	I5245<= not G925;
	I5248<= not G1110;
	I5251<= not G1424;
	I5254<= not G1700;
	I5258<= not G67;
	I5271<= not G70;
	I5276<= not G1411;
	I5279<= not G73;
	I5289<= not G49;
	I5292<= not G76;
	I5304<= not G79;
	I5308<= not G97;
	I5311<= not G98;
	I5332<= not G756;
	I5336<= not G1700;
	I5348<= not G746;
	I5378<= not G1857;
	I5383<= not G886;
	I5388<= not G889;
	I5391<= not G1101;
	I5395<= not G892;
	I5399<= not G895;
	I5403<= not G636;
	I5406<= not G898;
	I5410<= not G901;
	I5414<= not G904;
	I5418<= not G907;
	I5421<= not G549;
	I5424<= not G910;
	I5427<= not G913;
	I5430<= not G916;
	I5435<= not G18;
	I5438<= not G18;
	I5441<= not G919;
	I5445<= not G922;
	I5475<= not G1289;
	I5478<= not G1212;
	I5494<= not G1690;
	I5497<= not G587;
	I5510<= not G588;
	I5513<= not G255;
	I5525<= not G589;
	I5549<= not G868;
	I5555<= not G110;
	I5561<= not G869;
	I5565<= not G1713;
	I5579<= not G1197;
	I5584<= not G1200;
	I5588<= not G1203;
	I5632<= not G932;
	I5638<= not G936;
	I5641<= not G546;
	I5646<= not G940;
	I5652<= not G554;
	I5655<= not G557;
	I5658<= not G560;
	I5662<= not G563;
	I5667<= not G566;
	I5672<= not G569;
	I5684<= not G572;
	I5695<= not G575;
	I5704<= not G2056;
	I5707<= not G2418;
	I5710<= not G2431;
	I5713<= not G2436;
	I5716<= not G2068;
	I5719<= not G2072;
	I5722<= not G2075;
	I5725<= not G2079;
	I5728<= not G2084;
	I5731<= not G2089;
	I5734<= not G2097;
	I5737<= not G2100;
	I5740<= not G2341;
	I5751<= not G2296;
	I5754<= not G2304;
	I5765<= not G2004;
	I5789<= not G2162;
	I5792<= not G2080;
	I5795<= not G2462;
	I5798<= not G2085;
	I5801<= not G1984;
	I5809<= not G2356;
	I5812<= not G2090;
	I5815<= not G1994;
	I5818<= not G2098;
	I5821<= not G2101;
	I5824<= not G2502;
	I5827<= not G2271;
	I5830<= not G2067;
	I5833<= not G2103;
	I5837<= not G2507;
	I5840<= not G2432;
	I5843<= not G2509;
	I5847<= not G2275;
	I5850<= not G2273;
	I5854<= not G2523;
	I5858<= not G2529;
	I5862<= not G2537;
	I5909<= not G2207;
	I5913<= not G2169;
	I5916<= not G2217;
	I5919<= not G2530;
	I5922<= not G2170;
	I5926<= not G2172;
	I5929<= not G2225;
	I5932<= not G2539;
	I5935<= not G2174;
	I5940<= not G2175;
	I5943<= not G2233;
	I5946<= not G2176;
	I5949<= not G2540;
	I5952<= not G2506;
	I5957<= not G2178;
	I5960<= not G2239;
	I5963<= not G2179;
	I5966<= not G2541;
	I5970<= not G2185;
	I5973<= not G2247;
	I5976<= not G2186;
	I5979<= not G2543;
	I5982<= not G2510;
	I5986<= not G2194;
	I5989<= not G2252;
	I5992<= not G2195;
	I5995<= not G2196;
	I5998<= not G2197;
	I6001<= not G2548;
	I6007<= not G2199;
	I6010<= not G2256;
	I6013<= not G2200;
	I6016<= not G2201;
	I6019<= not G2554;
	I6022<= not G2258;
	I6025<= not G2259;
	I6028<= not G2208;
	I6031<= not G2209;
	I6034<= not G2210;
	I6037<= not G2560;
	I6040<= not G2216;
	I6043<= not G2267;
	I6046<= not G2218;
	I6049<= not G2219;
	I6052<= not G2220;
	I6055<= not G2569;
	I6061<= not G2246;
	I6065<= not G2226;
	I6068<= not G2227;
	I6071<= not G2269;
	I6074<= not G2228;
	I6077<= not G2349;
	I6080<= not G2108;
	I6085<= not G2234;
	I6088<= not G2235;
	I6091<= not G2270;
	I6094<= not G2110;
	I6097<= not G2391;
	I6102<= not G2240;
	I6106<= not G2116;
	I6118<= not G2248;
	I6121<= not G2121;
	I6133<= not G2253;
	I6150<= not G2122;
	I6156<= not G2119;
	I6159<= not G2123;
	I6163<= not G2547;
	I6173<= not G2125;
	I6183<= not G2131;
	I6193<= not G2155;
	I6196<= not G2462;
	I6217<= not G2302;
	I6220<= not G883;
	I6233<= not G2299;
	I6240<= not G878;
	I6247<= not G2462;
	I6256<= not G2462;
	I6260<= not G2025;
	I6264<= not G2118;
	I6273<= not G2482;
	I6277<= not G1206;
	I6282<= not G2231;
	I6294<= not G2238;
	I6299<= not G2242;
	I6302<= not G2243;
	I6343<= not G1963;
	I6347<= not G2462;
	I6356<= not G2459;
	I6360<= not G2261;
	I6363<= not G2459;
	I6367<= not G2045;
	I6370<= not G2356;
	I6373<= not G2024;
	I6381<= not G2257;
	I6385<= not G2260;
	I6388<= not G2329;
	I6391<= not G2478;
	I6395<= not G2334;
	I6398<= not G2335;
	I6403<= not G2337;
	I6406<= not G2339;
	I6409<= not G2356;
	I6414<= not G2342;
	I6417<= not G2344;
	I6421<= not G2346;
	I6424<= not G2462;
	I6428<= not G2348;
	I6432<= not G2350;
	I6436<= not G2351;
	I6439<= not G2352;
	I6443<= not G2363;
	I6454<= not G2368;
	I6461<= not G2261;
	I6474<= not G2297;
	I6477<= not G2069;
	I6480<= not G2462;
	I6484<= not G2073;
	I6495<= not G2076;
	I6498<= not G2958;
	I6501<= not G2578;
	I6504<= not G3214;
	I6507<= not G2808;
	I6510<= not G3267;
	I6513<= not G2812;
	I6517<= not G3271;
	I6520<= not G3186;
	I6523<= not G2819;
	I6528<= not G3274;
	I6531<= not G3186;
	I6535<= not G2826;
	I6538<= not G2827;
	I6543<= not G3186;
	I6546<= not G2987;
	I6549<= not G2838;
	I6553<= not G3186;
	I6557<= not G3086;
	I6560<= not G2845;
	I6565<= not G2614;
	I6569<= not G3186;
	I6572<= not G2853;
	I6576<= not G2617;
	I6580<= not G3186;
	I6587<= not G2620;
	I6590<= not G3186;
	I6598<= not G2623;
	I6601<= not G3186;
	I6611<= not G2626;
	I6616<= not G3186;
	I6624<= not G2629;
	I6639<= not G2632;
	I6643<= not G3008;
	I6648<= not G2635;
	I6654<= not G2952;
	I6661<= not G2752;
	I6671<= not G2757;
	I6676<= not G2759;
	I6679<= not G2902;
	I6686<= not G3015;
	I6690<= not G2743;
	I6694<= not G2749;
	I6702<= not G2801;
	I6726<= not G3306;
	I6733<= not G3321;
	I6738<= not G3113;
	I6742<= not G3326;
	I6754<= not G2906;
	I6757<= not G2732;
	I6767<= not G2914;
	I6784<= not G2742;
	I6789<= not G2748;
	I6799<= not G2750;
	I6802<= not G2751;
	I6812<= not G3290;
	I6815<= not G2755;
	I6818<= not G2758;
	I6821<= not G3015;
	I6832<= not G2909;
	I6844<= not G2915;
	I6851<= not G2937;
	I6856<= not G3318;
	I6861<= not G2942;
	I6867<= not G2949;
	I6870<= not G2852;
	I6876<= not G2956;
	I6888<= not G2960;
	I6891<= not G2962;
	I6894<= not G2813;
	I6898<= not G2964;
	I6901<= not G2818;
	I6904<= not G2820;
	I6907<= not G2994;
	I6911<= not G2825;
	I6914<= not G2828;
	I6917<= not G2832;
	I6921<= not G2839;
	I6924<= not G2843;
	I6929<= not G2846;
	I6932<= not G2850;
	I6938<= not G2854;
	I6941<= not G2858;
	I6944<= not G2859;
	I6947<= not G2860;
	I6952<= not G2867;
	I6955<= not G2871;
	I6958<= not G2872;
	I6962<= not G2791;
	I6965<= not G2880;
	I6968<= not G2881;
	I6971<= not G2882;
	I6976<= not G2884;
	I6979<= not G2888;
	I6982<= not G2889;
	I6985<= not G2890;
	I6996<= not G2904;
	I6999<= not G2905;
	I7002<= not G2907;
	I7006<= not G2912;
	I7009<= not G2913;
	I7014<= not G2919;
	I7017<= not G3068;
	I7022<= not G2941;
	I7029<= not G2946;
	I7043<= not G2908;
	I7048<= not G2807;
	I7054<= not G3093;
	I7061<= not G3050;
	I7064<= not G2984;
	I7070<= not G3138;
	I7076<= not G2985;
	I7086<= not G3142;
	I7096<= not G3186;
	I7099<= not G3228;
	I7104<= not G3186;
	I7109<= not G2970;
	I7112<= not G3186;
	I7118<= not G2979;
	I7131<= not G2640;
	I7140<= not G2641;
	I7143<= not G2614;
	I7151<= not G2642;
	I7154<= not G2617;
	I7157<= not G3015;
	I7163<= not G2643;
	I7166<= not G2620;
	I7173<= not G2644;
	I7176<= not G2623;
	I7182<= not G2645;
	I7185<= not G2626;
	I7191<= not G2646;
	I7194<= not G2629;
	I7202<= not G2647;
	I7205<= not G2632;
	I7210<= not G2798;
	I7213<= not G2635;
	I7216<= not G2952;
	I7220<= not G3213;
	I7233<= not G2817;
	I7236<= not G3219;
	I7240<= not G2824;
	I7244<= not G3226;
	I7249<= not G2833;
	I7255<= not G3227;
	I7260<= not G2844;
	I7264<= not G3252;
	I7269<= not G2851;
	I7272<= not G3253;
	I7276<= not G2861;
	I7280<= not G3208;
	I7284<= not G3255;
	I7288<= not G2873;
	I7291<= not G3212;
	I7295<= not G3260;
	I7300<= not G2883;
	I7303<= not G3262;
	I7308<= not G3070;
	I7311<= not G2803;
	I7315<= not G2891;
	I7318<= not G3266;
	I7330<= not G3761;
	I7333<= not G3729;
	I7336<= not G3997;
	I7339<= not G4004;
	I7342<= not G4011;
	I7345<= not G4050;
	I7348<= not G4056;
	I7351<= not G4061;
	I7354<= not G4066;
	I7357<= not G4077;
	I7360<= not G4081;
	I7363<= not G4005;
	I7366<= not G4012;
	I7369<= not G4051;
	I7372<= not G4057;
	I7375<= not G4062;
	I7378<= not G4067;
	I7381<= not G4078;
	I7384<= not G4082;
	I7387<= not G4083;
	I7390<= not G4087;
	I7393<= not G4096;
	I7396<= not G4102;
	I7399<= not G4113;
	I7402<= not G4121;
	I7405<= not G3861;
	I7408<= not G4125;
	I7411<= not G4140;
	I7414<= not G4156;
	I7417<= not G4160;
	I7420<= not G4167;
	I7423<= not G3331;
	I7426<= not G3334;
	I7429<= not G3344;
	I7432<= not G3663;
	I7435<= not G3459;
	I7438<= not G3461;
	I7441<= not G3473;
	I7444<= not G3683;
	I7447<= not G3694;
	I7450<= not G3704;
	I7453<= not G3708;
	I7456<= not G3716;
	I7459<= not G3720;
	I7462<= not G3721;
	I7465<= not G3726;
	I7468<= not G3697;
	I7478<= not G3566;
	I7487<= not G3371;
	I7509<= not G3566;
	I7513<= not G4144;
	I7523<= not G4095;
	I7536<= not G4098;
	I7546<= not G4105;
	I7556<= not G4080;
	I7559<= not G4116;
	I7577<= not G4124;
	I7586<= not G4127;
	I7593<= not G4142;
	I7600<= not G4159;
	I7606<= not G4166;
	I7612<= not G3817;
	I7625<= not G4164;
	I7630<= not G3524;
	I7633<= not G3474;
	I7636<= not G3330;
	I7639<= not G3722;
	I7642<= not G3440;
	I7648<= not G3727;
	I7651<= not G3332;
	I7654<= not G3728;
	I7659<= not G3731;
	I7662<= not G3336;
	I7665<= not G3732;
	I7668<= not G3733;
	I7671<= not G3351;
	I7674<= not G3352;
	I7677<= not G3735;
	I7680<= not G3736;
	I7691<= not G3363;
	I7694<= not G3742;
	I7697<= not G3743;
	I7701<= not G3513;
	I7707<= not G3370;
	I7710<= not G3749;
	I7713<= not G3750;
	I7716<= not G3751;
	I7719<= not G3752;
	I7726<= not G3378;
	I7729<= not G3757;
	I7732<= not G3758;
	I7735<= not G3759;
	I7743<= not G3762;
	I7746<= not G3763;
	I7749<= not G3764;
	I7752<= not G3407;
	I7757<= not G3767;
	I7760<= not G3768;
	I7763<= not G3769;
	I7766<= not G3770;
	I7771<= not G3418;
	I7776<= not G3773;
	I7779<= not G3774;
	I7782<= not G3775;
	I7790<= not G3782;
	I7793<= not G3783;
	I7800<= not G3791;
	I7803<= not G3820;
	I7810<= not G3799;
	I7817<= not G3399;
	I7820<= not G3811;
	I7825<= not G3414;
	I7829<= not G3425;
	I7833<= not G3585;
	I7837<= not G4158;
	I7840<= not G3431;
	I7843<= not G3440;
	I7847<= not G3435;
	I7852<= not G3438;
	I7858<= not G3631;
	I7886<= not G4076;
	I7889<= not G3373;
	I7899<= not G3380;
	I7906<= not G3907;
	I7909<= not G3387;
	I7916<= not G3664;
	I7920<= not G3440;
	I7923<= not G3394;
	I7931<= not G3624;
	I7935<= not G3440;
	I7938<= not G3406;
	I7946<= not G3417;
	I7952<= not G3664;
	I7956<= not G3428;
	I7964<= not G3433;
	I7973<= not G3437;
	I7984<= not G3621;
	I7996<= not G3462;
	I7999<= not G4114;
	I8004<= not G3967;
	I8007<= not G3829;
	I8011<= not G3820;
	I8024<= not G4117;
	I8031<= not G3540;
	I8036<= not G3820;
	I8039<= not G3506;
	I8050<= not G4089;
	I8061<= not G3381;
	I8080<= not G3538;
	I8085<= not G3664;
	I8089<= not G3545;
	I8098<= not G3583;
	I8109<= not G3622;
	I8116<= not G3627;
	I8123<= not G3630;
	I8126<= not G3662;
	I8133<= not G3632;
	I8136<= not G4144;
	I8139<= not G3681;
	I8147<= not G3633;
	I8154<= not G3636;
	I8161<= not G3637;
	I8164<= not G3566;
	I8192<= not G3566;
	I8199<= not G4013;
	I8204<= not G3976;
	I8211<= not G3566;
	I8215<= not G3981;
	I8228<= not G4468;
	I8231<= not G4170;
	I8234<= not G4232;
	I8237<= not G4295;
	I8240<= not G4380;
	I8247<= not G4615;
	I8250<= not G4589;
	I8253<= not G4637;
	I8256<= not G4711;
	I8259<= not G4590;
	I8262<= not G4636;
	I8265<= not G4602;
	I8268<= not G4674;
	I8275<= not G4351;
	I8278<= not G4495;
	I8282<= not G4770;
	I8285<= not G4771;
	I8290<= not G4778;
	I8293<= not G4779;
	I8298<= not G4437;
	I8303<= not G4784;
	I8308<= not G4443;
	I8311<= not G4794;
	I8315<= not G4788;
	I8320<= not G4452;
	I8324<= not G4794;
	I8328<= not G4801;
	I8333<= not G4456;
	I8337<= not G4352;
	I8340<= not G4804;
	I8351<= not G4794;
	I8358<= not G4794;
	I8379<= not G4231;
	I8385<= not G4238;
	I8388<= not G4239;
	I8396<= not G4255;
	I8403<= not G4264;
	I8406<= not G4274;
	I8410<= not G4283;
	I8414<= not G4293;
	I8418<= not G4794;
	I8421<= not G4309;
	I8429<= not G4458;
	I8436<= not G4462;
	I8442<= not G4464;
	I8449<= not G4469;
	I8456<= not G4472;
	I8462<= not G4475;
	I8465<= not G4807;
	I8473<= not G4577;
	I8476<= not G4577;
	I8487<= not G4526;
	I8490<= not G4526;
	I8495<= not G4325;
	I8499<= not G4330;
	I8503<= not G4445;
	I8506<= not G4334;
	I8520<= not G4338;
	I8535<= not G4340;
	I8551<= not G4342;
	I8611<= not G4562;
	I8614<= not G4414;
	I8631<= not G4425;
	I8647<= not G4219;
	I8711<= not G4530;
	I8724<= not G4791;
	I8811<= not G4465;
	I8815<= not G4471;
	I8820<= not G4473;
	I8827<= not G4477;
	I8831<= not G4480;
	I8835<= not G4791;
	I8839<= not G4484;
	I8842<= not G4556;
	I8848<= not G4490;
	I8851<= not G4498;
	I8854<= not G4500;
	I8858<= not G4506;
	I8865<= not G4518;
	I8869<= not G4421;
	I8872<= not G4529;
	I8877<= not G4421;
	I8880<= not G4537;
	I8885<= not G4548;
	I8889<= not G4553;
	I8892<= not G4554;
	I8900<= not G4560;
	I8903<= not G4561;
	I8911<= not G4565;
	I8919<= not G4576;
	I8929<= not G4582;
	I8934<= not G4271;
	I8943<= not G4585;
	I8967<= not G4482;
	I8973<= not G4488;
	I8982<= not G4728;
	I8985<= not G4733;
	I8989<= not G4746;
	I8996<= not G4757;
	I9001<= not G4762;
	I9013<= not G4767;
	I9016<= not G4722;
	I9020<= not G4773;
	I9023<= not G4727;
	I9029<= not G4781;
	I9032<= not G4732;
	I9040<= not G4794;
	I9043<= not G4786;
	I9046<= not G4736;
	I9053<= not G4752;
	I9056<= not G4753;
	I9062<= not G4759;
	I9065<= not G4760;
	I9068<= not G4768;
	I9074<= not G4764;
	I9077<= not G4765;
	I9080<= not G4775;
	I9084<= not G4886;
	I9087<= not G5113;
	I9090<= not G5567;
	I9093<= not G5397;
	I9096<= not G5568;
	I9099<= not G5572;
	I9102<= not G5586;
	I9105<= not G5589;
	I9108<= not G5593;
	I9111<= not G5596;
	I9114<= not G5603;
	I9117<= not G5615;
	I9120<= not G5218;
	I9123<= not G4890;
	I9126<= not G4891;
	I9129<= not G4892;
	I9132<= not G4893;
	I9135<= not G5198;
	I9138<= not G5210;
	I9141<= not G5402;
	I9144<= not G5007;
	I9147<= not G5011;
	I9150<= not G5012;
	I9153<= not G5027;
	I9156<= not G5032;
	I9159<= not G5033;
	I9162<= not G5035;
	I9165<= not G5037;
	I9168<= not G5040;
	I9171<= not G4902;
	I9174<= not G4903;
	I9177<= not G4904;
	I9180<= not G4905;
	I9185<= not G4915;
	I9188<= not G4908;
	I9191<= not G5546;
	I9194<= not G5236;
	I9199<= not G4935;
	I9202<= not G4915;
	I9205<= not G5309;
	I9208<= not G5047;
	I9213<= not G4944;
	I9216<= not G4935;
	I9221<= not G5236;
	I9224<= not G5063;
	I9229<= not G4954;
	I9232<= not G4944;
	I9237<= not G5205;
	I9240<= not G5069;
	I9243<= not G5245;
	I9248<= not G4954;
	I9253<= not G5052;
	I9256<= not G5078;
	I9259<= not G5301;
	I9265<= not G5085;
	I9268<= not G5305;
	I9273<= not G5091;
	I9276<= not G5241;
	I9279<= not G5314;
	I9282<= not G5633;
	I9287<= not G5576;
	I9290<= not G5052;
	I9293<= not G5486;
	I9296<= not G4908;
	I9302<= not G5576;
	I9305<= not G4970;
	I9308<= not G5494;
	I9311<= not G4915;
	I9317<= not G5576;
	I9320<= not G5013;
	I9323<= not G5620;
	I9326<= not G5320;
	I9329<= not G5504;
	I9332<= not G4935;
	I9338<= not G5576;
	I9341<= not G5013;
	I9346<= not G5281;
	I9349<= not G5515;
	I9352<= not G4944;
	I9359<= not G5576;
	I9362<= not G5013;
	I9365<= not G5392;
	I9368<= not G5288;
	I9371<= not G5075;
	I9377<= not G5576;
	I9380<= not G5013;
	I9383<= not G5296;
	I9388<= not G5576;
	I9391<= not G5013;
	I9394<= not G5195;
	I9399<= not G5013;
	I9402<= not G5107;
	I9409<= not G5013;
	I9415<= not G5047;
	I9421<= not G5063;
	I9424<= not G4963;
	I9427<= not G4963;
	I9433<= not G5069;
	I9440<= not G5078;
	I9443<= not G5557;
	I9446<= not G5052;
	I9452<= not G5085;
	I9458<= not G5091;
	I9461<= not G4940;
	I9475<= not G5445;
	I9479<= not G4954;
	I9483<= not G5050;
	I9486<= not G5066;
	I9491<= not G5072;
	I9498<= not G5081;
	I9505<= not G5088;
	I9510<= not G5421;
	I9514<= not G5094;
	I9519<= not G4998;
	I9525<= not G5001;
	I9531<= not G5004;
	I9536<= not G5008;
	I9539<= not G5354;
	I9544<= not G5024;
	I9550<= not G5030;
	I9564<= not G5109;
	I9567<= not G5556;
	I9571<= not G5509;
	I9581<= not G5111;
	I9585<= not G5241;
	I9588<= not G5114;
	I9591<= not G5095;
	I9594<= not G5083;
	I9598<= not G5120;
	I9602<= not G5013;
	I9605<= not G5620;
	I9608<= not G5127;
	I9612<= not G5149;
	I9617<= not G5405;
	I9620<= not G5189;
	I9625<= not G5405;
	I9632<= not G5557;
	I9639<= not G5126;
	I9642<= not G5229;
	I9647<= not G5148;
	I9652<= not G5426;
	I9655<= not G5173;
	I9658<= not G5150;
	I9662<= not G5319;
	I9665<= not G5174;
	I9669<= not G5426;
	I9673<= not G5182;
	I9677<= not G5190;
	I9680<= not G5194;
	I9684<= not G5426;
	I9688<= not G5201;
	I9695<= not G5212;
	I9699<= not G5426;
	I9706<= not G5221;
	I9712<= not G5230;
	I9717<= not G5426;
	I9720<= not G5248;
	I9727<= not G5250;
	I9731<= not G5255;
	I9734<= not G5257;
	I9737<= not G5258;
	I9744<= not G5263;
	I9749<= not G5266;
	I9754<= not G5271;
	I9759<= not G5344;
	I9762<= not G5276;
	I9766<= not G5348;
	I9769<= not G5287;
	I9773<= not G4934;
	I9776<= not G5353;
	I9779<= not G5391;
	I9783<= not G5395;
	I9786<= not G5396;
	I9789<= not G5401;
	I9792<= not G5403;
	I9795<= not G5404;
	I9798<= not G5415;
	I9801<= not G5416;
	I9804<= not G5417;
	I9807<= not G5419;
	I9810<= not G5576;
	I9813<= not G5241;
	I9816<= not G5576;
	I9822<= not G5219;
	I9826<= not G5390;
	I9829<= not G5013;
	I9833<= not G5197;
	I9836<= not G5405;
	I9839<= not G5226;
	I9842<= not G5405;
	I9845<= not G5405;
	I9848<= not G5557;
	I9851<= not G5405;
	I9854<= not G5557;
	I9857<= not G5269;
	I9860<= not G5405;
	I9863<= not G5557;
	I9866<= not G5274;
	I9869<= not G5405;
	I9872<= not G5557;
	I9875<= not G5278;
	I9880<= not G5405;
	I9883<= not G5557;
	I9886<= not G5286;
	I9893<= not G5557;
	I9896<= not G5295;
	I9901<= not G5557;
	I9905<= not G5300;
	I9915<= not G5304;
	I9923<= not G5308;
	I9930<= not G5317;
	I9935<= not G5477;
	I9938<= not G5478;
	I9953<= not G5484;
	I9956<= not G5485;
	I9965<= not G5493;
	I9973<= not G5502;
	I9981<= not G5514;
	I9984<= not G5529;
	I9988<= not G5526;
	I9992<= not G5633;
	I9995<= not G5536;
	I10003<= not G4908;
	I10006<= not G5633;
	I10009<= not G5542;
	I10012<= not G5543;
	I10015<= not G5641;
	I10018<= not G5862;
	I10021<= not G5692;
	I10024<= not G5700;
	I10027<= not G5751;
	I10030<= not G5685;
	I10033<= not G5693;
	I10036<= not G5701;
	I10039<= not G5718;
	I10042<= not G5723;
	I10045<= not G5727;
	I10048<= not G5734;
	I10051<= not G5702;
	I10054<= not G5728;
	I10057<= not G5741;
	I10060<= not G5752;
	I10063<= not G5766;
	I10066<= not G5778;
	I10069<= not G5787;
	I10072<= not G5719;
	I10075<= not G5724;
	I10078<= not G5729;
	I10081<= not G5735;
	I10084<= not G5742;
	I10087<= not G5753;
	I10090<= not G5767;
	I10093<= not G5779;
	I10096<= not G5794;
	I10099<= not G5800;
	I10102<= not G5730;
	I10105<= not G5736;
	I10108<= not G5743;
	I10111<= not G5754;
	I10114<= not G5768;
	I10117<= not G6241;
	I10120<= not G6248;
	I10123<= not G5676;
	I10126<= not G5682;
	I10129<= not G5688;
	I10132<= not G5696;
	I10135<= not G6249;
	I10138<= not G5677;
	I10141<= not G5683;
	I10144<= not G5689;
	I10147<= not G5697;
	I10150<= not G5705;
	I10153<= not G5947;
	I10156<= not G6100;
	I10159<= not G5936;
	I10162<= not G5943;
	I10165<= not G5948;
	I10168<= not G5982;
	I10171<= not G5992;
	I10174<= not G5994;
	I10177<= not G6103;
	I10180<= not G6107;
	I10183<= not G6108;
	I10186<= not G6110;
	I10189<= not G6112;
	I10192<= not G6115;
	I10195<= not G6116;
	I10198<= not G6118;
	I10201<= not G5998;
	I10204<= not G6031;
	I10221<= not G6117;
	I10228<= not G6113;
	I10231<= not G6111;
	I10234<= not G6114;
	I10237<= not G6120;
	I10240<= not G5937;
	I10243<= not G5918;
	I10248<= not G6125;
	I10251<= not G6126;
	I10258<= not G6134;
	I10274<= not G5811;
	I10278<= not G5815;
	I10282<= not G6163;
	I10286<= not G6237;
	I10289<= not G6003;
	I10293<= not G5863;
	I10296<= not G6242;
	I10299<= not G6243;
	I10302<= not G6179;
	I10305<= not G6180;
	I10308<= not G6003;
	I10314<= not G6251;
	I10317<= not G6003;
	I10322<= not G6193;
	I10325<= not G6003;
	I10331<= not G6198;
	I10334<= not G6003;
	I10340<= not G6205;
	I10343<= not G6003;
	I10349<= not G6215;
	I10352<= not G6216;
	I10355<= not G6003;
	I10362<= not G6224;
	I10367<= not G6234;
	I10370<= not G5857;
	I10374<= not G5852;
	I10378<= not G6244;
	I10381<= not G5847;
	I10384<= not G5842;
	I10388<= not G5830;
	I10391<= not G5838;
	I10394<= not G5824;
	I10398<= not G5820;
	I10412<= not G5821;
	I10421<= not G5826;
	I10427<= not G5839;
	I10434<= not G5843;
	I10437<= not G5755;
	I10445<= not G5770;
	I10456<= not G5844;
	I10461<= not G5849;
	I10477<= not G6049;
	I10484<= not G6155;
	I10495<= not G6144;
	I10499<= not G6149;
	I10503<= not G5858;
	I10514<= not G6154;
	I10526<= not G6161;
	I10531<= not G6169;
	I10535<= not G5867;
	I10538<= not G5910;
	I10541<= not G6176;
	I10546<= not G5914;
	I10549<= not G6184;
	I10553<= not G6192;
	I10557<= not G6197;
	I10560<= not G5887;
	I10563<= not G6043;
	I10566<= not G5904;
	I10573<= not G5980;
	I10584<= not G5864;
	I10589<= not G5763;
	I10592<= not G5865;
	I10598<= not G5874;
	I10601<= not G5996;
	I10607<= not G5763;
	I10610<= not G5879;
	I10613<= not G6000;
	I10620<= not G5884;
	I10623<= not G6002;
	I10630<= not G5889;
	I10633<= not G6015;
	I10639<= not G5830;
	I10643<= not G6026;
	I10648<= not G6030;
	I10651<= not G6035;
	I10655<= not G6036;
	I10659<= not G6038;
	I10663<= not G6040;
	I10666<= not G6042;
	I10671<= not G6045;
	I10678<= not G5777;
	I10682<= not G6051;
	I10685<= not G6054;
	I10689<= not G6059;
	I10693<= not G6068;
	I10698<= not G5856;
	I10702<= not G6071;
	I10706<= not G6080;
	I10710<= not G6088;
	I10713<= not G6003;
	I10716<= not G6093;
	I10719<= not G6003;
	I10724<= not G6096;
	I10729<= not G5935;
	I10733<= not G6099;
	I10736<= not G6104;
	I10739<= not G5942;
	I10753<= not G5814;
	I10756<= not G5810;
	I10759<= not G5803;
	I10762<= not G6127;
	I10789<= not G5867;
	I10795<= not G6123;
	I10801<= not G6536;
	I10804<= not G6388;
	I10807<= not G6396;
	I10810<= not G6539;
	I10813<= not G6397;
	I10816<= not G6406;
	I10819<= not G6706;
	I10822<= not G6584;
	I10825<= not G6588;
	I10828<= not G6708;
	I10831<= not G6710;
	I10834<= not G6715;
	I10837<= not G6717;
	I10840<= not G6719;
	I10843<= not G6723;
	I10846<= not G6729;
	I10849<= not G6734;
	I10852<= not G6751;
	I10855<= not G6685;
	I10858<= not G6688;
	I10861<= not G6694;
	I10864<= not G6634;
	I10873<= not G6331;
	I10885<= not G6332;
	I10888<= not G6333;
	I10891<= not G6334;
	I10898<= not G6735;
	I10901<= not G6620;
	I10904<= not G6558;
	I10907<= not G6705;
	I10910<= not G6703;
	I10914<= not G6728;
	I10917<= not G6732;
	I10920<= not G6733;
	I10924<= not G6736;
	I10927<= not G6755;
	I10937<= not G6552;
	I10941<= not G6555;
	I10946<= not G6548;
	I10949<= not G6747;
	I10952<= not G6556;
	I10958<= not G6559;
	I10963<= not G6793;
	I10966<= not G6561;
	I10971<= not G6344;
	I10974<= not G6563;
	I10979<= not G6565;
	I10984<= not G6757;
	I10991<= not G6759;
	I10996<= not G6786;
	I11005<= not G6386;
	I11008<= not G6795;
	I11011<= not G6340;
	I11021<= not G6398;
	I11024<= not G6399;
	I11029<= not G6485;
	I11034<= not G6629;
	I11037<= not G6629;
	I11043<= not G6412;
	I11046<= not G6635;
	I11049<= not G6635;
	I11055<= not G6419;
	I11058<= not G6641;
	I11061<= not G6641;
	I11065<= not G6750;
	I11068<= not G6426;
	I11071<= not G6656;
	I11076<= not G6649;
	I11079<= not G6649;
	I11082<= not G6749;
	I11085<= not G6433;
	I11088<= not G6434;
	I11091<= not G6657;
	I11094<= not G6657;
	I11097<= not G6748;
	I11100<= not G6442;
	I11103<= not G6667;
	I11106<= not G6667;
	I11109<= not G6464;
	I11112<= not G6445;
	I11115<= not G6462;
	I11119<= not G6461;
	I11122<= not G6450;
	I11127<= not G6452;
	I11132<= not G6451;
	I11135<= not G6679;
	I11140<= not G6448;
	I11143<= not G6446;
	I11146<= not G6439;
	I11149<= not G6468;
	I11152<= not G6469;
	I11155<= not G6470;
	I11159<= not G6478;
	I11162<= not G6479;
	I11166<= not G6480;
	I11169<= not G6481;
	I11173<= not G6500;
	I11176<= not G6501;
	I11180<= not G6506;
	I11183<= not G6507;
	I11188<= not G6513;
	I11191<= not G6514;
	I11194<= not G6515;
	I11198<= not G6521;
	I11201<= not G6522;
	I11204<= not G6523;
	I11207<= not G6524;
	I11211<= not G6527;
	I11214<= not G6528;
	I11217<= not G6529;
	I11222<= not G6533;
	I11225<= not G6534;
	I11228<= not G6471;
	I11232<= not G6537;
	I11235<= not G6538;
	I11238<= not G6543;
	I11249<= not G6541;
	I11252<= not G6542;
	I11255<= not G6547;
	I11269<= not G6545;
	I11272<= not G6546;
	I11275<= not G6502;
	I11286<= not G6551;
	I11289<= not G6508;
	I11293<= not G6516;
	I11296<= not G6525;
	I11299<= not G6727;
	I11303<= not G6526;
	I11306<= not G6731;
	I11309<= not G6531;
	I11312<= not G6488;
	I11315<= not G6644;
	I11318<= not G6488;
	I11322<= not G6652;
	I11326<= not G6660;
	I11330<= not G6571;
	I11333<= not G6670;
	I11338<= not G6680;
	I11342<= not G6686;
	I11345<= not G6692;
	I11348<= not G6695;
	I11351<= not G6698;
	I11354<= not G6553;
	I11357<= not G6594;
	I11360<= not G6351;
	I11363<= not G6595;
	I11367<= not G6392;
	I11383<= not G6385;
	I11387<= not G6672;
	I11391<= not G6387;
	I11394<= not G6621;
	I11397<= not G6713;
	I11405<= not G6627;
	I11408<= not G6405;
	I11412<= not G6411;
	I11417<= not G6638;
	I11420<= not G6417;
	I11423<= not G6488;
	I11427<= not G6573;
	I11433<= not G6424;
	I11436<= not G6488;
	I11440<= not G6577;
	I11444<= not G6653;
	I11447<= not G6431;
	I11450<= not G6488;
	I11456<= not G6440;
	I11459<= not G6488;
	I11464<= not G6443;
	I11467<= not G6488;
	I11472<= not G6488;
	I11477<= not G6488;
	I11483<= not G6567;
	I11489<= not G6569;
	I11494<= not G6574;
	I11498<= not G6578;
	I11501<= not G6581;
	I11505<= not G6585;
	I11515<= not G6589;
	I11519<= not G6591;
	I11524<= not G6593;
	I11528<= not G6796;
	I11531<= not G7126;
	I11534<= not G6917;
	I11537<= not G7144;
	I11540<= not G6877;
	I11543<= not G6881;
	I11560<= not G7037;
	I11563<= not G6819;
	I11566<= not G6820;
	I11569<= not G6821;
	I11572<= not G6822;
	I11575<= not G6823;
	I11578<= not G6824;
	I11581<= not G6826;
	I11584<= not G6827;
	I11587<= not G6828;
	I11590<= not G6829;
	I11593<= not G6830;
	I11596<= not G6831;
	I11599<= not G6832;
	I11602<= not G6833;
	I11605<= not G6834;
	I11608<= not G6903;
	I11611<= not G6913;
	I11614<= not G6838;
	I11617<= not G6839;
	I11620<= not G6840;
	I11623<= not G6841;
	I11626<= not G7042;
	I11629<= not G6914;
	I11632<= not G6931;
	I11635<= not G6947;
	I11638<= not G6948;
	I11641<= not G6960;
	I11644<= not G6970;
	I11647<= not G6925;
	I11650<= not G6938;
	I11653<= not G6954;
	I11656<= not G7122;
	I11659<= not G7097;
	I11662<= not G7033;
	I11665<= not G7038;
	I11668<= not G7043;
	I11671<= not G7047;
	I11674<= not G7051;
	I11677<= not G7056;
	I11680<= not G7064;
	I11683<= not G7069;
	I11686<= not G7039;
	I11689<= not G7044;
	I11692<= not G7048;
	I11695<= not G7052;
	I11698<= not G7057;
	I11701<= not G7065;
	I11704<= not G7008;
	I11707<= not G7009;
	I11710<= not G7020;
	I11713<= not G7023;
	I11716<= not G7026;
	I11719<= not G7029;
	I11722<= not G7034;
	I11725<= not G7040;
	I11728<= not G7010;
	I11731<= not G7021;
	I11734<= not G7024;
	I11737<= not G7027;
	I11740<= not G7030;
	I11743<= not G7035;
	I11746<= not G6857;
	I11752<= not G7032;
	I11756<= not G7191;
	I11759<= not G7244;
	I11767<= not G7201;
	I11770<= not G7202;
	I11773<= not G7257;
	I11778<= not G7210;
	I11783<= not G7246;
	I11786<= not G7246;
	I11790<= not G7246;
	I11794<= not G7188;
	I11797<= not G6852;
	I11800<= not G7246;
	I11804<= not G7190;
	I11807<= not G6854;
	I11810<= not G7246;
	I11814<= not G7196;
	I11817<= not G7246;
	I11821<= not G7205;
	I11824<= not G7246;
	I11829<= not G7213;
	I11833<= not G7077;
	I11836<= not G7220;
	I11841<= not G7226;
	I11845<= not G6869;
	I11858<= not G6888;
	I11869<= not G6894;
	I11873<= not G6863;
	I11879<= not G6893;
	I11882<= not G6895;
	I11889<= not G6898;
	I11898<= not G6896;
	I11901<= not G6897;
	I11904<= not G6902;
	I11921<= not G6904;
	I11926<= not G6900;
	I11929<= not G6901;
	I11932<= not G6908;
	I11942<= not G6909;
	I11947<= not G6905;
	I11950<= not G6906;
	I11953<= not G6907;
	I11956<= not G6912;
	I11961<= not G7053;
	I11964<= not G6910;
	I11967<= not G6911;
	I11970<= not G6918;
	I11989<= not G6919;
	I11992<= not G7058;
	I12009<= not G6915;
	I12012<= not G6916;
	I12015<= not G6924;
	I12026<= not G7119;
	I12029<= not G6922;
	I12032<= not G6923;
	I12035<= not G6930;
	I12053<= not G6928;
	I12056<= not G6929;
	I12081<= not G6934;
	I12099<= not G7258;
	I12103<= not G6859;
	I12120<= not G7106;
	I12123<= not G6861;
	I12133<= not G6870;
	I12150<= not G7074;
	I12153<= not G6874;
	I12156<= not G6878;
	I12159<= not G7243;
	I12162<= not G7146;
	I12165<= not G6882;
	I12168<= not G7256;
	I12171<= not G6885;
	I12174<= not G6939;
	I12177<= not G7259;
	I12180<= not G7263;
	I12183<= not G7007;
	I12186<= not G7264;
	I12190<= not G7268;
	I12193<= not G7270;
	I12196<= not G7272;
	I12199<= not G7278;
	I12202<= not G6983;
	I12205<= not G6993;
	I12208<= not G7124;
	I12223<= not G7049;
	I12226<= not G7066;
	I12229<= not G7070;
	I12232<= not G7072;
	I12235<= not G7082;
	I12239<= not G7073;
	I12242<= not G7089;
	I12245<= not G7093;
	I12248<= not G7098;
	I12251<= not G7076;
	I12255<= not G7203;
	I12258<= not G7103;
	I12261<= not G7078;
	I12265<= not G7211;
	I12268<= not G7107;
	I12271<= not G7218;
	I12274<= not G7110;
	I12279<= not G7225;
	I12282<= not G7113;
	I12286<= not G7231;
	I12289<= not G7142;
	I12293<= not G7116;
	I12296<= not G7236;
	I12300<= not G7240;
	I12303<= not G7242;
	I12307<= not G7245;
	I12318<= not G6862;
	I12322<= not G7246;
	I12326<= not G7246;
	I12335<= not G7133;
	I12339<= not G7054;
	I12344<= not G7062;
	I12354<= not G7143;
	I12357<= not G7147;
	I12360<= not G7183;
	I12363<= not G7187;
	I12366<= not G7134;
	I12369<= not G7189;
	I12372<= not G7137;
	I12376<= not G7195;
	I12380<= not G7204;
	I12384<= not G7212;
	I12388<= not G7219;
	I12397<= not G7284;
	I12400<= not G7537;
	I12403<= not G7611;
	I12406<= not G7464;
	I12409<= not G7501;
	I12412<= not G7520;
	I12415<= not G7631;
	I12418<= not G7568;
	I12421<= not G7634;
	I12424<= not G7635;
	I12427<= not G7636;
	I12430<= not G7649;
	I12433<= not G7657;
	I12436<= not G7659;
	I12439<= not G7663;
	I12442<= not G7672;
	I12445<= not G7521;
	I12448<= not G7530;
	I12451<= not G7538;
	I12454<= not G7544;
	I12457<= not G7559;
	I12460<= not G7569;
	I12463<= not G7579;
	I12466<= not G7585;
	I12469<= not G7531;
	I12472<= not G7539;
	I12475<= not G7545;
	I12478<= not G7560;
	I12481<= not G7570;
	I12484<= not G7580;
	I12487<= not G7723;
	I12490<= not G7637;
	I12493<= not G7650;
	I12496<= not G7724;
	I12499<= not G7725;
	I12502<= not G7726;
	I12505<= not G7728;
	I12508<= not G7731;
	I12511<= not G7733;
	I12514<= not G7735;
	I12517<= not G7737;
	I12520<= not G7415;
	I12523<= not G7421;
	I12526<= not G7648;
	I12529<= not G7589;
	I12532<= not G7594;
	I12535<= not G7656;
	I12538<= not G7658;
	I12541<= not G7662;
	I12544<= not G7669;
	I12547<= not G7673;
	I12550<= not G7675;
	I12553<= not G7676;
	I12556<= not G7678;
	I12559<= not G7477;
	I12562<= not G7377;
	I12565<= not G7388;
	I12568<= not G7502;
	I12571<= not G7509;
	I12574<= not G7522;
	I12577<= not G7532;
	I12580<= not G7540;
	I12583<= not G7546;
	I12586<= not G7561;
	I12589<= not G7571;
	I12592<= not G7445;
	I12595<= not G7706;
	I12598<= not G7628;
	I12601<= not G7629;
	I12604<= not G7630;
	I12607<= not G7633;
	I12610<= not G7627;
	I12613<= not G7525;
	I12616<= not G7534;
	I12627<= not G7697;
	I12631<= not G7705;
	I12634<= not G7727;
	I12638<= not G7708;
	I12641<= not G7709;
	I12644<= not G7729;
	I12647<= not G7711;
	I12652<= not G7458;
	I12655<= not G7402;
	I12678<= not G7376;
	I12683<= not G7387;
	I12690<= not G7555;
	I12694<= not G7374;
	I12712<= not G7441;
	I12751<= not G7626;
	I12759<= not G7702;
	I12762<= not G7541;
	I12765<= not G7638;
	I12770<= not G7638;
	I12773<= not G7581;
	I12776<= not G7586;
	I12779<= not G7608;
	I12783<= not G7590;
	I12786<= not G7622;
	I12790<= not G7618;
	I12793<= not G7619;
	I12796<= not G7543;
	I12799<= not G7556;
	I12805<= not G7684;
	I12809<= not G7686;
	I12813<= not G7688;
	I12817<= not G7692;
	I12822<= not G7677;
	I12825<= not G7696;
	I12829<= not G7680;
	I12832<= not G7681;
	I12835<= not G7660;
	I12838<= not G7682;
	I12843<= not G7683;
	I12846<= not G7685;
	I12849<= not G7632;
	I12853<= not G7638;
	I12857<= not G7638;
	I12862<= not G7638;
	I12867<= not G7638;
	I12871<= not G7638;
	I12875<= not G7638;
	I12878<= not G7638;
	I12901<= not G7984;
	I12904<= not G7985;
	I12907<= not G7959;
	I12910<= not G7922;
	I12913<= not G7845;
	I12916<= not G7849;
	I12919<= not G8003;
	I12930<= not G7896;
	I12933<= not G7899;
	I12936<= not G7983;
	I12939<= not G7977;
	I12942<= not G7982;
	I12948<= not G8019;
	I12953<= not G8024;
	I12971<= not G8039;
	I12978<= not G8040;
	I12981<= not G8041;
	I12986<= not G8042;
	I12989<= not G8043;
	I12993<= not G8044;
	I12999<= not G7844;
	I13002<= not G8045;
	I13005<= not G8046;
	I13010<= not G8047;
	I13013<= not G8048;
	I13017<= not G7848;
	I13020<= not G8049;
	I13023<= not G8050;
	I13027<= not G8051;
	I13030<= not G8052;
	I13036<= not G8053;
	I13039<= not G8054;
	I13043<= not G8055;
	I13048<= not G8059;
	I13051<= not G8060;
	I13057<= not G7843;
	I13068<= not G7906;
	I13083<= not G7921;
	I13086<= not G7924;
	I13096<= not G7925;
	I13099<= not G7927;
	I13102<= not G7928;
	I13105<= not G7929;
	I13109<= not G7981;
	I13114<= not G7930;
	I13117<= not G7904;
	I13122<= not G7966;
	I13125<= not G7975;
	I13128<= not G7976;
	I13131<= not G7979;
	I13166<= not G8009;
	I13185<= not G8192;
	I13188<= not G8171;
	I13191<= not G8132;
	I13194<= not G8140;
	I13197<= not G8186;
	I13200<= not G8251;
	I13203<= not G8196;
	I13206<= not G8197;
	I13209<= not G8198;
	I13212<= not G8195;
	I13224<= not G8261;
	I13227<= not G8264;
	I13230<= not G8244;
	I13233<= not G8265;
	I13236<= not G8245;
	I13239<= not G8266;
	I13242<= not G8267;
	I13245<= not G8269;
	I13255<= not G8270;
	I13280<= not G8250;
	I13290<= not G8254;
	I13314<= not G8260;
	I13317<= not G8093;
	I13320<= not G8096;
	I13323<= not G8203;
	I13326<= not G8203;
	I13329<= not G8116;
	I13332<= not G8206;
	I13335<= not G8206;
	I13338<= not G8210;
	I13341<= not G8210;
	I13344<= not G8121;
	I13347<= not G8122;
	I13351<= not G8214;
	I13354<= not G8214;
	I13357<= not G8125;
	I13360<= not G8126;
	I13364<= not G8221;
	I13367<= not G8221;
	I13370<= not G8128;
	I13373<= not G8226;
	I13376<= not G8226;
	I13379<= not G8133;
	I13382<= not G8134;
	I13385<= not G8230;
	I13388<= not G8230;
	I13391<= not G8178;
	I13394<= not G8137;
	I13397<= not G8138;
	I13400<= not G8236;
	I13403<= not G8236;
	I13406<= not G8179;
	I13409<= not G8141;
	I13412<= not G8142;
	I13415<= not G8144;
	I13418<= not G8145;
	I13421<= not G8200;
	I13424<= not G8200;
	I13427<= not G8241;
	I13430<= not G8241;
	I13433<= not G8181;
	I13436<= not G8187;
	I13439<= not G8187;
	I13442<= not G8182;
	I13445<= not G8149;
	I13448<= not G8150;
	I13451<= not G8152;
	I13454<= not G8183;
	I13457<= not G8184;
	I13460<= not G8155;
	I13463<= not G8156;
	I13466<= not G8160;
	I13469<= not G8147;
	I13475<= not G8173;
	I13478<= not G8191;
	I13482<= not G8193;
	I13485<= not G8194;
	I13489<= not G8233;
	I13568<= not G8343;
	I13571<= not G8355;
	I13574<= not G8360;
	I13577<= not G8330;
	I13580<= not G8338;
	I13583<= not G8344;
	I13586<= not G8356;
	I13589<= not G8361;
	I13592<= not G8362;
	I13595<= not G8339;
	I13606<= not G8311;
	I13609<= not G8312;
	I13612<= not G8325;
	I13615<= not G8333;
	I13618<= not G8345;
	I13621<= not G8315;
	I13624<= not G8320;
	I13627<= not G8326;
	I13630<= not G8334;
	I13633<= not G8346;
	I13636<= not G8357;
	I13639<= not G8321;
	I13642<= not G8378;
	I13645<= not G8379;
	I13648<= not G8376;
	I13666<= not G8292;
	I13669<= not G8294;
	I13674<= not G8304;
	I13678<= not G8306;
	I13682<= not G8310;
	I13695<= not G8363;
	I13708<= not G8337;
	I13711<= not G8342;
	I13714<= not G8351;
	I13717<= not G8354;
	I13720<= not G8358;
	I13723<= not G8359;
	I13726<= not G8375;
	I13729<= not G8290;
	I13732<= not G8291;
	I13735<= not G8293;
	I13738<= not G8295;
	I13741<= not G8296;
	I13744<= not G8297;
	I13747<= not G8299;
	I13773<= not G8384;
	I13776<= not G8513;
	I13779<= not G8514;
	I13782<= not G8515;
	I13785<= not G8516;
	I13788<= not G8517;
	I13791<= not G8518;
	I13794<= not G8472;
	I13797<= not G8473;
	I13800<= not G8500;
	I13803<= not G8476;
	I13806<= not G8478;
	I13809<= not G8480;
	I13812<= not G8519;
	I13816<= not G8559;
	I13819<= not G8488;
	I13822<= not G8488;
	I13825<= not G8488;
	I13828<= not G8488;
	I13831<= not G8560;
	I13834<= not G8488;
	I13837<= not G8488;
	I13840<= not G8488;
	I13915<= not G8451;
	I13918<= not G8451;
	I13933<= not G8505;
	I13941<= not G8488;
	I13945<= not G8488;
	I13949<= not G8451;
	I13952<= not G8451;
	I13956<= not G8451;
	I13959<= not G8451;
	I13962<= not G8451;
	I13965<= not G8451;
	I13969<= not G8451;
	I13975<= not G8588;
	I13978<= not G8575;
	I14005<= not G8631;
	I14010<= not G8642;
	I14040<= not G8649;
	I14045<= not G8603;
	I14055<= not G8650;
	I14077<= not G8758;
	I14080<= not G8714;
	I14083<= not G8747;
	I14087<= not G8770;
	I14090<= not G8771;
	I14094<= not G8700;
	I14097<= not G8773;
	I14101<= not G8774;
	I14105<= not G8776;
	I14109<= not G8765;
	I14112<= not G8777;
	I14116<= not G8766;
	I14119<= not G8779;
	I14123<= not G8767;
	I14127<= not G8768;
	I14130<= not G8769;
	I14133<= not G8772;
	I14136<= not G8775;
	I14140<= not G8717;
	I14176<= not G8784;
	I14179<= not G8785;
	I14182<= not G8788;
	I14185<= not G8790;
	I14188<= not G8792;
	I14191<= not G8795;
	I14194<= not G8798;
	I14224<= not G8794;
	I14228<= not G8797;
	I14232<= not G8800;
	I14236<= not G8802;
	I14239<= not G8803;
	I14242<= not G8787;
	I14249<= not G8804;
	I14252<= not G8783;
	I14257<= not G8805;
	I14295<= not G8806;
	I14299<= not G8810;
	I14303<= not G8811;
	I14306<= not G8812;
	I14309<= not G8813;
	I14312<= not G8814;
	I14315<= not G8815;
	I14319<= not G8816;
	I14323<= not G8817;
	I14326<= not G8818;
	I14330<= not G8819;
	I14340<= not G8820;
	I14349<= not G8958;
	I14352<= not G8946;
	I14355<= not G8948;
	I14358<= not G8950;
	I14361<= not G8951;
	I14364<= not G8952;
	I14367<= not G8953;
	I14370<= not G8954;
	I14373<= not G8956;
	I14376<= not G8959;
	I14379<= not G8961;
	I14382<= not G8886;
	I14385<= not G8890;
	I14388<= not G8924;
	I14391<= not G8928;
	I14394<= not G8884;
	I14397<= not G8888;
	I14400<= not G8891;
	I14405<= not G8937;
	I14409<= not G8938;
	I14412<= not G8939;
	I14415<= not G8940;
	I14418<= not G8941;
	I14421<= not G8944;
	I14424<= not G8945;
	I14439<= not G8969;
	I14449<= not G8973;
	I14452<= not G8922;
	I14473<= not G8921;
	I14477<= not G8943;
	I14485<= not G8883;
	I14490<= not G8885;
	I14494<= not G8887;
	I14499<= not G8889;
	I14503<= not G8920;
	I14506<= not G8923;
	I14509<= not G8926;
	I14519<= not G9106;
	I14522<= not G9108;
	I14525<= not G9109;
	I14528<= not G9270;
	I14531<= not G9273;
	I14534<= not G9290;
	I14537<= not G9308;
	I14540<= not G9310;
	I14543<= not G9311;
	I14546<= not G9312;
	I14549<= not G9262;
	I14552<= not G9264;
	I14555<= not G9009;
	I14558<= not G9024;
	I14561<= not G9025;
	I14564<= not G9026;
	I14567<= not G9027;
	I14570<= not G9028;
	I14573<= not G9029;
	I14579<= not G9272;
	I14642<= not G9088;
	I14645<= not G9088;
	I14668<= not G9309;
	I14672<= not G9261;
	I14675<= not G9263;
	I14678<= not G9265;
	I14681<= not G9110;
	I14684<= not G9124;
	I14687<= not G9258;
	I14690<= not G9150;
	I14694<= not G9259;
	I14697<= not G9260;
	I14701<= not G9291;
	I14709<= not G9267;
	I14713<= not G9052;
	I14786<= not G9266;
	I14793<= not G9269;
	I14799<= not G9661;
	I14802<= not G9666;
	I14805<= not G9360;
	I14873<= not G9525;
	I14876<= not G9526;
	I14884<= not G9454;
	I14888<= not G9454;
	I14903<= not G9507;
	I14906<= not G9508;
	I14910<= not G9532;
	I14914<= not G9533;
	I14918<= not G9535;
	I14933<= not G9454;
	I14939<= not G9454;
	I14944<= not G9454;
	I14948<= not G9555;
	I14955<= not G9765;
	I14958<= not G9767;
	I14961<= not G9769;
	I14964<= not G9762;
	I14967<= not G9763;
	I14970<= not G9732;
	I14973<= not G9733;
	I14976<= not G9670;
	I14979<= not G9671;
	I14982<= not G9672;
	I14989<= not G9813;
	I15036<= not G9721;
	I15060<= not G9696;
	I15063<= not G9699;
	I15068<= not G9710;
	I15072<= not G9713;
	I15075<= not G9761;
	I15079<= not G9745;
	I15082<= not G9719;
	I15085<= not G9720;
	I15088<= not G9832;
	I15114<= not G9875;
	I15127<= not G9919;
	I15157<= not G9931;
	I15162<= not G9958;
	I15181<= not G9968;
	I15184<= not G9974;
	I15187<= not G9968;
	I15190<= not G9974;
	I15193<= not G9968;
	I15196<= not G9974;
	I15229<= not G9968;
	I15232<= not G9974;
	I15235<= not G9968;
	I15238<= not G9974;
	I15241<= not G10013;
	I15244<= not G10031;
	I15247<= not G10032;
	I15250<= not G9980;
	I15253<= not G9987;
	I15263<= not G9995;
	I15266<= not G10001;
	I15269<= not G9993;
	I15272<= not G10019;
	I15275<= not G9994;
	I15278<= not G10033;
	I15281<= not G10025;
	I15284<= not G10034;
	I15287<= not G9980;
	I15290<= not G9984;
	I15293<= not G10001;
	I15296<= not G9995;
	I15299<= not G9995;
	I15302<= not G10007;
	I15305<= not G10001;
	I15308<= not G10019;
	I15311<= not G10013;
	I15314<= not G10007;
	I15317<= not G10025;
	I15320<= not G10013;
	I15323<= not G10019;
	I15326<= not G10025;
	I15329<= not G9995;
	I15332<= not G10001;
	I15335<= not G10007;
	I15338<= not G10013;
	I15341<= not G10019;
	I15344<= not G10025;
	I15347<= not G9995;
	I15350<= not G10001;
	I15353<= not G10007;
	I15356<= not G10013;
	I15359<= not G10019;
	I15362<= not G9987;
	I15365<= not G10025;
	I15368<= not G9990;
	I15371<= not G9990;
	I15374<= not G10007;
	I15377<= not G10104;
	I15380<= not G10098;
	I15383<= not G10107;
	I15386<= not G10101;
	I15389<= not G10110;
	I15392<= not G10104;
	I15395<= not G10058;
	I15400<= not G10069;
	I15403<= not G10069;
	I15406<= not G10065;
	I15409<= not G10065;
	I15412<= not G10075;
	I15415<= not G10075;
	I15418<= not G10083;
	I15421<= not G10083;
	I15424<= not G10080;
	I15427<= not G10088;
	I15437<= not G10050;
	I15448<= not G10056;
	I15458<= not G10069;
	I15461<= not G10074;
	I15464<= not G10094;
	I15467<= not G10079;
	I15470<= not G10111;
	I15473<= not G10087;
	I15476<= not G10114;
	I15479<= not G10091;
	I15482<= not G10115;
	I15485<= not G10092;
	I15488<= not G10116;
	I15491<= not G10093;
	I15494<= not G10117;
	I15497<= not G10119;
	I15500<= not G10051;
	I15503<= not G10044;
	I15507<= not G10047;
	I15510<= not G10035;
	I15514<= not G10122;
	I15517<= not G10051;
	I15520<= not G10035;
	I15523<= not G10058;
	I15526<= not G10051;
	I15530<= not G10107;
	I15536<= not G10111;
	I15539<= not G10069;
	I15542<= not G10065;
	I15545<= not G10075;
	I15548<= not G10083;
	I15551<= not G10080;
	I15554<= not G10088;
	I15559<= not G10094;
	I15562<= not G10098;
	I15565<= not G10101;
	I15568<= not G10094;
	I15580<= not G10155;
	I15583<= not G10157;
	I15586<= not G10159;
	I15589<= not G10161;
	I15592<= not G10163;
	I15595<= not G10165;
	I15598<= not G10170;
	I15601<= not G10173;
	I15604<= not G10148;
	I15632<= not G10184;
	I15635<= not G10185;
	I15639<= not G10179;
	I15665<= not G10193;
	I15669<= not G10194;
	I15672<= not G10132;
	I15675<= not G10133;
	I15688<= not G10207;
	I15691<= not G10233;
	I15694<= not G10234;
	I15698<= not G10235;
	I15701<= not G10236;
	I15704<= not G10238;
	I15708<= not G10241;
	I15725<= not G10251;
	I15729<= not G10254;
	I15733<= not G10257;
	I15736<= not G10258;
	I15741<= not G10260;
	I15744<= not G10261;
	I15749<= not G10263;
	I15752<= not G10264;
	I15756<= not G10266;
	I15759<= not G10267;
	I15763<= not G10244;
	I15768<= not G10249;
	I15771<= not G10250;
	I15775<= not G10253;
	I15778<= not G10255;
	I15782<= not G10259;
	I15787<= not G10269;
	I15792<= not G10279;
	I15795<= not G10280;
	I15798<= not G10281;
	I15801<= not G10282;
	I15804<= not G10283;
	I15807<= not G10284;
	I15811<= not G10200;
	I15814<= not G10202;
	I15817<= not G10199;
	I15820<= not G10204;
	I15823<= not G10201;
	I15826<= not G10205;
	I15829<= not G10203;
	I15832<= not G10206;
	I15855<= not G10336;
	I15858<= not G10336;
	I15861<= not G10339;
	I15864<= not G10339;
	I15956<= not G10402;
	I15959<= not G10402;
	I15962<= not G10405;
	I15965<= not G10405;
	I15968<= not G10408;
	I15971<= not G10408;
	I15974<= not G10411;
	I15977<= not G10411;
	I15980<= not G10414;
	I15983<= not G10414;
	I15986<= not G10417;
	I15989<= not G10417;
	I16095<= not G10401;
	I16098<= not G10369;
	I16101<= not G10381;
	I16105<= not G10382;
	I16108<= not G10383;
	I16111<= not G10385;
	I16114<= not G10387;
	I16121<= not G10396;
	I16124<= not G10396;
	I16169<= not G10448;
	I16172<= not G10498;
	I16175<= not G10488;
	I16178<= not G10490;
	I16181<= not G10491;
	I16184<= not G10484;
	I16187<= not G10492;
	I16190<= not G10493;
	I16193<= not G10485;
	I16196<= not G10496;
	I16200<= not G10494;
	I16203<= not G10454;
	I16206<= not G10453;
	I16209<= not G10452;
	I16214<= not G10500;
	I16217<= not G10501;
	I16220<= not G10502;
	I16236<= not G10535;
	I16239<= not G10525;
	I16252<= not G10515;
	I16255<= not G10554;
	I16258<= not G10555;
	I16261<= not G10556;
	I16264<= not G10557;
	I16269<= not G10558;
	I16273<= not G10559;
	I16277<= not G10536;
	I16280<= not G10537;
	I16283<= not G10538;
	I16286<= not G10540;
	I16289<= not G10541;
	I16292<= not G10551;
	I16295<= not G10552;
	I16298<= not G10553;
	I16307<= not G10589;
	I16311<= not G10584;
	I16356<= not G10597;
	I16360<= not G10590;
	I16363<= not G10599;
	I16366<= not G10591;
	I16370<= not G10592;
	I16373<= not G10593;
	I16376<= not G10596;
	I16379<= not G10598;
	I16387<= not G10629;
	I16407<= not G10696;
	I16413<= not G10663;
	I16416<= not G10664;
	I16432<= not G10702;
	I16439<= not G10702;
	I16458<= not G10734;
	I16461<= not G10735;
	I16475<= not G10765;
	I16479<= not G10767;
	I16484<= not G10770;
	I16487<= not G10771;
	I16492<= not G10773;
	I16496<= not G10707;
	I16500<= not G10711;
	I16507<= not G10712;
	I16510<= not G10712;
	I16514<= not G10717;
	I16518<= not G10718;
	I16525<= not G10719;
	I16528<= not G10732;
	I16531<= not G10720;
	I16534<= not G10747;
	I16537<= not G10721;
	I16540<= not G10722;
	I16543<= not G10747;
	I16546<= not G10724;
	I16550<= not G10726;
	I16553<= not G10754;
	I16571<= not G10819;
	I16574<= not G10821;
	I16577<= not G10825;
	I16580<= not G10826;
	I16583<= not G10848;
	I16586<= not G10850;
	I16589<= not G10820;
	I16592<= not G10781;
	I16595<= not G10783;
	I16598<= not G10804;
	I16601<= not G10806;
	I16604<= not G10786;
	I16607<= not G10787;
	I16610<= not G10792;
	I16613<= not G10794;
	I16616<= not G10796;
	I16623<= not G10858;
	I16626<= not G10859;
	I16629<= not G10860;
	I16632<= not G10861;
	I16635<= not G10862;
	I16638<= not G10863;
	I16641<= not G10864;
	I16644<= not G10865;
	I16647<= not G10866;
	I16650<= not G10776;
	I16656<= not G10791;
	I16660<= not G10793;
	I16664<= not G10795;
	I16667<= not G10780;
	I16670<= not G10797;
	I16673<= not G10782;
	I16676<= not G10798;
	I16679<= not G10784;
	I16682<= not G10799;
	I16685<= not G10785;
	I16688<= not G10800;
	I16691<= not G10788;
	I16708<= not G10822;
	I16717<= not G10779;
	I16720<= not G10854;
	I16723<= not G10851;
	I16735<= not G10855;
	I16739<= not G10856;
	I16742<= not G10857;
	I16760<= not G10888;
	I16763<= not G10890;
	I16766<= not G10892;
	I16769<= not G10894;
	I16772<= not G10887;
	I16775<= not G10889;
	I16778<= not G10891;
	I16781<= not G10893;
	I16784<= not G10895;
	I16787<= not G10896;
	I16790<= not G10900;
	I16793<= not G11014;
	I16796<= not G11016;
	I16799<= not G11017;
	I16802<= not G10902;
	I16805<= not G10904;
	I16808<= not G10906;
	I16811<= not G10908;
	I16814<= not G10910;
	I16817<= not G10912;
	I16843<= not G10898;
	I16847<= not G10886;
	I16850<= not G10905;
	I16853<= not G10907;
	I16856<= not G10909;
	I16859<= not G10911;
	I16863<= not G10972;
	I16867<= not G10913;
	I16871<= not G10973;
	I16879<= not G10936;
	I16897<= not G10947;
	I16920<= not G11084;
	I16938<= not G11086;
	I16941<= not G11076;
	I16944<= not G11079;
	I16947<= not G11080;
	I16950<= not G11081;
	I16953<= not G11082;
	I16956<= not G11096;
	I16979<= not G11088;
	I16982<= not G11088;
	I17070<= not G11233;
	I17084<= not G11249;
	I17092<= not G11217;
	I17096<= not G11219;
	I17100<= not G11221;
	I17104<= not G11223;
	I17108<= not G11225;
	I17112<= not G11227;
	I17116<= not G11229;
	I17121<= not G11231;
	I17124<= not G11232;
	I17142<= not G11301;
	I17146<= not G11305;
	I17149<= not G11306;
	I17152<= not G11308;
	I17155<= not G11310;
	I17158<= not G11312;
	I17161<= not G11314;
	I17164<= not G11320;
	I17170<= not G11294;
	I17173<= not G11293;
	I17176<= not G11286;
	I17179<= not G11307;
	I17182<= not G11309;
	I17185<= not G11311;
	I17188<= not G11313;
	I17191<= not G11315;
	I17194<= not G11317;
	I17198<= not G11319;
	I17202<= not G11322;
	I17206<= not G11323;
	I17209<= not G11289;
	I17213<= not G11290;
	I17216<= not G11291;
	I17219<= not G11292;
	I17225<= not G11298;
	I17228<= not G11300;
	I17231<= not G11303;
	I17234<= not G11353;
	I17237<= not G11394;
	I17240<= not G11395;
	I17243<= not G11396;
	I17246<= not G11341;
	I17249<= not G11342;
	I17252<= not G11343;
	I17255<= not G11344;
	I17258<= not G11345;
	I17261<= not G11346;
	I17265<= not G11352;
	I17268<= not G11351;
	I17271<= not G11388;
	I17274<= not G11389;
	I17277<= not G11390;
	I17302<= not G11391;
	I17312<= not G11392;
	I17315<= not G11393;
	I17318<= not G11340;
	I17321<= not G11348;
	I17324<= not G11347;
	I17327<= not G11349;
	I17331<= not G11357;
	I17334<= not G11360;
	I17337<= not G11363;
	I17340<= not G11366;
	I17344<= not G11369;
	I17347<= not G11373;
	I17350<= not G11377;
	I17353<= not G11381;
	I17356<= not G11384;
	I17359<= not G11372;
	I17362<= not G11376;
	I17365<= not G11380;
	I17368<= not G11423;
	I17371<= not G11410;
	I17374<= not G11411;
	I17377<= not G11412;
	I17381<= not G11436;
	I17384<= not G11437;
	I17387<= not G11438;
	I17390<= not G11430;
	I17407<= not G11417;
	I17410<= not G11419;
	I17413<= not G11425;
	I17416<= not G11420;
	I17419<= not G11421;
	I17424<= not G11424;
	I17435<= not G11454;
	I17438<= not G11444;
	I17441<= not G11445;
	I17444<= not G11446;
	I17447<= not G11457;
	I17450<= not G11450;
	I17453<= not G11451;
	I17456<= not G11453;
	I17466<= not G11447;
	I17470<= not G11452;
	I17482<= not G11479;
	I17500<= not G11478;
	I17510<= not G11481;
	I17513<= not G11482;
	I17516<= not G11483;
	I17519<= not G11484;
	I17522<= not G11485;
	I17525<= not G11486;
	I17528<= not G11487;
	I17531<= not G11488;
	I17534<= not G11495;
	I17537<= not G11497;
	I17540<= not G11498;
	I17543<= not G11499;
	I17546<= not G11500;
	I17549<= not G11501;
	I17552<= not G11502;
	I17555<= not G11503;
	I17558<= not G11504;
	I17563<= not G11492;
	I17591<= not G11514;
	I17610<= not G11549;
	I17613<= not G11550;
	I17616<= not G11561;
	I17633<= not G11578;
	I17636<= not G11577;
	I17642<= not G11579;
	I17657<= not G11598;
	I17662<= not G11602;
	I17666<= not G11603;
	I17669<= not G11604;
	I17672<= not G11605;
	I17675<= not G11606;
	I17678<= not G11607;
	I17681<= not G11608;
	I17684<= not G11609;
	I17687<= not G11610;
	I17692<= not G11596;
	I17695<= not G11614;
	I17698<= not G11616;
	I17701<= not G11617;
	I17704<= not G11618;
	I17707<= not G11619;
	I17710<= not G11620;
	I17713<= not G11621;
	I17716<= not G11622;
	I17719<= not G11623;
	I17724<= not G11625;
	I17730<= not G11638;
	I17733<= not G11639;
	I17736<= not G11640;
	I17739<= not G11641;
	I17742<= not G11636;
	I17746<= not G11643;
	I17749<= not G11644;
	I17752<= not G11645;
	I17755<= not G11646;
	I17758<= not G11647;
	I17761<= not G11652;
	I17764<= not G11651;
	I17767<= not G11648;
	I17770<= not G11649;
	I17773<= not G11650;
	G2081<=G932 and G928;
	G2091<=G976 and G971;
	G2132<=G1872 and G1882;
	G2160<=G745 and G746;
	G2161<=I5084 and I5085;
	G2264<=G1771 and G1766;
	G2276<=G1765 and G1610;
	G2306<=G1223 and G1218;
	G2379<=G744 and G743;
	G2496<=G374 and G369;
	G2511<=G461 and G456;
	G2525<=G762 and G758;
	G2531<=G658 and G668;
	G2534<=G798 and G794;
	G2544<=G1341 and G1336;
	G2561<=G742 and G741;
	G2563<=I5689 and I5690;
	G2756<=G936 and G2081;
	G2760<=G981 and G2091;
	G2794<=I5886 and I5887;
	G2800<=G2399 and G2369 and G591;
	G2804<=G2132 and G1891;
	G2892<=G1980 and G1976;
	G2895<=G2411 and G1678;
	G2910<=G2424 and G1660;
	G2911<=G2411 and G1675;
	G2917<=G2424 and G1657;
	G2918<=G2411 and G1672;
	G2939<=G2411 and G1687;
	G2940<=G2424 and G1654;
	G2944<=G2424 and G1669;
	G2945<=G2411 and G1684;
	G2950<=G2424 and G1666;
	G2951<=G2411 and G1681;
	G2957<=G2424 and G1663;
	G2981<=G1776 and G2264;
	G2990<=G2061 and G2557 and G1814;
	G3015<=G2028 and G2191;
	G3047<=G1227 and G2306;
	G3089<=G2054 and G2050;
	G3098<=G2331 and G2198;
	G3101<=I6309 and I6310;
	G3104<=I6316 and I6317;
	G3108<=I6330 and I6331;
	G3111<=I6337 and I6338;
	G3257<=G378 and G2496;
	G3263<=G2503 and G2328;
	G3268<=G466 and G2511;
	G3275<=G115 and G2356;
	G3281<=G766 and G2525;
	G3284<=G2531 and G677;
	G3287<=G802 and G2534;
	G3301<=G1346 and G2544;
	G3374<=G1231 and G3047;
	G3381<=G940 and G2756;
	G3383<=G186 and G3228;
	G3389<=G207 and G3228;
	G3396<=G213 and G3228;
	G3400<=G115 and G3164;
	G3407<=G2561 and G3012;
	G3412<=G219 and G3228;
	G3418<=G2379 and G3012;
	G3422<=G225 and G3228;
	G3423<=I6630 and I6631;
	G3429<=G231 and G3228;
	G3434<=G237 and G3228;
	G3497<=G2804 and G1900;
	G3506<=G986 and G2760;
	G3512<=G2050 and G2971;
	G3516<=G1209 and G3015;
	G3533<=G1981 and G2892;
	G3536<=G2390 and G3103;
	G3563<=G3275 and G2126;
	G3586<=G3323 and G2191;
	G3661<=G382 and G3257;
	G3684<=G1710 and G3015;
	G3685<=G1781 and G2981;
	G3695<=G1712 and G3015;
	G3696<=G1713 and G3015;
	G3706<=G471 and G3268;
	G3714<=G1690 and G2991;
	G3718<=G192 and G3164;
	G3772<=G2542 and G3089;
	G3804<=G3098 and G2203;
	G3807<=G3003 and G3062;
	G3829<=G2028 and G2728;
	G3863<=G3323 and G2728;
	G3880<=G3186 and G2023;
	G3904<=G2948 and G2779;
	G3908<=G186 and G3164;
	G3912<=G207 and G3164;
	G3939<=G213 and G3164;
	G3942<=G219 and G3164;
	G3970<=G225 and G3164;
	G3974<=G231 and G3164;
	G3979<=G237 and G3164;
	G3987<=G243 and G3164;
	G3989<=G248 and G3164;
	G3991<=G1738 and G2774;
	G3998<=G2677 and G2276;
	G3999<=G1741 and G2777;
	G4000<=G1744 and G2778;
	G4006<=G201 and G3228;
	G4007<=G2683 and G2276;
	G4008<=G2689 and G2276;
	G4009<=G1747 and G2789;
	G4047<=G2695 and G2276;
	G4048<=G1750 and G2790;
	G4053<=G2701 and G2276;
	G4054<=G1753 and G2793;
	G4058<=G2707 and G2276;
	G4059<=G1756 and G2796;
	G4063<=G2713 and G2276;
	G4064<=G1759 and G2799;
	G4068<=G2719 and G2276;
	G4069<=G1762 and G2802;
	G4070<=G3263 and G2330;
	G4073<=G3200 and G3222;
	G4079<=G2765 and G2276;
	G4097<=G2677 and G2989;
	G4099<=G770 and G3281;
	G4103<=G2683 and G2997;
	G4106<=G3284 and G686;
	G4109<=G806 and G3287;
	G4114<=G1351 and G3301;
	G4115<=G2689 and G3009;
	G4123<=G2695 and G3037;
	G4126<=G2701 and G3040;
	G4128<=G1976 and G2779;
	G4141<=G2707 and G3051;
	G4157<=G2713 and G3055;
	G4161<=G2719 and G3060;
	G4162<=G3106 and G2971;
	G4169<=G2765 and G3066;
	G4220<=G105 and G3539;
	G4223<=G1003 and G3914;
	G4224<=G1092 and G3638;
	G4229<=G999 and G3914;
	G4230<=G1095 and G3638;
	G4235<=G1011 and G3914;
	G4236<=G1098 and G3638;
	G4252<=G1007 and G3914;
	G4253<=G1074 and G3638;
	G4261<=G1019 and G3914;
	G4269<=G1015 and G3914;
	G4316<=G1965 and G3400;
	G4325<=G1166 and G3682;
	G4330<=G1163 and G3693;
	G4334<=G1160 and G3703;
	G4338<=G1157 and G3707;
	G4340<=G1153 and G3715;
	G4341<=G339 and G3586;
	G4342<=G1149 and G3719;
	G4343<=G345 and G3586;
	G4345<=G1169 and G3730;
	G4348<=G3497 and G1909;
	G4358<=G1209 and G3747;
	G4360<=G1861 and G3748;
	G4364<=G1215 and G3756;
	G4383<=G2517 and G3829;
	G4389<=G3529 and G3092;
	G4392<=G3273 and G3829;
	G4397<=G3475 and G2181;
	G4400<=G4088 and G3829;
	G4401<=G2971 and G3772;
	G4421<=G4112 and G2980;
	G4431<=G2268 and G3533;
	G4432<=G3723 and G1975;
	G4465<=G1117 and G3828;
	G4471<=G1121 and G3862;
	G4473<=G1125 and G3874;
	G4477<=G1129 and G3878;
	G4480<=G1133 and G3905;
	G4481<=G1713 and G3906;
	G4483<=G336 and G3586;
	G4484<=G1137 and G3909;
	G4486<=G1711 and G3910;
	G4487<=G1718 and G3911;
	G4489<=G348 and G3586;
	G4490<=G1141 and G3913;
	G4492<=G1786 and G3685;
	G4497<=G351 and G3586;
	G4498<=G1145 and G3940;
	G4500<=G1357 and G3941;
	G4502<=G2031 and G3938;
	G4503<=G654 and G3943;
	G4505<=G354 and G3586;
	G4506<=G1113 and G3944;
	G4512<=G357 and G3586;
	G4518<=G452 and G3975;
	G4522<=G360 and G3586;
	G4529<=G448 and G3980;
	G4534<=G363 and G3586;
	G4537<=G444 and G3988;
	G4542<=G366 and G3586;
	G4548<=G440 and G3990;
	G4550<=G342 and G3586;
	G4553<=G435 and G3995;
	G4554<=G542 and G3996;
	G4559<=G2034 and G3829;
	G4560<=G431 and G4002;
	G4561<=G538 and G4003;
	G4565<=G534 and G4010;
	G4576<=G530 and G4049;
	G4581<=G3766 and G3254;
	G4582<=G525 and G4055;
	G4584<=G3710 and G2322;
	G4585<=G521 and G4060;
	G4604<=G3056 and G3753 and G2325;
	G4610<=G3804 and G2212;
	G4617<=G3275 and G3879;
	G4670<=G192 and G3946;
	G4712<=G1071 and G3638;
	G4714<=G646 and G3333;
	G4715<=G1077 and G3638;
	G4718<=G650 and G3343;
	G4720<=G1023 and G3914;
	G4722<=G426 and G3353;
	G4723<=G3626 and G2779;
	G4725<=G1032 and G3914;
	G4727<=G386 and G3364;
	G4732<=G391 and G3372;
	G4736<=G396 and G3379;
	G4752<=G401 and G3385;
	G4753<=G481 and G3386;
	G4759<=G406 and G3392;
	G4760<=G486 and G3393;
	G4764<=G411 and G3404;
	G4765<=G491 and G3405;
	G4770<=G416 and G3415;
	G4771<=G496 and G3416;
	G4778<=G421 and G3426;
	G4779<=G501 and G3427;
	G4784<=G506 and G3432;
	G4788<=G511 and G3436;
	G4801<=G516 and G3439;
	G4804<=G476 and G3458;
	G4806<=G3215 and G3992 and G2493;
	G4807<=G3015 and G1289 and G3937;
	G4816<=G4070 and G2336;
	G4820<=G186 and G3946;
	G4823<=G207 and G3946;
	G4824<=G774 and G4099;
	G4827<=G213 and G3946;
	G4828<=G4106 and G695;
	G4831<=G810 and G4109;
	G4834<=G219 and G3946;
	G4836<=G643 and G3520;
	G4837<=G1068 and G3638;
	G4838<=G3275 and G4122;
	G4839<=G225 and G3946;
	G4865<=G1080 and G3638;
	G4866<=G231 and G3946;
	G4868<=G1027 and G3914;
	G4869<=G1083 and G3638;
	G4870<=G237 and G3946;
	G4871<=G1864 and G3523;
	G4875<=G995 and G3914;
	G4876<=G1086 and G3638;
	G4877<=G243 and G3946;
	G4878<=G1868 and G3531;
	G4881<=G991 and G3914;
	G4882<=G1089 and G3638;
	G4883<=G248 and G3946;
	G4884<=G3813 and G2971;
	G4890<=G630 and G4739;
	G4891<=G631 and G4739;
	G4892<=G632 and G4739;
	G4893<=G635 and G4739;
	G4902<=G1848 and G4243;
	G4903<=G1849 and G4243;
	G4904<=G1850 and G4243;
	G4905<=G1853 and G4243;
	G4914<=G1062 and G4436;
	G4921<=G2779 and G4431;
	G4932<=G1065 and G4442;
	G4940<=G3500 and G4440;
	G4941<=G1038 and G4451;
	G4949<=G3505 and G4449;
	G4950<=G1415 and G4682;
	G4952<=G1648 and G4457;
	G4959<=G1520 and G4682;
	G4960<=G1403 and G4682;
	G4962<=G1651 and G4461;
	G4967<=G1515 and G4682;
	G4968<=G1432 and G4682;
	G4969<=G1642 and G4463;
	G4971<=G1419 and G4682;
	G4972<=G1436 and G4682;
	G4973<=G1645 and G4467;
	G4977<=G4567 and G4807;
	G4986<=G1411 and G4682;
	G4987<=G1440 and G4682;
	G4989<=G1424 and G4682;
	G4990<=G1444 and G4682;
	G4991<=G1508 and G4640;
	G4992<=G1407 and G4682;
	G4993<=G1448 and G4682;
	G4994<=G1504 and G4640;
	G4995<=G1474 and G4640;
	G4996<=G1428 and G4682;
	G4998<=G1304 and G4485;
	G4999<=G1499 and G4640;
	G5000<=G1470 and G4640;
	G5001<=G1300 and G4491;
	G5002<=G1494 and G4640;
	G5003<=G1466 and G4640;
	G5004<=G1296 and G4499;
	G5005<=G1490 and G4640;
	G5006<=G1462 and G4640;
	G5008<=G1292 and G4507;
	G5009<=G1486 and G4640;
	G5010<=G1458 and G4640;
	G5023<=G1071 and G4511;
	G5024<=G1284 and G4513;
	G5025<=G1482 and G4640;
	G5026<=G1453 and G4640;
	G5029<=G1077 and G4521;
	G5030<=G1280 and G4523;
	G5031<=G1478 and G4640;
	G5041<=G3983 and G4401;
	G5044<=G4348 and G1918;
	G5051<=G4432 and G2834;
	G5067<=G305 and G4811;
	G5074<=G1771 and G4587;
	G5083<=G3709 and G4586;
	G5084<=G1776 and G4591;
	G5090<=G1781 and G4592;
	G5097<=G1786 and G4603;
	G5099<=G4821 and G3829;
	G5100<=G1791 and G4606;
	G5104<=G1796 and G4608;
	G5108<=G1801 and G4614;
	G5110<=G1806 and G4618;
	G5115<=G1394 and G4572;
	G5123<=G1618 and G4669;
	G5126<=G3076 and G4638;
	G5128<=G4474 and G2733;
	G5145<=G1639 and G4673;
	G5148<=G3088 and G4671;
	G5150<=G1275 and G4678;
	G5151<=G4478 and G2733;
	G5168<=G1512 and G4679;
	G5170<=G1811 and G4680;
	G5172<=G4555 and G4549;
	G5173<=G3094 and G4676;
	G5174<=G1235 and G4681;
	G5178<=G2047 and G4401 and G4104;
	G5180<=G4541 and G4533;
	G5181<=G4520 and G4510;
	G5182<=G1240 and G4713;
	G5188<=G4504 and G4496;
	G5190<=G1245 and G4716;
	G5194<=G1610 and G4717;
	G5199<=G1068 and G4719;
	G5201<=G1250 and G4721;
	G5204<=G4838 and G2126;
	G5211<=G1080 and G4724;
	G5212<=G1255 and G4726;
	G5215<=G4276 and G3400;
	G5220<=G1083 and G4729;
	G5221<=G1260 and G4730;
	G5228<=G1086 and G4734;
	G5230<=G1265 and G4735;
	G5233<=G1791 and G4492;
	G5248<=G673 and G4738;
	G5249<=G1089 and G4747;
	G5250<=G1270 and G4748;
	G5254<=G4335 and G4165;
	G5255<=G682 and G4754;
	G5256<=G4297 and G2779;
	G5257<=G691 and G4755;
	G5258<=G700 and G4756;
	G5259<=G627 and G4739;
	G5260<=G1092 and G4758;
	G5263<=G709 and G4761;
	G5264<=G1095 and G4763;
	G5266<=G718 and G4766;
	G5268<=G1098 and G4769;
	G5271<=G727 and G4772;
	G5273<=G1074 and G4776;
	G5276<=G736 and G4780;
	G5279<=G1766 and G4783;
	G5280<=G4593 and G3052;
	G5287<=G3876 and G4782;
	G5318<=G4401 and G1857;
	G5349<=G2126 and G4617;
	G5354<=G2733 and G4460;
	G5390<=G3220 and G4819;
	G5398<=G4610 and G2224;
	G5418<=G1512 and G4344;
	G5421<=G4631 and G2733 and G3819;
	G5444<=G1041 and G4880;
	G5445<=G4631 and G3875 and G2733;
	G5470<=G1044 and G4222;
	G5473<=G4268 and G3518;
	G5476<=G1615 and G4237;
	G5477<=G1887 and G4241;
	G5478<=G1905 and G4242;
	G5479<=G1845 and G4243;
	G5480<=G4279 and G3519;
	G5483<=G1621 and G4254;
	G5484<=G1896 and G4256;
	G5485<=G1914 and G4257;
	G5489<=G4287 and G3521;
	G5491<=G1624 and G4262;
	G5492<=G1654 and G4263;
	G5493<=G1923 and G4265;
	G5497<=G4296 and G3522;
	G5499<=G1627 and G4270;
	G5500<=G1657 and G4272;
	G5501<=G1672 and G4273;
	G5502<=G1932 and G4275;
	G5507<=G4310 and G3528;
	G5510<=G1630 and G4280;
	G5512<=G1660 and G4281;
	G5513<=G1675 and G4282;
	G5514<=G1941 and G4284;
	G5518<=G4317 and G3532;
	G5522<=G1633 and G4289;
	G5523<=G1663 and G4290;
	G5524<=G1678 and G4291;
	G5525<=G1721 and G4292;
	G5526<=G1950 and G4294;
	G5528<=G4322 and G3537;
	G5529<=G4129 and G4288;
	G5530<=G1636 and G4305;
	G5531<=G1666 and G4306;
	G5532<=G1681 and G4307;
	G5533<=G1724 and G4308;
	G5535<=G4327 and G3544;
	G5536<=G4867 and G4298;
	G5537<=G4143 and G4299;
	G5538<=G1669 and G4313;
	G5539<=G1684 and G4314;
	G5540<=G1727 and G4315;
	G5541<=G4331 and G3582;
	G5543<=G4874 and G4312;
	G5544<=G1687 and G4320;
	G5545<=G1730 and G4321;
	G5547<=G1733 and G4326;
	G5569<=G4816 and G2338;
	G5575<=G1618 and G4501;
	G5588<=G1639 and G4508;
	G5591<=G1615 and G4514;
	G5595<=G1621 and G4524;
	G5598<=G778 and G4824;
	G5601<=G1035 and G4375;
	G5602<=G1624 and G4535;
	G5605<=G4828 and G704;
	G5608<=G814 and G4831;
	G5611<=G1047 and G4382;
	G5612<=G1627 and G4543;
	G5617<=G1050 and G4391;
	G5618<=G1630 and G4551;
	G5625<=G1053 and G4399;
	G5626<=G1633 and G4557;
	G5631<=G1056 and G4416;
	G5632<=G1636 and G4563;
	G5640<=G1059 and G4427;
	G5674<=G148 and G5361;
	G5675<=G131 and G5361;
	G5680<=G153 and G5361;
	G5681<=G135 and G5361;
	G5686<=G158 and G5361;
	G5687<=G139 and G5361;
	G5690<=G1567 and G5112;
	G5694<=G162 and G5361;
	G5695<=G166 and G5361;
	G5698<=G1571 and G5116;
	G5699<=G1592 and G5117;
	G5703<=G174 and G5361;
	G5704<=G143 and G5361;
	G5706<=G1574 and G5121;
	G5707<=G1595 and G5122;
	G5720<=G170 and G5361;
	G5721<=G1577 and G5143;
	G5722<=G1598 and G5144;
	G5725<=G1580 and G5166;
	G5726<=G1601 and G5167;
	G5731<=G1583 and G5175;
	G5732<=G1604 and G5176;
	G5737<=G1524 and G5183;
	G5738<=G1586 and G5184;
	G5739<=G1607 and G5185;
	G5744<=G1528 and G5191;
	G5745<=G1549 and G5192;
	G5746<=G1589 and G5193;
	G5755<=G5103 and G5354;
	G5756<=G1531 and G5202;
	G5757<=G1552 and G5203;
	G5769<=G2112 and G4921 and G3818;
	G5770<=G4466 and G5128;
	G5771<=G1534 and G5213;
	G5772<=G1555 and G5214;
	G5781<=G1537 and G5222;
	G5782<=G1558 and G5223;
	G5788<=G1540 and G5231;
	G5789<=G1561 and G5232;
	G5795<=G1543 and G5251;
	G5796<=G1564 and G5252;
	G5804<=G1546 and G5261;
	G5825<=G3204 and G5318;
	G5848<=G3860 and G5519;
	G5853<=G5044 and G1927;
	G5863<=G5272 and G2173;
	G5877<=G4921 and G639;
	G5882<=G5592 and G3829;
	G5897<=G2204 and G5354;
	G5902<=G2555 and G4977;
	G5911<=G3322 and G4977;
	G5913<=G1041 and G5320;
	G5915<=G4168 and G4977;
	G5917<=G1044 and G5320;
	G5918<=G2965 and G5292 and G4609;
	G5919<=G5216 and G2965;
	G5934<=G5215 and G1965;
	G5944<=G1796 and G5233;
	G6047<=G2017 and G4977;
	G6058<=G1035 and G5320;
	G6064<=G5398 and G2230;
	G6067<=G1047 and G5320;
	G6070<=G1050 and G5320;
	G6075<=G549 and G5613;
	G6079<=G1053 and G5320;
	G6083<=G552 and G5619;
	G6087<=G1056 and G5320;
	G6090<=G553 and G5627;
	G6092<=G1059 and G5320;
	G6095<=G1062 and G5320;
	G6098<=G1065 and G5320;
	G6102<=G1038 and G5320;
	G6123<=G5630 and G4311;
	G6126<=G5639 and G4319;
	G6162<=G3584 and G5200;
	G6163<=G4572 and G5354;
	G6179<=G5115 and G5354;
	G6180<=G2190 and G5128;
	G6186<=G546 and G5042;
	G6187<=G5569 and G2340;
	G6193<=G2206 and G5151;
	G6194<=G554 and G5043;
	G6198<=G1499 and G5128;
	G6199<=G557 and G5062;
	G6204<=G3738 and G4921;
	G6205<=G1515 and G5151;
	G6206<=G560 and G5068;
	G6215<=G1504 and G5128;
	G6216<=G2232 and G5151;
	G6217<=G563 and G5073;
	G6221<=G782 and G5598;
	G6224<=G1520 and G5151;
	G6225<=G566 and G5082;
	G6228<=G5605 and G713;
	G6231<=G818 and G5608;
	G6234<=G2244 and G5151;
	G6235<=G569 and G5089;
	G6238<=G572 and G5096;
	G6240<=G182 and G5361;
	G6244<=G2255 and G5151;
	G6245<=G575 and G5098;
	G6246<=G178 and G5361;
	G6247<=G127 and G5361;
	G6316<=G1270 and G5949;
	G6317<=G1304 and G5949;
	G6318<=G1300 and G5949;
	G6319<=G1296 and G5949;
	G6320<=G1292 and G5949;
	G6321<=G1284 and G5949;
	G6322<=G1275 and G5949;
	G6323<=G1235 and G5949;
	G6324<=G1240 and G5949;
	G6325<=G1245 and G5949;
	G6326<=G1250 and G5949;
	G6327<=G1255 and G5949;
	G6328<=G1260 and G5949;
	G6329<=G1265 and G5949;
	G6331<=G201 and G5904;
	G6332<=G1374 and G5904;
	G6333<=G197 and G5904;
	G6334<=G1389 and G5904;
	G6341<=G272 and G5885;
	G6342<=G293 and G5886;
	G6345<=G5823 and G4426;
	G6346<=G5038 and G5883;
	G6347<=G275 and G5890;
	G6348<=G296 and G5891;
	G6350<=G5837 and G4435;
	G6351<=G6210 and G5052;
	G6352<=G278 and G5894;
	G6353<=G299 and G5895;
	G6358<=G5841 and G4441;
	G6359<=G281 and G5898;
	G6360<=G302 and G5899;
	G6362<=G5846 and G4450;
	G6363<=G284 and G5901;
	G6364<=G5851 and G4454;
	G6404<=G2132 and G5748;
	G6410<=G2804 and G5759;
	G6416<=G3497 and G5774;
	G6423<=G4348 and G5784;
	G6430<=G5044 and G5791;
	G6438<=G5853 and G5797;
	G6439<=G4479 and G5919;
	G6463<=G5052 and G6210;
	G6471<=G5224 and G6014;
	G6472<=G5853 and G1936;
	G6502<=G5981 and G3095;
	G6508<=G5983 and G3096;
	G6516<=G5993 and G3097;
	G6525<=G5995 and G3102;
	G6526<=G76 and G6052;
	G6530<=G6207 and G3829;
	G6531<=G79 and G6056;
	G6532<=G339 and G6057;
	G6535<=G345 and G6063;
	G6540<=G1223 and G6072;
	G6544<=G1227 and G6081;
	G6549<=G5515 and G6175;
	G6550<=G1231 and G6089;
	G6554<=G5075 and G6183;
	G6576<=G5762 and G5503;
	G6580<=G1801 and G5944;
	G6616<=G6105 and G3246;
	G6618<=G658 and G6016;
	G6619<=G49 and G6156;
	G6621<=G52 and G6164;
	G6622<=G336 and G6165;
	G6623<=G55 and G6170;
	G6624<=G348 and G6171;
	G6625<=G1218 and G6178;
	G6627<=G58 and G6181;
	G6628<=G351 and G6182;
	G6632<=G61 and G6190;
	G6633<=G354 and G6191;
	G6638<=G64 and G6195;
	G6639<=G357 and G6196;
	G6640<=G5281 and G5801;
	G6645<=G67 and G6202;
	G6646<=G360 and G6203;
	G6647<=G5288 and G5808;
	G6653<=G70 and G6213;
	G6654<=G363 and G6214;
	G6655<=G5296 and G5812;
	G6656<=G2733 and G6061 and G4631;
	G6661<=G73 and G6219;
	G6662<=G366 and G6220;
	G6663<=G6064 and G2237;
	G6666<=G5301 and G5818;
	G6671<=G342 and G6227;
	G6673<=G5305 and G5822;
	G6679<=G4631 and G6074 and G2733;
	G6684<=G5314 and G5836;
	G6687<=G5486 and G5840;
	G6693<=G5494 and G5845;
	G6696<=G5504 and G5850;
	G6699<=G6177 and G4221;
	G6701<=G6185 and G4228;
	G6728<=G6250 and G4318;
	G6730<=G1872 and G6128;
	G6733<=G5678 and G4324;
	G6738<=G2531 and G6137;
	G6741<=G3284 and G6141;
	G6743<=G4106 and G6146;
	G6744<=G4828 and G6151;
	G6745<=G5605 and G6158;
	G6746<=G6228 and G6166;
	G6747<=G2214 and G5897;
	G6752<=G6187 and G2343;
	G6756<=G3010 and G5877;
	G6757<=G2221 and G5919;
	G6759<=G148 and G5919;
	G6760<=G786 and G6221;
	G6763<=G5802 and G4381;
	G6771<=G263 and G5866;
	G6772<=G6228 and G722;
	G6775<=G822 and G6231;
	G6776<=G5809 and G4390;
	G6786<=G178 and G5919;
	G6787<=G266 and G5875;
	G6788<=G287 and G5876;
	G6790<=G5813 and G4398;
	G6791<=G269 and G5880;
	G6792<=G290 and G5881;
	G6794<=G5819 and G4415;
	G6795<=G5036 and G5878;
	G6819<=G243 and G6596;
	G6820<=G1362 and G6596;
	G6821<=G237 and G6596;
	G6822<=G231 and G6596;
	G6823<=G1368 and G6596;
	G6824<=G1371 and G6596;
	G6826<=G225 and G6596;
	G6827<=G219 and G6596;
	G6828<=G1377 and G6596;
	G6829<=G213 and G6596;
	G6830<=G1380 and G6596;
	G6831<=G207 and G6596;
	G6832<=G1383 and G6596;
	G6833<=G186 and G6596;
	G6834<=G1365 and G6596;
	G6838<=G192 and G6596;
	G6839<=G1397 and G6596;
	G6840<=G248 and G6596;
	G6841<=G1400 and G6596;
	G6855<=G1964 and G6392;
	G6872<=G1896 and G6389;
	G6873<=G3263 and G6557;
	G6875<=G1905 and G6400;
	G6876<=G4070 and G6560;
	G6879<=G1914 and G6407;
	G6880<=G4816 and G6562;
	G6883<=G1923 and G6413;
	G6884<=G5569 and G6564;
	G6886<=G1932 and G6420;
	G6887<=G6187 and G6566;
	G6889<=G1941 and G6427;
	G6890<=G6752 and G6568;
	G6891<=G1950 and G6435;
	G6892<=G6472 and G5805;
	G6940<=G6472 and G1945;
	G6983<=G6592 and G3105;
	G6994<=G6758 and G3829;
	G7032<=G2965 and G6626 and G5292;
	G7046<=G5892 and G6570;
	G7050<=G5896 and G6575;
	G7055<=G5900 and G6579;
	G7059<=G6078 and G6714;
	G7060<=G6739 and G5521;
	G7061<=G790 and G6760;
	G7063<=G5903 and G6582;
	G7068<=G5912 and G6586;
	G7071<=G5916 and G6590;
	G7088<=G2331 and G6737;
	G7125<=G1212 and G6648;
	G7127<=G6663 and G2241;
	G7130<=G6041 and G6697;
	G7131<=G6044 and G6700;
	G7132<=G6048 and G6702;
	G7134<=G5587 and G6354;
	G7135<=G869 and G6355;
	G7136<=G6050 and G6704;
	G7137<=G5590 and G6361;
	G7138<=G6055 and G6707;
	G7139<=G6060 and G6709;
	G7140<=G6069 and G6711;
	G7141<=G6073 and G6716;
	G7145<=G6082 and G6718;
	G7182<=G1878 and G6720;
	G7185<=G1887 and G6724;
	G7186<=G2503 and G6403;
	G7191<=G6343 and G4323;
	G7200<=G3098 and G6418;
	G7202<=G6349 and G4329;
	G7209<=G3804 and G6425;
	G7217<=G4610 and G6432;
	G7224<=G5398 and G6441;
	G7230<=G6064 and G6444;
	G7235<=G6663 and G6447;
	G7241<=G6772 and G6172;
	G7260<=G6752 and G2345;
	G7271<=G5028 and G6499;
	G7277<=G6772 and G731;
	G7368<=G6980 and G3880;
	G7378<=G6990 and G3880;
	G7389<=G7001 and G3880;
	G7409<=G4976 and G632 and G6858;
	G7435<=G7260 and G6572;
	G7444<=G7277 and G5827;
	G7449<=G6868 and G4355;
	G7453<=G7148 and G2809;
	G7459<=G7148 and G2814;
	G7466<=G7148 and G2821;
	G7472<=G7148 and G2829;
	G7496<=G7148 and G2840;
	G7504<=G7148 and G2847;
	G7515<=G7148 and G2855;
	G7526<=G7148 and G2868;
	G7535<=G7148 and G2874;
	G7536<=G7148 and G2877;
	G7541<=G7075 and G3109;
	G7542<=G7148 and G2885;
	G7549<=G7269 and G3829;
	G7581<=G7092 and G5420;
	G7586<=G7096 and G5423;
	G7590<=G7102 and G5425;
	G7613<=G6940 and G5984;
	G7623<=G664 and G7079;
	G7625<=G673 and G7085;
	G7632<=G7184 and G5574;
	G7661<=G7127 and G2251;
	G7674<=G7004 and G3880;
	G7679<=G1950 and G6863;
	G7704<=G682 and G7197;
	G7705<=G6853 and G4328;
	G7707<=G691 and G7206;
	G7709<=G6856 and G4333;
	G7710<=G700 and G7214;
	G7718<=G709 and G7221;
	G7719<=G718 and G7227;
	G7720<=G727 and G7232;
	G7721<=G736 and G7237;
	G7722<=G7127 and G6449;
	G7730<=G7260 and G2347;
	G7732<=G6935 and G3880;
	G7734<=G6944 and G3880;
	G7736<=G6951 and G3880;
	G7739<=G6957 and G3880;
	G7741<=G6961 and G3880;
	G7743<=G6967 and G3880;
	G7818<=G1878 and G7479;
	G7819<=G1887 and G7479;
	G7820<=G1896 and G7479;
	G7821<=G1905 and G7479;
	G7822<=G1914 and G7479;
	G7823<=G1923 and G7479;
	G7824<=G1932 and G7479;
	G7825<=G1941 and G7479;
	G7843<=G7599 and G5919;
	G7876<=G7609 and G3790;
	G7879<=G7610 and G3798;
	G7881<=G7612 and G3810;
	G7884<=G7457 and G7022;
	G7885<=G7614 and G3812;
	G7888<=G7465 and G7025;
	G7889<=G7615 and G3814;
	G7891<=G7471 and G7028;
	G7892<=G7616 and G3815;
	G7893<=G7478 and G7031;
	G7894<=G7617 and G3816;
	G7895<=G7503 and G7036;
	G7898<=G7511 and G7041;
	G7902<=G7661 and G6587;
	G7930<=G7621 and G3110;
	G7931<=G2809 and G7446;
	G7933<=G2814 and G7450;
	G7935<=G2821 and G7454;
	G7937<=G7606 and G4013;
	G7939<=G2829 and G7460;
	G7940<=G7620 and G4013;
	G7943<=G2840 and G7467;
	G7945<=G2847 and G7473;
	G7948<=G2855 and G7497;
	G7951<=G2868 and G7505;
	G7954<=G2874 and G7512;
	G7955<=G2877 and G7516;
	G7957<=G2885 and G7527;
	G7958<=G736 and G7697;
	G7962<=G7730 and G6712;
	G7970<=G7384 and G7703;
	G7988<=G1878 and G7379;
	G8005<=G7510 and G6871;
	G8010<=G7738 and G7413;
	G8014<=G7740 and G7419;
	G8018<=G7742 and G7425;
	G8019<=G7386 and G4332;
	G8023<=G7367 and G7430;
	G8024<=G7394 and G4337;
	G8028<=G7375 and G7436;
	G8032<=G7385 and G7438;
	G8039<=G7587 and G5128;
	G8040<=G7523 and G5128;
	G8041<=G7524 and G5128;
	G8042<=G7533 and G5128;
	G8043<=G7582 and G5128;
	G8044<=G7598 and G5919;
	G8045<=G7547 and G5128;
	G8046<=G7548 and G5128;
	G8047<=G7557 and G5919;
	G8048<=G7558 and G5919;
	G8049<=G7567 and G5919;
	G8050<=G7596 and G5919;
	G8051<=G7572 and G5128;
	G8052<=G7573 and G5128;
	G8053<=G7583 and G5919;
	G8054<=G7584 and G5919;
	G8055<=G7588 and G5128;
	G8059<=G7592 and G5919;
	G8060<=G7593 and G5919;
	G8068<=G664 and G7826;
	G8069<=G673 and G7826;
	G8070<=G682 and G7826;
	G8071<=G691 and G7826;
	G8072<=G700 and G7826;
	G8073<=G709 and G7826;
	G8074<=G718 and G7826;
	G8075<=G727 and G7826;
	G8097<=G6200 and G7851;
	G8098<=G6201 and G7852;
	G8101<=G6208 and G7877;
	G8102<=G6209 and G7878;
	G8104<=G6218 and G7880;
	G8107<=G6226 and G7882;
	G8108<=G1891 and G7938;
	G8117<=G6236 and G7886;
	G8118<=G1900 and G7941;
	G8119<=G6239 and G7890;
	G8120<=G1909 and G7944;
	G8123<=G1918 and G7946;
	G8127<=G1927 and G7949;
	G8130<=G1936 and G7952;
	G8135<=G1945 and G7956;
	G8136<=G7926 and G7045;
	G8147<=G2955 and G7961;
	G8163<=G7960 and G3737;
	G8167<=G5253 and G7853;
	G8168<=G5262 and G7853;
	G8169<=G5265 and G7853;
	G8170<=G5270 and G7853;
	G8172<=G5275 and G7853;
	G8173<=G7971 and G3112;
	G8174<=G5284 and G7853;
	G8175<=G5291 and G7853;
	G8176<=G5299 and G7853;
	G8185<=G664 and G7997;
	G8209<=G4094 and G3792 and G7980;
	G8217<=G1872 and G7883;
	G8224<=G1882 and G7887;
	G8244<=G7847 and G4336;
	G8245<=G7850 and G4339;
	G8246<=G7846 and G7442;
	G8250<=G2771 and G7907;
	G8254<=G2773 and G7909;
	G8260<=G2775 and G7911;
	G8289<=G6777 and G8109 and G6475;
	G8364<=G658 and G8235;
	G8365<=G668 and G8240;
	G8366<=G8199 and G7265;
	G8380<=G8252 and G4240;
	G8382<=G6077 and G8213;
	G8384<=G8180 and G3397;
	G8385<=G6084 and G8218;
	G8386<=G6085 and G8219;
	G8387<=G6086 and G8220;
	G8388<=G8177 and G7689;
	G8389<=G6091 and G8225;
	G8390<=G8268 and G6465;
	G8399<=G6094 and G8229;
	G8400<=G6097 and G8234;
	G8401<=G677 and G8124;
	G8403<=G6101 and G8239;
	G8404<=G686 and G8129;
	G8406<=G695 and G8131;
	G8408<=G704 and G8139;
	G8410<=G713 and G8143;
	G8413<=G722 and G8146;
	G8416<=G731 and G8151;
	G8461<=G8298 and G7403;
	G8462<=G8300 and G7406;
	G8463<=G8301 and G7410;
	G8464<=G8302 and G7416;
	G8469<=G8305 and G7422;
	G8470<=G8308 and G7427;
	G8474<=G8383 and G5285;
	G8499<=G8377 and G4737;
	G8505<=G8309 and G4789;
	G8508<=G8411 and G7967;
	G8510<=G8414 and G7972;
	G8547<=G8307 and G7693;
	G8550<=G8402 and G8011;
	G8553<=G8405 and G8015;
	G8554<=G8407 and G8020;
	G8555<=G8409 and G8025;
	G8556<=G8412 and G8029;
	G8557<=G8415 and G8033;
	G8598<=G8471 and G7432;
	G8603<=G3983 and G8548;
	G8648<=G4588 and G8511;
	G8651<=G8520 and G4013;
	G8652<=G8523 and G4013;
	G8653<=G8526 and G4013;
	G8654<=G8529 and G4013;
	G8655<=G8532 and G4013;
	G8659<=G8535 and G4013;
	G8663<=G8538 and G4013;
	G8683<=G4803 and G8549;
	G8687<=G8558 and G8036;
	G8693<=G3738 and G8509;
	G8698<=G7591 and G8576;
	G8699<=G7595 and G8579;
	G8701<=G7597 and G8582;
	G8703<=G7601 and G8585;
	G8706<=G7602 and G8589;
	G8708<=G7605 and G8592;
	G8710<=G7607 and G8595;
	G8718<=G8600 and G7903;
	G8720<=G8601 and G7905;
	G8722<=G8604 and G7908;
	G8724<=G8606 and G7910;
	G8726<=G8608 and G7913;
	G8728<=G8610 and G7915;
	G8730<=G8613 and G7917;
	G8731<=G8622 and G7918;
	G8732<=G8624 and G7919;
	G8733<=G8625 and G7920;
	G8734<=G8626 and G7923;
	G8735<=G7600 and G8632;
	G8736<=G7439 and G8635;
	G8748<=G7670 and G8656;
	G8749<=G7604 and G8660;
	G8753<=G7414 and G8664;
	G8754<=G7420 and G8667;
	G8755<=G7426 and G8671;
	G8756<=G7431 and G8674;
	G8759<=G7437 and G8677;
	G8763<=G7440 and G8680;
	G8764<=G7443 and G8684;
	G8765<=G8630 and G5151;
	G8766<=G8612 and G5151;
	G8767<=G8616 and G5151;
	G8768<=G8623 and G5151;
	G8769<=G8629 and G5151;
	G8772<=G8627 and G5151;
	G8775<=G8628 and G5151;
	G8778<=G8688 and G2317;
	G8786<=G8638 and G8716;
	G8789<=G8639 and G8719;
	G8791<=G8641 and G8721;
	G8793<=G8644 and G8723;
	G8796<=G8645 and G8725;
	G8799<=G8647 and G8727;
	G8801<=G8742 and G8729;
	G8820<=G8705 and G5422;
	G8821<=G8643 and G8751;
	G8822<=G8614 and G8752;
	G8827<=G8552 and G8696;
	G8837<=G8646 and G8697;
	G8838<=G8602 and G8702;
	G8841<=G8605 and G8704;
	G8842<=G8607 and G8707;
	G8844<=G8609 and G8709;
	G8845<=G8611 and G8711;
	G8846<=G8615 and G8712;
	G8848<=G8715 and G8713;
	G8875<=G8255 and G6368 and G8858;
	G8876<=G8105 and G6764 and G8858;
	G8877<=G8103 and G6764 and G8858;
	G8878<=G8099 and G6368 and G8858;
	G8879<=G8110 and G6764 and G8858;
	G8927<=G7872 and G8807;
	G8929<=G8095 and G6368 and G8828;
	G8930<=G8100 and G6368 and G8828;
	G8931<=G8807 and G8164;
	G8935<=G8106 and G6778 and G8849;
	G8936<=G8115 and G6778 and G8849;
	G8947<=G8056 and G6368 and G8828;
	G8949<=G8255 and G6368 and G8828;
	G8955<=G8110 and G6368 and G8828;
	G8957<=G8081 and G6368 and G8828;
	G8960<=G8085 and G6368 and G8828;
	G8962<=G8089 and G6368 and G8828;
	G8963<=G8056 and G6368 and G8849;
	G8964<=G8255 and G6368 and G8849;
	G8965<=G8110 and G6778 and G8849;
	G8966<=G8081 and G6778 and G8849;
	G8967<=G8085 and G6778 and G8849;
	G8968<=G8089 and G6778 and G8849;
	G8971<=G8081 and G6764 and G8858;
	G8972<=G8085 and G6764 and G8858;
	G8974<=G8094 and G6368 and G8858;
	G8975<=G8089 and G6764 and G8858;
	G8994<=G8110 and G6778 and G8925;
	G8995<=G6454 and G8929;
	G9010<=G6454 and G8930;
	G9030<=G8935 and G7192;
	G9052<=G8936 and G7192;
	G9110<=G8880 and G4790;
	G9111<=G8965 and G6674;
	G9124<=G8881 and G4802;
	G9125<=G8966 and G6674;
	G9150<=G8882 and G4805;
	G9151<=G8967 and G6674;
	G9173<=G8968 and G6674;
	G9192<=G6454 and G8955;
	G9205<=G6454 and G8957;
	G9223<=G6454 and G8960;
	G9240<=G6454 and G8962;
	G9256<=G6689 and G8963;
	G9257<=G6689 and G8964;
	G9266<=G8932 and G3398;
	G9268<=G6681 and G8947;
	G9269<=G8933 and G3413;
	G9271<=G6681 and G8949;
	G9272<=G8934 and G3424;
	G9274<=G8974 and G5708;
	G9292<=G8878 and G5708;
	G9313<=G8876 and G5708;
	G9316<=G8877 and G5708;
	G9317<=G6109 and G8875;
	G9324<=G8879 and G5708;
	G9328<=G8971 and G5708;
	G9331<=G8972 and G5708;
	G9335<=G8975 and G5708;
	G9357<=G962 and G9223;
	G9358<=G1318 and G9151;
	G9359<=G1308 and G9173;
	G9364<=G965 and G9223;
	G9365<=G1321 and G9151;
	G9366<=G1311 and G9173;
	G9384<=G968 and G9223;
	G9385<=G1324 and G9151;
	G9386<=G1327 and G9151;
	G9389<=G1330 and G9151;
	G9390<=G1333 and G9151;
	G9409<=G1721 and G9052;
	G9411<=G1724 and G9052;
	G9412<=G1727 and G9052;
	G9414<=G1730 and G9052;
	G9415<=G1733 and G9052;
	G9417<=G1738 and G9052;
	G9418<=G1741 and G9052;
	G9419<=G1744 and G9030;
	G9420<=G1747 and G9030;
	G9422<=G1750 and G9030;
	G9425<=G1753 and G9030;
	G9428<=G1756 and G9030;
	G9430<=G1759 and G9030;
	G9447<=G1762 and G9030;
	G9454<=G8994 and G5708;
	G9555<=G9107 and G3391;
	G9582<=G2725 and G9173;
	G9583<=G886 and G8995;
	G9584<=G2726 and G9173;
	G9585<=G889 and G8995;
	G9586<=G2727 and G9173;
	G9587<=G892 and G8995;
	G9588<=G3272 and G9173;
	G9590<=G895 and G8995;
	G9592<=G4 and G9292;
	G9593<=G898 and G9205;
	G9594<=G1 and G9292;
	G9595<=G901 and G9205;
	G9596<=G2649 and G9010;
	G9597<=G1170 and G9125;
	G9598<=G2086 and G9274;
	G9599<=G8 and G9292;
	G9600<=G904 and G9205;
	G9601<=G922 and G9192;
	G9602<=G2650 and G9010;
	G9603<=G1173 and G9125;
	G9604<=G1194 and G9111;
	G9607<=G12 and G9274;
	G9608<=G7 and G9292;
	G9609<=G907 and G9205;
	G9610<=G925 and G9192;
	G9611<=G2651 and G9010;
	G9612<=G2652 and G9240;
	G9613<=G1176 and G9125;
	G9614<=G1197 and G9111;
	G9617<=G9 and G9274;
	G9618<=G910 and G9205;
	G9619<=G2772 and G9010;
	G9620<=G2653 and G9240;
	G9621<=G1179 and G9125;
	G9622<=G1200 and G9111;
	G9623<=G17 and G9274;
	G9641<=G913 and G9205;
	G9642<=G2654 and G9240;
	G9643<=G950 and G9223;
	G9644<=G1182 and G9125;
	G9645<=G1203 and G9111;
	G9648<=G16 and G9274;
	G9649<=G916 and G9205;
	G9650<=G2797 and G9240;
	G9651<=G944 and G9240;
	G9652<=G953 and G9223;
	G9653<=G1185 and G9125;
	G9657<=G919 and G9205;
	G9658<=G947 and G9240;
	G9659<=G956 and G9223;
	G9660<=G1188 and G9125;
	G9662<=G2094 and G9292;
	G9663<=G959 and G9223;
	G9664<=G1191 and G9125;
	G9665<=G1314 and G9151;
	G9689<=G263 and G9432;
	G9690<=G266 and G9432;
	G9691<=G269 and G9432;
	G9692<=G272 and G9432;
	G9693<=G275 and G9432;
	G9694<=G278 and G9432;
	G9695<=G1567 and G9474;
	G9696<=G281 and G9432;
	G9698<=G1571 and G9474;
	G9699<=G284 and G9432;
	G9701<=G1574 and G9474;
	G9703<=G1577 and G9474;
	G9705<=G1580 and G9474;
	G9707<=G1583 and G9474;
	G9709<=G1524 and G9490;
	G9710<=G1586 and G9474;
	G9712<=G1528 and G9490;
	G9713<=G1589 and G9474;
	G9715<=G1531 and G9490;
	G9716<=G1534 and G9490;
	G9717<=G1537 and G9490;
	G9718<=G1540 and G9490;
	G9719<=G1543 and G9490;
	G9720<=G1546 and G9490;
	G9721<=G9413 and G4785;
	G9828<=G9722 and G9785;
	G9829<=G9723 and G9785;
	G9830<=G9725 and G9785;
	G9831<=G9727 and G9785;
	G9833<=G9729 and G9785;
	G9834<=G9731 and G9785;
	G9835<=G9735 and G9785;
	G9836<=G9737 and G9785;
	G9837<=G9697 and G9751;
	G9838<=G9700 and G9754;
	G9839<=G9702 and G9742;
	G9840<=G9704 and G9747;
	G9841<=G9706 and G9512;
	G9842<=G9708 and G9516;
	G9843<=G9711 and G9519;
	G9844<=G9714 and G9522;
	G9846<=G287 and G9764;
	G9847<=G290 and G9766;
	G9848<=G9724 and G9557;
	G9849<=G293 and G9768;
	G9850<=G9726 and G9560;
	G9851<=G296 and G9770;
	G9852<=G9728 and G9563;
	G9853<=G299 and G9771;
	G9854<=G9730 and G9566;
	G9855<=G302 and G9772;
	G9856<=G1592 and G9773;
	G9857<=G9734 and G9569;
	G9858<=G1595 and G9774;
	G9859<=G9736 and G9573;
	G9860<=G1598 and G9775;
	G9861<=G9738 and G9579;
	G9862<=G1601 and G9777;
	G9863<=G9740 and G9576;
	G9864<=G1604 and G9778;
	G9865<=G1607 and G9780;
	G9866<=G1549 and G9802;
	G9867<=G1552 and G9807;
	G9868<=G1555 and G9812;
	G9869<=G1558 and G9814;
	G9870<=G1561 and G9816;
	G9871<=G1564 and G9668;
	G9896<=G9883 and G9624;
	G9897<=G9884 and G9624;
	G9898<=G9887 and G9367;
	G9899<=G9889 and G9367;
	G9900<=G9845 and G8327;
	G9901<=G9893 and G9392;
	G9902<=G9894 and G9392;
	G9903<=G9885 and G9673;
	G9904<=G9886 and G9676;
	G9905<=G9872 and G9680;
	G9906<=G9873 and G9683;
	G9907<=G9888 and G9686;
	G9908<=G9890 and G9782;
	G9909<=G9891 and G9804;
	G9910<=G9892 and G9809;
	G9932<=G9911 and G9624;
	G9933<=G9912 and G9624;
	G9934<=G9913 and G9624;
	G9935<=G9914 and G9624;
	G9936<=G9915 and G9624;
	G9937<=G9916 and G9624;
	G9938<=G9917 and G9367;
	G9939<=G9918 and G9367;
	G9940<=G9920 and G9367;
	G9941<=G9921 and G9367;
	G9942<=G9922 and G9367;
	G9943<=G9923 and G9367;
	G9944<=G9924 and G9392;
	G9945<=G9925 and G9392;
	G9946<=G9926 and G9392;
	G9947<=G9927 and G9392;
	G9948<=G9928 and G9392;
	G9949<=G9929 and G9392;
	G9959<=G9950 and G9536;
	G9960<=G9951 and G9536;
	G9962<=G9952 and G9536;
	G9963<=G9953 and G9536;
	G9964<=G9954 and G9536;
	G9965<=G9955 and G9536;
	G9966<=G9956 and G9536;
	G9967<=G9957 and G9536;
	G10230<=G8892 and G10145;
	G10232<=G8892 and G10150;
	G10237<=G10145 and G9100;
	G10240<=G10150 and G9103;
	G10268<=G10183 and G3307;
	G10295<=G8892 and G10208;
	G10297<=G8892 and G10211;
	G10298<=G8892 and G10214;
	G10299<=G8892 and G10217;
	G10300<=G8892 and G10220;
	G10301<=G8892 and G10223;
	G10303<=G10208 and G9076;
	G10304<=G10211 and G9079;
	G10306<=G10214 and G9082;
	G10308<=G10217 and G9085;
	G10312<=G10220 and G9094;
	G10316<=G10223 and G9097;
	G10325<=G10248 and G3307;
	G10328<=G10252 and G3307;
	G10331<=G10256 and G3307;
	G10333<=G10262 and G3307;
	G10334<=G10265 and G3307;
	G10348<=G10272 and G3705;
	G10357<=G10278 and G2462;
	G10365<=G10319 and G2135;
	G10367<=G10362 and G3375;
	G10369<=G10361 and G3382;
	G10442<=G10311 and G2135;
	G10445<=G10315 and G2135;
	G10448<=G10421 and G3335;
	G10449<=G10420 and G3345;
	G10450<=G10364 and G3359;
	G10451<=G10444 and G3365;
	G10452<=G10439 and G3388;
	G10453<=G10437 and G3395;
	G10454<=G10435 and G3411;
	G10494<=G10433 and G3945;
	G10495<=G10431 and G3971;
	G10496<=G10429 and G3977;
	G10503<=G10388 and G2135;
	G10504<=G10389 and G2135;
	G10506<=G10390 and G2135;
	G10508<=G10391 and G2135;
	G10510<=G10393 and G2135;
	G10512<=G10395 and G2135;
	G10514<=G10489 and G4580;
	G10515<=G10505 and G10469 and I16142;
	G10518<=G10513 and G10440 and I16145;
	G10560<=G10487 and G4575;
	G10561<=G10549 and G4583;
	G10581<=G10531 and G9453;
	G10582<=G10532 and G9473;
	G10583<=G10518 and G10515;
	G10595<=G10550 and G4347;
	G10597<=G10533 and G4359;
	G10599<=G10534 and G4365;
	G10622<=G10543 and G4525;
	G10623<=G10544 and G4536;
	G10624<=G10545 and G4544;
	G10625<=G10546 and G4552;
	G10626<=G10547 and G4558;
	G10627<=G10548 and G4564;
	G10633<=G10600 and G3829;
	G10634<=G10604 and G3829;
	G10638<=G10608 and G3829;
	G10642<=G10612 and G3829;
	G10661<=G10594 and G3015;
	G10662<=G8892 and G10571;
	G10666<=G10575 and G9424;
	G10667<=G10576 and G9427;
	G10669<=G10577 and G9429;
	G10670<=G10571 and G9091;
	G10671<=G10578 and G9431;
	G10672<=G10579 and G9449;
	G10673<=G10580 and G9450;
	G10680<=G10564 and G3586;
	G10681<=G10567 and G3586;
	G10682<=G10600 and G3863;
	G10684<=G10604 and G3863;
	G10685<=G10608 and G3863;
	G10686<=G10612 and G3863;
	G10690<=G10616 and G3863;
	G10701<=G10620 and G10619;
	G10705<=G10564 and G4840;
	G10706<=G10567 and G4840;
	G10715<=G2272 and G10630;
	G10716<=G10497 and G10675;
	G10731<=G5118 and G1850 and G10665;
	G10736<=G10658 and G4840;
	G10737<=G10687 and G4840;
	G10738<=G10692 and G4840;
	G10739<=G10676 and G3368;
	G10740<=G10676 and G3384;
	G10741<=G10635 and G4013;
	G10742<=G10655 and G3586;
	G10743<=G10639 and G4013;
	G10745<=G10658 and G3586;
	G10746<=G10643 and G4013;
	G10750<=G10687 and G3586;
	G10751<=G10646 and G4013;
	G10752<=G10692 and G3586;
	G10753<=G10649 and G4013;
	G10758<=G10652 and G4013;
	G10759<=G10698 and G10697;
	G10760<=G10695 and G10691;
	G10761<=G10700 and G10699;
	G10762<=G10635 and G4840;
	G10763<=G10639 and G4840;
	G10764<=G10643 and G4840;
	G10766<=G10646 and G4840;
	G10768<=G10649 and G4840;
	G10769<=G10652 and G4840;
	G10772<=G10655 and G4840;
	G10777<=G10733 and G3015;
	G10778<=G1027 and G10729;
	G10780<=G10723 and G5124;
	G10782<=G10725 and G5146;
	G10784<=G10727 and G5169;
	G10785<=G10728 and G5177;
	G10788<=G8303 and G10754;
	G10808<=G10744 and G3829;
	G10809<=G4811 and G10754;
	G10818<=G10730 and G4545;
	G10933<=G10853 and G3982;
	G10937<=G4822 and G10822;
	G10946<=G5225 and G10827;
	G10948<=G2223 and G10809;
	G10949<=G2947 and G10809;
	G10950<=G10788 and G6355;
	G10969<=G3625 and G10809;
	G10970<=G10852 and G3390;
	G10971<=G10849 and G3161;
	G11005<=G5119 and G10827;
	G11006<=G5125 and G10827;
	G11007<=G5147 and G10827;
	G11008<=G5171 and G10827;
	G11009<=G5179 and G10827;
	G11010<=G5187 and G10827;
	G11011<=G1968 and G10809;
	G11012<=G5196 and G10827;
	G11013<=G5209 and G10827;
	G11015<=G5217 and G10827;
	G11018<=G7286 and G10974;
	G11019<=G421 and G10974;
	G11020<=G452 and G10974;
	G11021<=G448 and G10974;
	G11022<=G444 and G10974;
	G11023<=G440 and G10974;
	G11024<=G435 and G10974;
	G11025<=G426 and G10974;
	G11026<=G386 and G10974;
	G11027<=G391 and G10974;
	G11028<=G396 and G10974;
	G11029<=G401 and G10974;
	G11030<=G406 and G10974;
	G11031<=G411 and G10974;
	G11032<=G416 and G10974;
	G11070<=G2008 and G10913;
	G11085<=G312 and G10897;
	G11087<=G829 and G10950;
	G11091<=G833 and G10950;
	G11092<=G837 and G10950;
	G11093<=G841 and G10950;
	G11094<=G374 and G10883;
	G11095<=G845 and G10950;
	G11097<=G378 and G10884;
	G11098<=G849 and G10950;
	G11099<=G382 and G10885;
	G11100<=G853 and G10950;
	G11101<=G857 and G10950;
	G11102<=G861 and G10950;
	G11103<=G2250 and G10937;
	G11104<=G2963 and G10937;
	G11105<=G3634 and G10937;
	G11143<=G10923 and G4567;
	G11144<=G305 and G10926;
	G11145<=G315 and G10927;
	G11146<=G318 and G10928;
	G11147<=G321 and G10929;
	G11148<=G2321 and G10913;
	G11149<=G324 and G10930;
	G11150<=G3087 and G10913;
	G11151<=G327 and G10931;
	G11152<=G369 and G10903;
	G11153<=G3771 and G10913;
	G11154<=G330 and G10932;
	G11156<=G333 and G10934;
	G11158<=G309 and G10935;
	G11161<=G1969 and G10937;
	G11164<=G4889 and G11112;
	G11165<=G476 and G11112;
	G11166<=G542 and G11112;
	G11167<=G538 and G11112;
	G11168<=G534 and G11112;
	G11169<=G530 and G11112;
	G11170<=G525 and G11112;
	G11171<=G481 and G11112;
	G11172<=G486 and G11112;
	G11173<=G491 and G11112;
	G11174<=G496 and G11112;
	G11175<=G501 and G11112;
	G11176<=G506 and G11112;
	G11177<=G511 and G11112;
	G11178<=G516 and G11112;
	G11186<=G5594 and G11059;
	G11187<=G5597 and G11061;
	G11188<=G5604 and G11063;
	G11189<=G5616 and G11064;
	G11190<=G5623 and G11065;
	G11192<=G5628 and G11066;
	G11194<=G5637 and G11067;
	G11196<=G4912 and G11068;
	G11198<=G4919 and G11069;
	G11204<=G971 and G11083;
	G11209<=G11074 and G9448;
	G11210<=G11078 and G4515;
	G11211<=G11058 and G5534;
	G11212<=G944 and G11155;
	G11213<=G947 and G11157;
	G11214<=G950 and G11159;
	G11215<=G953 and G11160;
	G11216<=G956 and G11162;
	G11218<=G959 and G11053;
	G11220<=G962 and G11054;
	G11222<=G965 and G11055;
	G11224<=G968 and G11056;
	G11226<=G461 and G11057;
	G11228<=G466 and G11060;
	G11230<=G471 and G11062;
	G11234<=G5424 and G11106;
	G11235<=G5443 and G11107;
	G11236<=G5469 and G11108;
	G11237<=G5472 and G11109;
	G11238<=G5474 and G11110;
	G11240<=G5481 and G11111;
	G11248<=G976 and G11071;
	G11253<=G981 and G11072;
	G11254<=G986 and G11073;
	G11255<=G456 and G11075;
	G11271<=G5624 and G11191;
	G11272<=G5629 and G11193;
	G11273<=G5638 and G11195;
	G11274<=G4913 and G11197;
	G11277<=G4920 and G11199;
	G11279<=G4939 and G11200;
	G11281<=G4948 and G11202;
	G11282<=G4958 and G11203;
	G11283<=G4966 and G11205;
	G11290<=G11246 and G4226;
	G11291<=G11247 and G4233;
	G11292<=G11252 and G4250;
	G11295<=G5475 and G11239;
	G11296<=G5482 and G11241;
	G11297<=G5490 and G11242;
	G11299<=G5498 and G11243;
	G11302<=G5508 and G11244;
	G11304<=G5520 and G11245;
	G11320<=G11201 and G4379;
	G11340<=G11285 and G4424;
	G11349<=G11288 and G7964;
	G11372<=G11316 and G4266;
	G11376<=G11318 and G4277;
	G11380<=G11321 and G4285;
	G11387<=G11284 and G3629;
	G11391<=G11275 and G7912;
	G11392<=G11278 and G7914;
	G11393<=G11280 and G7916;
	G11407<=G11339 and G5949;
	G11413<=G11354 and G10679;
	G11425<=G11350 and G10899;
	G11455<=G11435 and G5446;
	G11456<=G3765 and G3517 and G11422;
	G11458<=G11426 and G5446;
	G11459<=G11427 and G5446;
	G11460<=G11428 and G5446;
	G11461<=G11429 and G5446;
	G11462<=G11431 and G5446;
	G11463<=G11432 and G5446;
	G11464<=G11433 and G5446;
	G11465<=G11434 and G5446;
	G11492<=G11480 and G4807;
	G11514<=G11491 and G5151;
	G11519<=G1317 and G3015 and G11492;
	G11544<=G11515 and G10584;
	G11551<=G11538 and G4013;
	G11552<=G2677 and G11519;
	G11553<=G2683 and G11519;
	G11554<=G2689 and G11519;
	G11555<=G2695 and G11519;
	G11556<=G2701 and G11519;
	G11557<=G2707 and G11519;
	G11558<=G2713 and G11519;
	G11559<=G2719 and G11519;
	G11560<=G2765 and G11519;
	G11561<=G11518 and G3015;
	G11571<=G2018 and G11561;
	G11581<=G1308 and G11539;
	G11582<=G1311 and G11540;
	G11583<=G1314 and G11541;
	G11584<=G1318 and G11542;
	G11585<=G1321 and G11543;
	G11586<=G1324 and G11545;
	G11587<=G1327 and G11546;
	G11588<=G1330 and G11547;
	G11589<=G1333 and G11548;
	G11590<=G2274 and G11561;
	G11591<=G2988 and G11561;
	G11592<=G3717 and G11561;
	G11595<=G1336 and G11575;
	G11597<=G11576 and G5446;
	G11599<=G1341 and G11572;
	G11600<=G1346 and G11573;
	G11601<=G1351 and G11574;
	G11636<=G11624 and G7936;
	G11637<=G11626 and G5446;
	G11639<=G11612 and G7897;
	G11640<=G11613 and G7900;
	G11641<=G11615 and G7901;
	I5084<=G1462 and G1470 and G1474 and G1478;
	I5085<=G1490 and G1494 and G1504 and G1508;
	I5689<=G1419 and G1424 and G1428 and G1432;
	I5690<=G1436 and G1440 and G1444 and G1448;
	I5886<=G174 and G170 and G2249 and G2254;
	I5887<=G2078 and G2083 and G166 and G2095;
	I6309<=G2446 and G2451 and G2456 and G2475;
	I6310<=G2396 and G2407 and G2421 and G2435;
	I6316<=G2082 and G2087 and G2381 and G2395;
	I6317<=G2406 and G2420 and G2434 and G2438;
	I6330<=G2549 and G2556 and G2562 and G2570;
	I6331<=G2060 and G2070 and G2074 and G2077;
	I6337<=G201 and G2421 and G2407 and G2396;
	I6338<=G2475 and G2456 and G2451 and G2446;
	I6630<=G2677 and G2683 and G2689 and G2701;
	I6631<=G2707 and G2713 and G2719 and G2765;
	I16142<=G10511 and G10509 and G10507;
	I16145<=G10366 and G10447 and G10446;
	G2088<= not (I4911 and I4912);
	G2096<= not (I4929 and I4930);
	G2099<= not (I4942 and I4943);
	G2102<= not (I4955 and I4956);
	G2104<= not (I4965 and I4966);
	G2105<= not (I4972 and I4973);
	G2106<= not (I4979 and I4980);
	G2107<= not (I4986 and I4987);
	G2109<= not (I4996 and I4997);
	G2111<= not (I5006 and I5007);
	G2115<= not (I5014 and I5015);
	G2117<= not (I5024 and I5025);
	G2120<= not (I5035 and I5036);
	G2167<= not (I5105 and I5106);
	G2177<= not (I5127 and I5128);
	G2180<= not (I5136 and I5137);
	G2205<= not (I5165 and I5166);
	G2215<= not (I5185 and I5186);
	G2223<= not (I5203 and I5204);
	G2236<= not (I5230 and I5231);
	G2250<= not (I5264 and I5265);
	G2257<= not (I5283 and I5284);
	G2260<= not (I5296 and I5297);
	G2272<= not (I5316 and I5317);
	G2274<= not (I5324 and I5325);
	G2303<= not (I5342 and I5343);
	G2310<= not (G591 and G605);
	G2321<= not (I5372 and I5373);
	G2325<= not (G611 and G617);
	G2354<= not (G1515 and G1520);
	G2372<= not (I5450 and I5451);
	G2380<= not (I5460 and I5461);
	G2389<= not (I5469 and I5470);
	G2405<= not (I5485 and I5486);
	G2419<= not (I5501 and I5502);
	G2433<= not (I5517 and I5518);
	G2437<= not (I5529 and I5530);
	G2439<= not (G1814 and G1828);
	G2445<= not (I5539 and I5540);
	G2493<= not (G1834 and G1840);
	G2500<= not (G178 and G182);
	G2510<= not (I5592 and I5593);
	G2515<= not (I5605 and I5606);
	G2516<= not (I5612 and I5613);
	G2517<= not (I5619 and I5620);
	G2555<= not (I5676 and I5677);
	G2776<= not (I5866 and I5867);
	G2792<= not (I5879 and I5880);
	G2795<= not (I5892 and I5893);
	G2938<= not (I6110 and I6111);
	G2943<= not (I6125 and I6126);
	G2947<= not (I6137 and I6138);
	G2948<= not (I6144 and I6145);
	G2959<= not (I6167 and I6168);
	G2961<= not (I6177 and I6178);
	G2963<= not (I6187 and I6188);
	G2970<= not (I6200 and I6201);
	G2979<= not (I6208 and I6209);
	G2987<= not (G2481 and G883);
	G2988<= not (I6225 and I6226);
	G3003<= not (G599 and G2399);
	G3008<= not (G2444 and G878);
	G3010<= not (G2382 and G2399);
	G3011<= not (G591 and G2382);
	G3041<= not (G2364 and G2399 and G2374 and G2382);
	G3056<= not (G2374 and G599);
	G3061<= not (G611 and G2374);
	G3062<= not (G2369 and G591 and G611);
	G3070<= not (G2016 and G1206);
	G3071<= not (G605 and G2374 and G2382);
	G3087<= not (I6288 and I6289);
	G3106<= not (I6323 and I6324);
	G3200<= not (G1822 and G2061);
	G3204<= not (G2571 and G2061);
	G3205<= not (G1814 and G2571);
	G3209<= not (G2550 and G2061 and G2564 and G2571);
	G3215<= not (G2564 and G1822);
	G3221<= not (G1834 and G2564);
	G3222<= not (G2557 and G1814 and G1834);
	G3247<= not (G1828 and G2564 and G2571);
	G3261<= not (G2229 and G2222 and G2211 and G2202);
	G3273<= not (I6448 and I6449);
	G3304<= not (I6468 and I6469);
	G3322<= not (I6488 and I6489);
	G3460<= not (I6665 and I6666);
	G3524<= not (G3209 and G3221);
	G3529<= not (G2310 and G3062 and G2325);
	G3530<= not (I6715 and I6716);
	G3585<= not (I6747 and I6748);
	G3623<= not (I6761 and I6762);
	G3625<= not (I6771 and I6772);
	G3626<= not (I6778 and I6779);
	G3631<= not (I6793 and I6794);
	G3634<= not (I6806 and I6807);
	G3662<= not (I6826 and I6827);
	G3681<= not (I6837 and I6838);
	G3717<= not (I6880 and I6881);
	G3734<= not (G3039 and G599);
	G3753<= not (G2382 and G2364 and G2800);
	G3766<= not (G2439 and G3222 and G2493);
	G3771<= not (I6989 and I6990);
	G3813<= not (I7034 and I7035);
	G3818<= not (G3056 and G3071 and G2310 and G3003);
	G3978<= not (G3207 and G1822);
	G3992<= not (G2571 and G2550 and G2990);
	G4088<= not (I7224 and I7225);
	G4104<= not (G3215 and G3247 and G2439 and G3200);
	G4117<= not (G3041 and G3061);
	G4130<= not (G3044 and G2518);
	G4144<= not (G2160 and G3044);
	G4168<= not (I7322 and I7323);
	G4297<= not (I7563 and I7564);
	G4374<= not (I7684 and I7685);
	G4476<= not (G3807 and G3071);
	G4482<= not (I7864 and I7865);
	G4488<= not (I7876 and I7877);
	G4538<= not (G3475 and G2399);
	G4588<= not (G3440 and G2745);
	G4675<= not (G4073 and G3247);
	G4749<= not (G3710 and G2061);
	G4803<= not (G3664 and G2356);
	G4821<= not (I8179 and I8180);
	G4976<= not (G2310 and G4604 and G3807);
	G5013<= not (G4749 and G3247 and G3205);
	G5103<= not (I8480 and I8481);
	G5118<= not (G2439 and G4806 and G4073);
	G5119<= not (I8514 and I8515);
	G5125<= not (I8528 and I8529);
	G5147<= not (I8544 and I8545);
	G5171<= not (I8562 and I8563);
	G5179<= not (I8576 and I8577);
	G5187<= not (I8590 and I8591);
	G5196<= not (I8605 and I8606);
	G5209<= not (I8625 and I8626);
	G5217<= not (I8641 and I8642);
	G5219<= not (I8651 and I8652);
	G5225<= not (I8663 and I8664);
	G5226<= not (I8670 and I8671);
	G5227<= not (I8677 and I8678);
	G5269<= not (I8716 and I8717);
	G5274<= not (I8729 and I8730);
	G5277<= not (G3734 and G4538);
	G5278<= not (I8739 and I8740);
	G5286<= not (I8751 and I8752);
	G5295<= not (I8762 and I8763);
	G5300<= not (I8771 and I8772);
	G5304<= not (I8779 and I8780);
	G5308<= not (I8787 and I8788);
	G5317<= not (I8796 and I8797);
	G5319<= not (I8804 and I8805);
	G5527<= not (G3978 and G4749);
	G5548<= not (G1840 and G4401);
	G5552<= not (G4777 and G4401);
	G5557<= not (G4538 and G3071 and G3011);
	G5592<= not (I9007 and I9008);
	G5935<= not (I9558 and I9559);
	G5942<= not (I9575 and I9576);
	G6003<= not (G5552 and G5548);
	G6019<= not (G617 and G4921);
	G6027<= not (G4566 and G4921);
	G6207<= not (I9947 and I9948);
	G6488<= not (G6027 and G6019);
	G6548<= not (G6132 and G6124 and G6122);
	G6573<= not (I10508 and I10509);
	G6577<= not (I10520 and I10521);
	G6740<= not (G6131 and G2550);
	G6758<= not (I10770 and I10771);
	G6858<= not (I10931 and I10932);
	G7054<= not (I11242 and I11243);
	G7062<= not (I11262 and I11263);
	G7067<= not (I11279 and I11280);
	G7101<= not (G6617 and G2364);
	G7269<= not (I11509 and I11510);
	G7523<= not (I11908 and I11909);
	G7524<= not (I11915 and I11916);
	G7533<= not (I11936 and I11937);
	G7547<= not (I11974 and I11975);
	G7548<= not (I11981 and I11982);
	G7557<= not (I11996 and I11997);
	G7558<= not (I12003 and I12004);
	G7567<= not (I12020 and I12021);
	G7572<= not (I12039 and I12040);
	G7573<= not (I12046 and I12047);
	G7582<= not (I12061 and I12062);
	G7583<= not (I12068 and I12069);
	G7584<= not (I12075 and I12076);
	G7587<= not (I12086 and I12087);
	G7588<= not (I12093 and I12094);
	G7592<= not (I12107 and I12108);
	G7593<= not (I12114 and I12115);
	G7596<= not (I12127 and I12128);
	G7598<= not (I12137 and I12138);
	G7599<= not (I12144 and I12145);
	G7624<= not (I12215 and I12216);
	G7671<= not (G7011 and G6995 and G6984 and G6974);
	G7717<= not (G6863 and G3206);
	G7932<= not (G7395 and G6847 and G7279 and G7273);
	G7934<= not (G7395 and G6847 and G7279 and G7369);
	G7942<= not (G7395 and G6847 and G7380 and G7369);
	G7947<= not (G7395 and G7390 and G7279 and G7369);
	G7950<= not (G7395 and G7390 and G7380 and G7273);
	G7953<= not (G7395 and G7390 and G7380 and G7369);
	G7960<= not (G7409 and G5573);
	G7978<= not (G7697 and G3038);
	G7986<= not (G7011 and G6995 and G6984 and G7550);
	G7987<= not (G7011 and G6995 and G7562 and G6974);
	G7990<= not (G7011 and G6995 and G7562 and G7550);
	G7992<= not (G7011 and G7574 and G6984 and G6974);
	G7994<= not (G7011 and G7574 and G6984 and G7550);
	G7996<= not (G7011 and G7574 and G7562 and G6974);
	G8000<= not (G7011 and G7574 and G7562 and G7550);
	G8006<= not (G5552 and G7717);
	G8109<= not (G5052 and G7853);
	G8177<= not (I13077 and I13078);
	G8180<= not (I13090 and I13091);
	G8190<= not (G6027 and G7978);
	G8298<= not (I13249 and I13250);
	G8300<= not (I13259 and I13260);
	G8301<= not (I13266 and I13267);
	G8302<= not (I13273 and I13274);
	G8305<= not (I13284 and I13285);
	G8307<= not (I13294 and I13295);
	G8308<= not (I13301 and I13302);
	G8309<= not (I13308 and I13309);
	G8402<= not (I13505 and I13506);
	G8405<= not (I13514 and I13515);
	G8407<= not (I13522 and I13523);
	G8409<= not (I13530 and I13531);
	G8411<= not (I13538 and I13539);
	G8412<= not (I13545 and I13546);
	G8414<= not (I13553 and I13554);
	G8415<= not (I13560 and I13561);
	G8471<= not (I13660 and I13661);
	G8501<= not (G3760 and G8366);
	G8502<= not (G2382 and G605 and G591 and G8366);
	G8506<= not (G3475 and G8366);
	G8507<= not (G3738 and G8366);
	G8511<= not (G5277 and G8366);
	G8512<= not (G3723 and G8366);
	G8541<= not (G4001 and G8390);
	G8542<= not (G2571 and G1828 and G1814 and G8390);
	G8545<= not (G3710 and G8390);
	G8546<= not (G3983 and G8390);
	G8549<= not (G5527 and G8390);
	G8551<= not (G3967 and G8390);
	G8558<= not (I13766 and I13767);
	G8612<= not (I13858 and I13859);
	G8616<= not (I13868 and I13869);
	G8623<= not (I13877 and I13878);
	G8627<= not (I13887 and I13888);
	G8628<= not (I13894 and I13895);
	G8629<= not (I13901 and I13902);
	G8630<= not (I13908 and I13909);
	G8705<= not (I13991 and I13992);
	G8737<= not (G2317 and G4921 and G8688);
	G8738<= not (G8688 and G4921);
	G8743<= not (G8617 and G6971 and G6964);
	G8744<= not (G8617 and G6509 and G6971);
	G8745<= not (G8617 and G6517 and G6964);
	G8746<= not (G8617 and G6517 and G6509);
	G8757<= not (G8599 and G4401);
	G8824<= not (G8502 and G8501 and G8739);
	G8825<= not (G8502 and G8738 and G8506);
	G8826<= not (G8739 and G8737 and G8648);
	G8839<= not (G8750 and G4401);
	G8840<= not (G8542 and G8541 and G8760);
	G8843<= not (G8542 and G8757 and G8545);
	G8847<= not (G8760 and G8683);
	G8880<= not (I14203 and I14204);
	G8881<= not (I14210 and I14211);
	G8882<= not (I14217 and I14218);
	G8932<= not (I14264 and I14265);
	G8933<= not (I14271 and I14272);
	G8934<= not (I14278 and I14279);
	G8942<= not (G8823 and G4921);
	G8970<= not (G5548 and G8839);
	G9107<= not (I14443 and I14444);
	G9204<= not (G6019 and G8942);
	G9413<= not (I14613 and I14614);
	G10043<= not (I15257 and I15258);
	G10144<= not (I15431 and I15432);
	G10149<= not (I15442 and I15443);
	G10153<= not (I15452 and I15453);
	G10229<= not (I15608 and I15609);
	G10231<= not (I15616 and I15617);
	G10302<= not (I15717 and I15718);
	G10366<= not (G10285 and G5392);
	G10384<= not (I15871 and I15872);
	G10386<= not (I15879 and I15880);
	G10392<= not (I15891 and I15892);
	G10394<= not (I15899 and I15900);
	G10396<= not (I15907 and I15908);
	G10440<= not (G10360 and G6037);
	G10446<= not (G10443 and G5350);
	G10447<= not (G10363 and G5360);
	G10467<= not (I15993 and I15994);
	G10468<= not (I16000 and I16001);
	G10469<= not (G10430 and G5999);
	G10470<= not (I16008 and I16009);
	G10472<= not (I16016 and I16017);
	G10474<= not (I16024 and I16025);
	G10475<= not (I16031 and I16032);
	G10476<= not (I16038 and I16039);
	G10477<= not (I16045 and I16046);
	G10478<= not (I16052 and I16053);
	G10479<= not (I16059 and I16060);
	G10480<= not (I16066 and I16067);
	G10481<= not (I16073 and I16074);
	G10482<= not (I16080 and I16081);
	G10483<= not (I16087 and I16088);
	G10505<= not (G10432 and G5938);
	G10507<= not (G10434 and G5859);
	G10509<= not (G10436 and G6023);
	G10511<= not (G10438 and G6032);
	G10513<= not (G10441 and G5345);
	G10665<= not (I16331 and I16332);
	G10779<= not (I16468 and I16469);
	G10853<= not (G10731 and G5034);
	G10886<= not (G10807 and G10805);
	G11276<= not (I17052 and I17053);
	G11414<= not (I17282 and I17283);
	G11415<= not (I17289 and I17290);
	G11416<= not (I17296 and I17297);
	G11418<= not (I17306 and I17307);
	G11448<= not (I17394 and I17395);
	G11449<= not (I17401 and I17402);
	G11474<= not (I17460 and I17461);
	G11490<= not (I17486 and I17487);
	G11491<= not (I17493 and I17494);
	G11496<= not (I17504 and I17505);
	G11538<= not (I17568 and I17569);
	G11549<= not (I17585 and I17586);
	I4910<= not (G386 and G318);
	I4911<= not (G386 and I4910);
	I4912<= not (G318 and I4910);
	I4928<= not (G391 and G321);
	I4929<= not (G391 and I4928);
	I4930<= not (G321 and I4928);
	I4941<= not (G396 and G324);
	I4942<= not (G396 and I4941);
	I4943<= not (G324 and I4941);
	I4954<= not (G401 and G327);
	I4955<= not (G401 and I4954);
	I4956<= not (G327 and I4954);
	I4964<= not (G406 and G330);
	I4965<= not (G406 and I4964);
	I4966<= not (G330 and I4964);
	I4971<= not (G991 and G995);
	I4972<= not (G991 and I4971);
	I4973<= not (G995 and I4971);
	I4978<= not (G411 and G333);
	I4979<= not (G411 and I4978);
	I4980<= not (G333 and I4978);
	I4985<= not (G999 and G1003);
	I4986<= not (G999 and I4985);
	I4987<= not (G1003 and I4985);
	I4995<= not (G416 and G309);
	I4996<= not (G416 and I4995);
	I4997<= not (G309 and I4995);
	I5005<= not (G421 and G312);
	I5006<= not (G421 and I5005);
	I5007<= not (G312 and I5005);
	I5013<= not (G1007 and G1011);
	I5014<= not (G1007 and I5013);
	I5015<= not (G1011 and I5013);
	I5023<= not (G995 and G1275);
	I5024<= not (G995 and I5023);
	I5025<= not (G1275 and I5023);
	I5034<= not (G1015 and G1019);
	I5035<= not (G1015 and I5034);
	I5036<= not (G1019 and I5034);
	I5104<= not (G431 and G435);
	I5105<= not (G431 and I5104);
	I5106<= not (G435 and I5104);
	I5126<= not (G1386 and G1389);
	I5127<= not (G1386 and I5126);
	I5128<= not (G1389 and I5126);
	I5135<= not (G521 and G525);
	I5136<= not (G521 and I5135);
	I5137<= not (G525 and I5135);
	I5164<= not (G1508 and G1499);
	I5165<= not (G1508 and I5164);
	I5166<= not (G1499 and I5164);
	I5184<= not (G1415 and G1515);
	I5185<= not (G1415 and I5184);
	I5186<= not (G1515 and I5184);
	I5202<= not (G369 and G374);
	I5203<= not (G369 and I5202);
	I5204<= not (G374 and I5202);
	I5229<= not (G182 and G148);
	I5230<= not (G182 and I5229);
	I5231<= not (G148 and I5229);
	I5263<= not (G456 and G461);
	I5264<= not (G456 and I5263);
	I5265<= not (G461 and I5263);
	I5282<= not (G758 and G762);
	I5283<= not (G758 and I5282);
	I5284<= not (G762 and I5282);
	I5295<= not (G794 and G798);
	I5296<= not (G794 and I5295);
	I5297<= not (G798 and I5295);
	I5315<= not (G1032 and G1027);
	I5316<= not (G1032 and I5315);
	I5317<= not (G1027 and I5315);
	I5323<= not (G1336 and G1341);
	I5324<= not (G1336 and I5323);
	I5325<= not (G1341 and I5323);
	I5341<= not (G315 and G426);
	I5342<= not (G315 and I5341);
	I5343<= not (G426 and I5341);
	I5371<= not (G971 and G976);
	I5372<= not (G971 and I5371);
	I5373<= not (G976 and I5371);
	I5449<= not (G1235 and G991);
	I5450<= not (G1235 and I5449);
	I5451<= not (G991 and I5449);
	I5459<= not (G1240 and G1003);
	I5460<= not (G1240 and I5459);
	I5461<= not (G1003 and I5459);
	I5468<= not (G1245 and G999);
	I5469<= not (G1245 and I5468);
	I5470<= not (G999 and I5468);
	I5484<= not (G1250 and G1011);
	I5485<= not (G1250 and I5484);
	I5486<= not (G1011 and I5484);
	I5500<= not (G1255 and G1007);
	I5501<= not (G1255 and I5500);
	I5502<= not (G1007 and I5500);
	I5516<= not (G1260 and G1019);
	I5517<= not (G1260 and I5516);
	I5518<= not (G1019 and I5516);
	I5528<= not (G1265 and G1015);
	I5529<= not (G1265 and I5528);
	I5530<= not (G1015 and I5528);
	I5538<= not (G1270 and G1023);
	I5539<= not (G1270 and I5538);
	I5540<= not (G1023 and I5538);
	I5591<= not (G1696 and G1703);
	I5592<= not (G1696 and I5591);
	I5593<= not (G1703 and I5591);
	I5604<= not (G1149 and G1153);
	I5605<= not (G1149 and I5604);
	I5606<= not (G1153 and I5604);
	I5611<= not (G1280 and G1284);
	I5612<= not (G1280 and I5611);
	I5613<= not (G1284 and I5611);
	I5618<= not (G1766 and G1771);
	I5619<= not (G1766 and I5618);
	I5620<= not (G1771 and I5618);
	I5675<= not (G1218 and G1223);
	I5676<= not (G1218 and I5675);
	I5677<= not (G1223 and I5675);
	I5865<= not (G2107 and G2105);
	I5866<= not (G2107 and I5865);
	I5867<= not (G2105 and I5865);
	I5878<= not (G2120 and G2115);
	I5879<= not (G2120 and I5878);
	I5880<= not (G2115 and I5878);
	I5891<= not (G750 and G2057);
	I5892<= not (G750 and I5891);
	I5893<= not (G2057 and I5891);
	I6109<= not (G2205 and G1494);
	I6110<= not (G2205 and I6109);
	I6111<= not (G1494 and I6109);
	I6124<= not (G2215 and G1419);
	I6125<= not (G2215 and I6124);
	I6126<= not (G1419 and I6124);
	I6136<= not (G2496 and G378);
	I6137<= not (G2496 and I6136);
	I6138<= not (G378 and I6136);
	I6143<= not (G1976 and G646);
	I6144<= not (G1976 and I6143);
	I6145<= not (G646 and I6143);
	I6166<= not (G2236 and G153);
	I6167<= not (G2236 and I6166);
	I6168<= not (G153 and I6166);
	I6176<= not (G2177 and G197);
	I6177<= not (G2177 and I6176);
	I6178<= not (G197 and I6176);
	I6186<= not (G2511 and G466);
	I6187<= not (G2511 and I6186);
	I6188<= not (G466 and I6186);
	I6199<= not (G2525 and G766);
	I6200<= not (G2525 and I6199);
	I6201<= not (G766 and I6199);
	I6207<= not (G2534 and G802);
	I6208<= not (G2534 and I6207);
	I6209<= not (G802 and I6207);
	I6224<= not (G2544 and G1346);
	I6225<= not (G2544 and I6224);
	I6226<= not (G1346 and I6224);
	I6287<= not (G2091 and G981);
	I6288<= not (G2091 and I6287);
	I6289<= not (G981 and I6287);
	I6322<= not (G2050 and G1864);
	I6323<= not (G2050 and I6322);
	I6324<= not (G1864 and I6322);
	I6447<= not (G2264 and G1776);
	I6448<= not (G2264 and I6447);
	I6449<= not (G1776 and I6447);
	I6467<= not (G23 and G2479);
	I6468<= not (G23 and I6467);
	I6469<= not (G2479 and I6467);
	I6487<= not (G2306 and G1227);
	I6488<= not (G2306 and I6487);
	I6489<= not (G1227 and I6487);
	I6664<= not (G2792 and G2776);
	I6665<= not (G2792 and I6664);
	I6666<= not (G2776 and I6664);
	I6714<= not (G2961 and G201);
	I6715<= not (G2961 and I6714);
	I6716<= not (G201 and I6714);
	I6746<= not (G2938 and G1453);
	I6747<= not (G2938 and I6746);
	I6748<= not (G1453 and I6746);
	I6760<= not (G2943 and G1448);
	I6761<= not (G2943 and I6760);
	I6762<= not (G1448 and I6760);
	I6770<= not (G3257 and G382);
	I6771<= not (G3257 and I6770);
	I6772<= not (G382 and I6770);
	I6777<= not (G2892 and G650);
	I6778<= not (G2892 and I6777);
	I6779<= not (G650 and I6777);
	I6792<= not (G2959 and G143);
	I6793<= not (G2959 and I6792);
	I6794<= not (G143 and I6792);
	I6805<= not (G3268 and G471);
	I6806<= not (G3268 and I6805);
	I6807<= not (G471 and I6805);
	I6825<= not (G3281 and G770);
	I6826<= not (G3281 and I6825);
	I6827<= not (G770 and I6825);
	I6836<= not (G3287 and G806);
	I6837<= not (G3287 and I6836);
	I6838<= not (G806 and I6836);
	I6879<= not (G3301 and G1351);
	I6880<= not (G3301 and I6879);
	I6881<= not (G1351 and I6879);
	I6988<= not (G2760 and G986);
	I6989<= not (G2760 and I6988);
	I6990<= not (G986 and I6988);
	I7033<= not (G3089 and G1868);
	I7034<= not (G3089 and I7033);
	I7035<= not (G1868 and I7033);
	I7223<= not (G2981 and G1781);
	I7224<= not (G2981 and I7223);
	I7225<= not (G1781 and I7223);
	I7321<= not (G3047 and G1231);
	I7322<= not (G3047 and I7321);
	I7323<= not (G1231 and I7321);
	I7562<= not (G3533 and G654);
	I7563<= not (G3533 and I7562);
	I7564<= not (G654 and I7562);
	I7683<= not (G1023 and G3460);
	I7684<= not (G1023 and I7683);
	I7685<= not (G3460 and I7683);
	I7863<= not (G4099 and G774);
	I7864<= not (G4099 and I7863);
	I7865<= not (G774 and I7863);
	I7875<= not (G4109 and G810);
	I7876<= not (G4109 and I7875);
	I7877<= not (G810 and I7875);
	I8178<= not (G3685 and G1786);
	I8179<= not (G3685 and I8178);
	I8180<= not (G1786 and I8178);
	I8479<= not (G4455 and G3530);
	I8480<= not (G4455 and I8479);
	I8481<= not (G3530 and I8479);
	I8513<= not (G4873 and G3513);
	I8514<= not (G4873 and I8513);
	I8515<= not (G3513 and I8513);
	I8527<= not (G4879 and G481);
	I8528<= not (G4879 and I8527);
	I8529<= not (G481 and I8527);
	I8543<= not (G4218 and G486);
	I8544<= not (G4218 and I8543);
	I8545<= not (G486 and I8543);
	I8561<= not (G4227 and G491);
	I8562<= not (G4227 and I8561);
	I8563<= not (G491 and I8561);
	I8575<= not (G4234 and G496);
	I8576<= not (G4234 and I8575);
	I8577<= not (G496 and I8575);
	I8589<= not (G4251 and G501);
	I8590<= not (G4251 and I8589);
	I8591<= not (G501 and I8589);
	I8604<= not (G4259 and G506);
	I8605<= not (G4259 and I8604);
	I8606<= not (G506 and I8604);
	I8624<= not (G4267 and G511);
	I8625<= not (G4267 and I8624);
	I8626<= not (G511 and I8624);
	I8640<= not (G4278 and G516);
	I8641<= not (G4278 and I8640);
	I8642<= not (G516 and I8640);
	I8650<= not (G4824 and G778);
	I8651<= not (G4824 and I8650);
	I8652<= not (G778 and I8650);
	I8662<= not (G4286 and G476);
	I8663<= not (G4286 and I8662);
	I8664<= not (G476 and I8662);
	I8669<= not (G4831 and G814);
	I8670<= not (G4831 and I8669);
	I8671<= not (G814 and I8669);
	I8676<= not (G4374 and G1027);
	I8677<= not (G4374 and I8676);
	I8678<= not (G1027 and I8676);
	I8715<= not (G4601 and G4052);
	I8716<= not (G4601 and I8715);
	I8717<= not (G4052 and I8715);
	I8728<= not (G4605 and G1117);
	I8729<= not (G4605 and I8728);
	I8730<= not (G1117 and I8728);
	I8738<= not (G4607 and G1121);
	I8739<= not (G4607 and I8738);
	I8740<= not (G1121 and I8738);
	I8750<= not (G4613 and G1125);
	I8751<= not (G4613 and I8750);
	I8752<= not (G1125 and I8750);
	I8761<= not (G4616 and G1129);
	I8762<= not (G4616 and I8761);
	I8763<= not (G1129 and I8761);
	I8770<= not (G4619 and G1133);
	I8771<= not (G4619 and I8770);
	I8772<= not (G1133 and I8770);
	I8778<= not (G4630 and G1137);
	I8779<= not (G4630 and I8778);
	I8780<= not (G1137 and I8778);
	I8786<= not (G4639 and G1141);
	I8787<= not (G4639 and I8786);
	I8788<= not (G1141 and I8786);
	I8795<= not (G4672 and G1145);
	I8796<= not (G4672 and I8795);
	I8797<= not (G1145 and I8795);
	I8803<= not (G4677 and G1113);
	I8804<= not (G4677 and I8803);
	I8805<= not (G1113 and I8803);
	I9006<= not (G4492 and G1791);
	I9007<= not (G4492 and I9006);
	I9008<= not (G1791 and I9006);
	I9557<= not (G5598 and G782);
	I9558<= not (G5598 and I9557);
	I9559<= not (G782 and I9557);
	I9574<= not (G5608 and G818);
	I9575<= not (G5608 and I9574);
	I9576<= not (G818 and I9574);
	I9946<= not (G5233 and G1796);
	I9947<= not (G5233 and I9946);
	I9948<= not (G1796 and I9946);
	I10507<= not (G6221 and G786);
	I10508<= not (G6221 and I10507);
	I10509<= not (G786 and I10507);
	I10519<= not (G6231 and G822);
	I10520<= not (G6231 and I10519);
	I10521<= not (G822 and I10519);
	I10769<= not (G5944 and G1801);
	I10770<= not (G5944 and I10769);
	I10771<= not (G1801 and I10769);
	I10930<= not (G6395 and G5555);
	I10931<= not (G6395 and I10930);
	I10932<= not (G5555 and I10930);
	I11241<= not (G6760 and G790);
	I11242<= not (G6760 and I11241);
	I11243<= not (G790 and I11241);
	I11261<= not (G6775 and G826);
	I11262<= not (G6775 and I11261);
	I11263<= not (G826 and I11261);
	I11278<= not (G305 and G6485);
	I11279<= not (G305 and I11278);
	I11280<= not (G6485 and I11278);
	I11508<= not (G6580 and G1806);
	I11509<= not (G6580 and I11508);
	I11510<= not (G1806 and I11508);
	I11907<= not (G6967 and G1474);
	I11908<= not (G6967 and I11907);
	I11909<= not (G1474 and I11907);
	I11914<= not (G6935 and G1494);
	I11915<= not (G6935 and I11914);
	I11916<= not (G1494 and I11914);
	I11935<= not (G7004 and G1458);
	I11936<= not (G7004 and I11935);
	I11937<= not (G1458 and I11935);
	I11973<= not (G7001 and G1462);
	I11974<= not (G7001 and I11973);
	I11975<= not (G1462 and I11973);
	I11980<= not (G6957 and G1482);
	I11981<= not (G6957 and I11980);
	I11982<= not (G1482 and I11980);
	I11995<= not (G7107 and G127);
	I11996<= not (G7107 and I11995);
	I11997<= not (G127 and I11995);
	I12002<= not (G7082 and G153);
	I12003<= not (G7082 and I12002);
	I12004<= not (G153 and I12002);
	I12019<= not (G7119 and G166);
	I12020<= not (G7119 and I12019);
	I12021<= not (G166 and I12019);
	I12038<= not (G6990 and G1466);
	I12039<= not (G6990 and I12038);
	I12040<= not (G1466 and I12038);
	I12045<= not (G6951 and G1486);
	I12046<= not (G6951 and I12045);
	I12047<= not (G1486 and I12045);
	I12060<= not (G6961 and G1478);
	I12061<= not (G6961 and I12060);
	I12062<= not (G1478 and I12060);
	I12067<= not (G7116 and G139);
	I12068<= not (G7116 and I12067);
	I12069<= not (G139 and I12067);
	I12074<= not (G7098 and G174);
	I12075<= not (G7098 and I12074);
	I12076<= not (G174 and I12074);
	I12085<= not (G6980 and G1470);
	I12086<= not (G6980 and I12085);
	I12087<= not (G1470 and I12085);
	I12092<= not (G6944 and G1490);
	I12093<= not (G6944 and I12092);
	I12094<= not (G1490 and I12092);
	I12106<= not (G7113 and G135);
	I12107<= not (G7113 and I12106);
	I12108<= not (G135 and I12106);
	I12113<= not (G7093 and G162);
	I12114<= not (G7093 and I12113);
	I12115<= not (G162 and I12113);
	I12126<= not (G7103 and G170);
	I12127<= not (G7103 and I12126);
	I12128<= not (G170 and I12126);
	I12136<= not (G7110 and G131);
	I12137<= not (G7110 and I12136);
	I12138<= not (G131 and I12136);
	I12143<= not (G7089 and G158);
	I12144<= not (G7089 and I12143);
	I12145<= not (G158 and I12143);
	I12214<= not (G7061 and G2518);
	I12215<= not (G7061 and I12214);
	I12216<= not (G2518 and I12214);
	I13076<= not (G1872 and G7963);
	I13077<= not (G1872 and I13076);
	I13078<= not (G7963 and I13076);
	I13089<= not (G8006 and G1840);
	I13090<= not (G8006 and I13089);
	I13091<= not (G1840 and I13089);
	I13248<= not (G1891 and G8148);
	I13249<= not (G1891 and I13248);
	I13250<= not (G8148 and I13248);
	I13258<= not (G1900 and G8153);
	I13259<= not (G1900 and I13258);
	I13260<= not (G8153 and I13258);
	I13265<= not (G1909 and G8154);
	I13266<= not (G1909 and I13265);
	I13267<= not (G8154 and I13265);
	I13272<= not (G1918 and G8158);
	I13273<= not (G1918 and I13272);
	I13274<= not (G8158 and I13272);
	I13283<= not (G1927 and G8159);
	I13284<= not (G1927 and I13283);
	I13285<= not (G8159 and I13283);
	I13293<= not (G1882 and G8161);
	I13294<= not (G1882 and I13293);
	I13295<= not (G8161 and I13293);
	I13300<= not (G1936 and G8162);
	I13301<= not (G1936 and I13300);
	I13302<= not (G8162 and I13300);
	I13307<= not (G8190 and G617);
	I13308<= not (G8190 and I13307);
	I13309<= not (G617 and I13307);
	I13504<= not (G677 and G8247);
	I13505<= not (G677 and I13504);
	I13506<= not (G8247 and I13504);
	I13513<= not (G686 and G8248);
	I13514<= not (G686 and I13513);
	I13515<= not (G8248 and I13513);
	I13521<= not (G695 and G8249);
	I13522<= not (G695 and I13521);
	I13523<= not (G8249 and I13521);
	I13529<= not (G704 and G8253);
	I13530<= not (G704 and I13529);
	I13531<= not (G8253 and I13529);
	I13537<= not (G658 and G8157);
	I13538<= not (G658 and I13537);
	I13539<= not (G8157 and I13537);
	I13544<= not (G713 and G8259);
	I13545<= not (G713 and I13544);
	I13546<= not (G8259 and I13544);
	I13552<= not (G668 and G8262);
	I13553<= not (G668 and I13552);
	I13554<= not (G8262 and I13552);
	I13559<= not (G722 and G8263);
	I13560<= not (G722 and I13559);
	I13561<= not (G8263 and I13559);
	I13659<= not (G1945 and G8322);
	I13660<= not (G1945 and I13659);
	I13661<= not (G8322 and I13659);
	I13765<= not (G731 and G8417);
	I13766<= not (G731 and I13765);
	I13767<= not (G8417 and I13765);
	I13857<= not (G8538 and G1448);
	I13858<= not (G8538 and I13857);
	I13859<= not (G1448 and I13857);
	I13867<= not (G8523 and G1403);
	I13868<= not (G8523 and I13867);
	I13869<= not (G1403 and I13867);
	I13876<= not (G8535 and G1444);
	I13877<= not (G8535 and I13876);
	I13878<= not (G1444 and I13876);
	I13886<= not (G8532 and G1440);
	I13887<= not (G8532 and I13886);
	I13888<= not (G1440 and I13886);
	I13893<= not (G8529 and G1436);
	I13894<= not (G8529 and I13893);
	I13895<= not (G1436 and I13893);
	I13900<= not (G8520 and G1428);
	I13901<= not (G8520 and I13900);
	I13902<= not (G1428 and I13900);
	I13907<= not (G8526 and G1432);
	I13908<= not (G8526 and I13907);
	I13909<= not (G1432 and I13907);
	I13990<= not (G622 and G8688);
	I13991<= not (G622 and I13990);
	I13992<= not (G8688 and I13990);
	I14202<= not (G8825 and G591);
	I14203<= not (G8825 and I14202);
	I14204<= not (G591 and I14202);
	I14209<= not (G8824 and G599);
	I14210<= not (G8824 and I14209);
	I14211<= not (G599 and I14209);
	I14216<= not (G8826 and G605);
	I14217<= not (G8826 and I14216);
	I14218<= not (G605 and I14216);
	I14263<= not (G8843 and G1814);
	I14264<= not (G8843 and I14263);
	I14265<= not (G1814 and I14263);
	I14270<= not (G8840 and G1822);
	I14271<= not (G8840 and I14270);
	I14272<= not (G1822 and I14270);
	I14277<= not (G8847 and G1828);
	I14278<= not (G8847 and I14277);
	I14279<= not (G1828 and I14277);
	I14442<= not (G8970 and G1834);
	I14443<= not (G8970 and I14442);
	I14444<= not (G1834 and I14442);
	I14612<= not (G9204 and G611);
	I14613<= not (G9204 and I14612);
	I14614<= not (G611 and I14612);
	I15256<= not (G9984 and G9980);
	I15257<= not (G9984 and I15256);
	I15258<= not (G9980 and I15256);
	I15430<= not (G10047 and G10044);
	I15431<= not (G10047 and I15430);
	I15432<= not (G10044 and I15430);
	I15441<= not (G10035 and G10122);
	I15442<= not (G10035 and I15441);
	I15443<= not (G10122 and I15441);
	I15451<= not (G10058 and G10051);
	I15452<= not (G10058 and I15451);
	I15453<= not (G10051 and I15451);
	I15607<= not (G10149 and G10144);
	I15608<= not (G10149 and I15607);
	I15609<= not (G10144 and I15607);
	I15615<= not (G10043 and G10153);
	I15616<= not (G10043 and I15615);
	I15617<= not (G10153 and I15615);
	I15716<= not (G10231 and G10229);
	I15717<= not (G10231 and I15716);
	I15718<= not (G10229 and I15716);
	I15870<= not (G10358 and G2713);
	I15871<= not (G10358 and I15870);
	I15872<= not (G2713 and I15870);
	I15878<= not (G10359 and G2719);
	I15879<= not (G10359 and I15878);
	I15880<= not (G2719 and I15878);
	I15890<= not (G853 and G10286);
	I15891<= not (G853 and I15890);
	I15892<= not (G10286 and I15890);
	I15898<= not (G857 and G10287);
	I15899<= not (G857 and I15898);
	I15900<= not (G10287 and I15898);
	I15906<= not (G6899 and G10302);
	I15907<= not (G6899 and I15906);
	I15908<= not (G10302 and I15906);
	I15992<= not (G10422 and G2677);
	I15993<= not (G10422 and I15992);
	I15994<= not (G2677 and I15992);
	I15999<= not (G10423 and G2683);
	I16000<= not (G10423 and I15999);
	I16001<= not (G2683 and I15999);
	I16007<= not (G10424 and G2689);
	I16008<= not (G10424 and I16007);
	I16009<= not (G2689 and I16007);
	I16015<= not (G10425 and G2695);
	I16016<= not (G10425 and I16015);
	I16017<= not (G2695 and I16015);
	I16023<= not (G10426 and G2701);
	I16024<= not (G10426 and I16023);
	I16025<= not (G2701 and I16023);
	I16030<= not (G829 and G10368);
	I16031<= not (G829 and I16030);
	I16032<= not (G10368 and I16030);
	I16037<= not (G10427 and G2707);
	I16038<= not (G10427 and I16037);
	I16039<= not (G2707 and I16037);
	I16044<= not (G833 and G10370);
	I16045<= not (G833 and I16044);
	I16046<= not (G10370 and I16044);
	I16051<= not (G837 and G10371);
	I16052<= not (G837 and I16051);
	I16053<= not (G10371 and I16051);
	I16058<= not (G841 and G10372);
	I16059<= not (G841 and I16058);
	I16060<= not (G10372 and I16058);
	I16065<= not (G10428 and G2765);
	I16066<= not (G10428 and I16065);
	I16067<= not (G2765 and I16065);
	I16072<= not (G845 and G10373);
	I16073<= not (G845 and I16072);
	I16074<= not (G10373 and I16072);
	I16079<= not (G849 and G10374);
	I16080<= not (G849 and I16079);
	I16081<= not (G10374 and I16079);
	I16086<= not (G861 and G10375);
	I16087<= not (G861 and I16086);
	I16088<= not (G10375 and I16086);
	I16330<= not (G10616 and G4997);
	I16331<= not (G10616 and I16330);
	I16332<= not (G4997 and I16330);
	I16467<= not (G10716 and G10518);
	I16468<= not (G10716 and I16467);
	I16469<= not (G10518 and I16467);
	I17051<= not (G10923 and G11249);
	I17052<= not (G10923 and I17051);
	I17053<= not (G11249 and I17051);
	I17281<= not (G11360 and G11357);
	I17282<= not (G11360 and I17281);
	I17283<= not (G11357 and I17281);
	I17288<= not (G11366 and G11363);
	I17289<= not (G11366 and I17288);
	I17290<= not (G11363 and I17288);
	I17295<= not (G11373 and G11369);
	I17296<= not (G11373 and I17295);
	I17297<= not (G11369 and I17295);
	I17305<= not (G11381 and G11377);
	I17306<= not (G11381 and I17305);
	I17307<= not (G11377 and I17305);
	I17393<= not (G11415 and G11414);
	I17394<= not (G11415 and I17393);
	I17395<= not (G11414 and I17393);
	I17400<= not (G11418 and G11416);
	I17401<= not (G11418 and I17400);
	I17402<= not (G11416 and I17400);
	I17459<= not (G11449 and G11448);
	I17460<= not (G11449 and I17459);
	I17461<= not (G11448 and I17459);
	I17485<= not (G11384 and G11474);
	I17486<= not (G11384 and I17485);
	I17487<= not (G11474 and I17485);
	I17492<= not (G11475 and G3623);
	I17493<= not (G11475 and I17492);
	I17494<= not (G3623 and I17492);
	I17503<= not (G11475 and G7603);
	I17504<= not (G11475 and I17503);
	I17505<= not (G7603 and I17503);
	I17567<= not (G11496 and G1610);
	I17568<= not (G11496 and I17567);
	I17569<= not (G1610 and I17567);
	I17584<= not (G11354 and G11515);
	I17585<= not (G11354 and I17584);
	I17586<= not (G11515 and I17584);
	G2204<=G1393 or G1394;
	G2305<=I5351 or I5352;
	G2309<=I5357 or I5358;
	G2315<=G1163 or G1166 or G1113 or I5363;
	G2316<=G1300 or G1304 or G1270 or I5366;
	G2353<=G1403 or G1407 or G1411 or G1415;
	G2499<=I5570 or I5571;
	G2501<=G448 or G452 or G421 or I5576;
	G2514<=I5599 or I5600;
	G2521<=G538 or G542 or G476 or I5626;
	G2522<=G833 or G829 or I5629;
	G2528<=G861 or G857 or G853 or G849;
	G2538<=G1466 or G1458 or I5649;
	G2744<=I5804 or I5805;
	G2984<=G2528 or G2522;
	G3120<=I6350 or I6351;
	G3354<=G2920 or G2124;
	G3399<=G2918 or G2940;
	G3414<=G2911 or G2917;
	G3425<=G2895 or G2910;
	G3431<=G2951 or G2957;
	G3435<=G2945 or G2950;
	G3438<=G2939 or G2944;
	G3513<=G3118 or G2180;
	G3584<=G2863 or G2516;
	G3688<=G3144 or G2454;
	G3698<=G3121 or G2480;
	G3819<=G3275 or G9;
	G3860<=G3107 or G2167;
	G3875<=G3275 or G12;
	G4052<=G2862 or G2515;
	G4089<=G1959 or G3318;
	G4231<=G3991 or G3998;
	G4238<=G3999 or G4007;
	G4239<=G4000 or G4008;
	G4255<=G4009 or G4047;
	G4264<=G4048 or G4053;
	G4274<=G4054 or G4058;
	G4283<=G4059 or G4063;
	G4293<=G4064 or G4068;
	G4300<=G3546 or G2391;
	G4309<=G4069 or G4079;
	G4556<=G3536 or G2916;
	G4609<=G3400 or G119;
	G4640<=G3348 or G3563 or G1527;
	G4682<=G3563 or G3348 or G1570;
	G4997<=G4581 or G4584;
	G5028<=G4836 or G4128;
	G5036<=G4871 or G4162;
	G5038<=G4878 or G4884;
	G5189<=G4345 or G3496;
	G5224<=G4360 or G3512;
	G5229<=G4364 or G3516;
	G5309<=G3664 or G4401;
	G5361<=G4316 or G4093 or G126;
	G5396<=G4481 or G3684;
	G5403<=G4486 or G3695;
	G5404<=G4487 or G3696;
	G5405<=G4476 or G3440;
	G5555<=G4389 or G4397;
	G5576<=G4675 or G3664;
	G5587<=G4714 or G3904;
	G5590<=G4718 or G4723;
	G5762<=G5178 or G5186;
	G5802<=G5601 or G4837;
	G5803<=G5575 or G4820;
	G5809<=G5611 or G4865;
	G5810<=G5588 or G4823;
	G5813<=G5617 or G4869;
	G5814<=G5591 or G4827;
	G5819<=G5625 or G4876;
	G5820<=G5595 or G4834;
	G5823<=G5631 or G4882;
	G5824<=G5602 or G4839;
	G5837<=G5640 or G4224;
	G5838<=G5612 or G4866;
	G5841<=G4914 or G4230;
	G5842<=G5618 or G4870;
	G5846<=G4932 or G4236;
	G5847<=G5626 or G4877;
	G5849<=G4949 or G4260;
	G5851<=G4941 or G4253;
	G5852<=G5632 or G4883;
	G5857<=G5418 or G4670;
	G5867<=G3440 or G4921;
	G5910<=G5023 or G4341;
	G5914<=G5029 or G4343;
	G5981<=G5074 or G4383;
	G5983<=G5084 or G4392;
	G5993<=G5090 or G4400;
	G5995<=G5097 or G5099;
	G5996<=G5473 or G3908;
	G6000<=G5480 or G3912;
	G6002<=G5489 or G3939;
	G6015<=G5497 or G3942;
	G6026<=G5507 or G3970;
	G6035<=G5518 or G3974;
	G6038<=G5528 or G3979;
	G6042<=G5535 or G3987;
	G6045<=G5541 or G3989;
	G6049<=G5254 or G3718;
	G6054<=G5199 or G4483;
	G6059<=G5211 or G4489;
	G6061<=G5204 or G4;
	G6068<=G5220 or G4497;
	G6071<=G5228 or G4505;
	G6074<=G5349 or G1;
	G6078<=G4503 or G5256;
	G6080<=G5249 or G4512;
	G6088<=G5260 or G4522;
	G6093<=G5264 or G4534;
	G6096<=G5268 or G4542;
	G6099<=G5273 or G4550;
	G6105<=G5279 or G4559;
	G6122<=G5172 or G5180;
	G6124<=G5181 or G5188;
	G6177<=G5444 or G4712;
	G6185<=G5470 or G4715;
	G6243<=G5537 or G4774;
	G6465<=G5825 or G5041;
	G6468<=G5690 or G4950;
	G6469<=G5698 or G4959;
	G6470<=G5699 or G4960;
	G6478<=G5706 or G4967;
	G6479<=G5707 or G4968;
	G6480<=G5721 or G4971;
	G6481<=G5722 or G4972;
	G6485<=G5848 or G5067;
	G6500<=G5725 or G4986;
	G6501<=G5726 or G4987;
	G6506<=G5731 or G4989;
	G6507<=G5732 or G4990;
	G6513<=G5737 or G4991;
	G6514<=G5738 or G4992;
	G6515<=G5739 or G4993;
	G6522<=G5744 or G4994;
	G6523<=G5745 or G4995;
	G6524<=G5746 or G4996;
	G6528<=G5756 or G4999;
	G6529<=G5757 or G5000;
	G6533<=G5771 or G5002;
	G6534<=G5772 or G5003;
	G6537<=G5781 or G5005;
	G6538<=G5782 or G5006;
	G6541<=G5788 or G5009;
	G6542<=G5789 or G5010;
	G6545<=G5795 or G5025;
	G6546<=G5796 or G5026;
	G6551<=G5804 or G5031;
	G6592<=G5100 or G5882;
	G6626<=G5934 or G123;
	G6672<=G5941 or G5259;
	G6739<=G5769 or G5780;
	G6755<=G6106 or G5479;
	G6777<=G5691 or G5052;
	G6894<=G6763 or G4868;
	G6895<=G6776 or G4875;
	G6897<=G6771 or G6240;
	G6898<=G6790 or G4881;
	G6899<=G6463 or G5471;
	G6900<=G6787 or G6246;
	G6901<=G6788 or G6247;
	G6902<=G6794 or G4223;
	G6906<=G6791 or G5674;
	G6907<=G6792 or G5675;
	G6908<=G6345 or G4229;
	G6909<=G6346 or G5684;
	G6910<=G6341 or G5680;
	G6911<=G6342 or G5681;
	G6912<=G6350 or G4235;
	G6915<=G6347 or G5686;
	G6916<=G6348 or G5687;
	G6918<=G6358 or G4252;
	G6922<=G6352 or G5694;
	G6923<=G6353 or G5695;
	G6924<=G6362 or G4261;
	G6928<=G6359 or G5703;
	G6929<=G6360 or G5704;
	G6930<=G6364 or G4269;
	G6934<=G6363 or G5720;
	G7075<=G5104 or G6530;
	G7092<=G6540 or G5902;
	G7096<=G6544 or G5911;
	G7102<=G6550 or G5915;
	G7106<=G6554 or G5917;
	G7133<=G6616 or G3067;
	G7143<=G6619 or G6039;
	G7183<=G6623 or G6046;
	G7184<=G6625 or G6047;
	G7189<=G6632 or G6053;
	G7203<=G6640 or G6058;
	G7204<=G6645 or G6062;
	G7211<=G6647 or G6067;
	G7218<=G6655 or G6070;
	G7219<=G6661 or G6076;
	G7225<=G6666 or G6079;
	G7231<=G6673 or G6087;
	G7236<=G6684 or G6092;
	G7240<=G6687 or G6095;
	G7242<=G6693 or G6098;
	G7244<=G6699 or G4720;
	G7245<=G6696 or G6102;
	G7246<=G6465 or G6003;
	G7257<=G6701 or G4725;
	G7258<=G6549 or G5913;
	G7265<=G6756 or G6204;
	G7290<=G7046 or G6316;
	G7291<=G7050 or G6317;
	G7292<=G7055 or G6318;
	G7293<=G7063 or G6319;
	G7294<=G7068 or G6320;
	G7295<=G7071 or G6321;
	G7296<=G7131 or G6322;
	G7297<=G7132 or G6323;
	G7298<=G7136 or G6324;
	G7299<=G7138 or G6325;
	G7300<=G7139 or G6326;
	G7301<=G7140 or G6327;
	G7302<=G7141 or G6328;
	G7303<=G7145 or G6329;
	G7367<=G7224 or G6744;
	G7375<=G7230 or G6745;
	G7384<=G7088 or G6618;
	G7385<=G7235 or G6746;
	G7441<=G7271 or G6789;
	G7457<=G6873 or G6404;
	G7465<=G6876 or G6410;
	G7471<=G6880 or G6416;
	G7478<=G6884 or G6423;
	G7503<=G6887 or G6430;
	G7510<=G7186 or G6730;
	G7511<=G6890 or G6438;
	G7621<=G5108 or G6994;
	G7626<=G7060 or G5267;
	G7638<=G7265 or G6488;
	G7651<=G7135 or G4084;
	G7660<=G7059 or G6583;
	G7664<=G6855 or G4084;
	G7712<=G7125 or G3540;
	G7738<=G7200 or G6738;
	G7740<=G7209 or G6741;
	G7742<=G7217 or G6743;
	G7846<=G7722 or G7241;
	G7926<=G7435 or G6892;
	G7963<=G7687 or G7182;
	G7971<=G5110 or G7549;
	G8148<=G7884 or G6872;
	G8153<=G7888 or G6875;
	G8154<=G7891 or G6879;
	G8157<=G7965 or G7623;
	G8158<=G7893 or G6883;
	G8159<=G7895 or G6886;
	G8161<=G8005 or G7185;
	G8162<=G7898 or G6889;
	G8187<=G7542 or G7998;
	G8193<=G5145 or G7937;
	G8194<=G5168 or G7940;
	G8199<=G7902 or G7444;
	G8200<=G7535 or G8008;
	G8203<=G7453 or G7999;
	G8206<=G7459 or G8007;
	G8210<=G7466 or G7995;
	G8214<=G7472 or G8004;
	G8221<=G7496 or G7993;
	G8226<=G7504 or G8002;
	G8230<=G7515 or G7991;
	G8236<=G7526 or G8001;
	G8241<=G7536 or G7989;
	G8247<=G8010 or G7704;
	G8248<=G8014 or G7707;
	G8249<=G8018 or G7710;
	G8252<=G7988 or G7679;
	G8253<=G8023 or G7718;
	G8259<=G8028 or G7719;
	G8261<=G7876 or G3383;
	G8262<=G7970 or G7625;
	G8263<=G8032 or G7720;
	G8264<=G7879 or G3389;
	G8265<=G7881 or G3396;
	G8266<=G7885 or G3412;
	G8267<=G7889 or G3422;
	G8268<=G7962 or G7613;
	G8269<=G7892 or G3429;
	G8270<=G7894 or G3434;
	G8281<=G8097 or G7818;
	G8282<=G8101 or G7819;
	G8283<=G8098 or G7820;
	G8284<=G8102 or G7821;
	G8285<=G8104 or G7822;
	G8286<=G8107 or G7823;
	G8287<=G8117 or G7824;
	G8288<=G8119 or G7825;
	G8322<=G8136 or G6891;
	G8377<=G8185 or G7958;
	G8383<=G8163 or G5051;
	G8417<=G8246 or G7721;
	G8428<=G8382 or G8068;
	G8429<=G8385 or G8069;
	G8430<=G8386 or G8070;
	G8431<=G8387 or G8071;
	G8432<=G8389 or G8072;
	G8433<=G8399 or G8073;
	G8434<=G8400 or G8074;
	G8435<=G8403 or G8075;
	G8451<=G3440 or G8366;
	G8488<=G3664 or G8390;
	G8552<=G8217 or G8388;
	G8559<=G8380 or G4731;
	G8574<=G5679 or G7853 or G8465;
	G8602<=G8401 or G8550;
	G8605<=G8404 or G8553;
	G8607<=G8406 or G8554;
	G8609<=G8408 or G8555;
	G8611<=G8410 or G8556;
	G8614<=G8365 or G8510;
	G8615<=G8413 or G8557;
	G8631<=G8474 or G7449;
	G8638<=G8108 or G8461;
	G8639<=G8118 or G8462;
	G8641<=G8120 or G8463;
	G8642<=G5236 or G5205 or G8465;
	G8643<=G8364 or G8508;
	G8644<=G8123 or G8464;
	G8645<=G8127 or G8469;
	G8646<=G8224 or G8547;
	G8647<=G8130 or G8470;
	G8649<=G8499 or G4519;
	G8715<=G8416 or G8687;
	G8742<=G8135 or G8598;
	G8770<=G5476 or G8651;
	G8771<=G5483 or G8652;
	G8773<=G5491 or G8653;
	G8774<=G5499 or G8654;
	G8776<=G5510 or G8655;
	G8777<=G5522 or G8659;
	G8779<=G5530 or G8663;
	G8806<=G7931 or G8718;
	G8810<=G7933 or G8720;
	G8811<=G7935 or G8722;
	G8812<=G7939 or G8724;
	G8813<=G7943 or G8726;
	G8814<=G7945 or G8728;
	G8815<=G7948 or G8730;
	G8816<=G7951 or G8731;
	G8817<=G7954 or G8732;
	G8818<=G7955 or G8733;
	G8819<=G7957 or G8734;
	G8823<=G8778 or G8693;
	G8883<=G8838 or G8753;
	G8885<=G8841 or G8754;
	G8887<=G8842 or G8755;
	G8889<=G8844 or G8756;
	G8920<=G8845 or G8759;
	G8921<=G8827 or G8748;
	G8922<=G8822 or G8736;
	G8923<=G8846 or G8763;
	G8926<=G8848 or G8764;
	G8937<=G8786 or G8698;
	G8938<=G8789 or G8699;
	G8939<=G8791 or G8701;
	G8940<=G8793 or G8703;
	G8941<=G8796 or G8706;
	G8943<=G8837 or G8749;
	G8944<=G8799 or G8708;
	G8945<=G8801 or G8710;
	G8973<=G8821 or G8735;
	G9088<=G8927 or G8381;
	G9363<=G9205 or G9192;
	G9367<=G9335 or G9331;
	G9388<=G9240 or G9223;
	G9392<=G9328 or G9324;
	G9509<=G9151 or G9125 or G9111;
	G9510<=G9125 or G9111;
	G9511<=G9151 or G9125 or G9111;
	G9512<=G9151 or G9125;
	G9515<=G9173 or G9151;
	G9516<=G9151 or G9125;
	G9519<=G9173 or G9151 or G9125;
	G9522<=G9173 or G9125;
	G9528<=G9151 or G9125 or G9111;
	G9536<=G9335 or G9331 or G9328 or G9324;
	G9557<=G9052 or G9030;
	G9560<=G9052 or G9030;
	G9563<=G9052 or G9030;
	G9566<=G9052 or G9030;
	G9569<=G9052 or G9030;
	G9573<=G9052 or G9030;
	G9579<=G9052 or G9030;
	G9624<=G9316 or G9313;
	G9673<=G9454 or G9292 or G9274;
	G9676<=G9454 or G9292 or G9274;
	G9680<=G9454 or G9292 or G9274;
	G9683<=G9454 or G9292 or G9274;
	G9686<=G9454 or G9292 or G9274;
	G9697<=G9665 or G9606 or I14822;
	G9700<=G9358 or G9667 or I14827;
	G9702<=G9365 or G9647 or I14831;
	G9704<=G9385 or G9605 or I14835;
	G9706<=G9644 or G9386 or G9591;
	G9708<=G9653 or G9389 or G9646;
	G9711<=G9660 or G9390 or G9359 or G9589;
	G9714<=G9664 or G9366 or G9654;
	G9722<=G9612 or G9643 or G9410 or I14855;
	G9723<=G9620 or G9652 or G9391 or I14858;
	G9724<=G9409 or G9419 or G9615;
	G9725<=G9642 or G9659 or G9616 or I14862;
	G9726<=G9411 or G9420 or G9489;
	G9727<=G9650 or G9663 or G9362 or I14866;
	G9728<=G9412 or G9422 or G9426;
	G9729<=G9618 or G9357 or G9656;
	G9730<=G9414 or G9425 or G9423;
	G9731<=G9641 or G9364 or G9387;
	G9734<=G9415 or G9428 or G9421;
	G9735<=G9649 or G9651 or G9384 or G9361;
	G9736<=G9430 or G9416;
	G9737<=G9657 or G9658 or G9655;
	G9738<=G9417 or G9447 or G9506;
	G9740<=G9418 or G9505;
	G9742<=G9173 or G9528;
	G9747<=G9173 or G9509;
	G9751<=G9515 or G9510;
	G9754<=G9173 or G9511;
	G9785<=G9010 or G8995 or G9388 or G9363;
	G9872<=G9617 or G9594 or G9750;
	G9873<=G9623 or G9599 or G9758;
	G9885<=G9739 or G9598 or G9662 or G9746;
	G9886<=G9607 or G9592 or G9759;
	G9888<=G9648 or G9608 or G9757;
	G9891<=G9741 or G9760;
	G9911<=G9846 or G9689;
	G9912<=G9847 or G9690;
	G9913<=G9849 or G9691;
	G9914<=G9851 or G9692;
	G9915<=G9853 or G9693;
	G9916<=G9855 or G9694;
	G9917<=G9856 or G9695;
	G9918<=G9858 or G9698;
	G9920<=G9860 or G9701;
	G9921<=G9862 or G9703;
	G9922<=G9864 or G9705;
	G9923<=G9865 or G9707;
	G9924<=G9866 or G9709;
	G9925<=G9867 or G9712;
	G9926<=G9868 or G9715;
	G9927<=G9869 or G9716;
	G9928<=G9870 or G9717;
	G9929<=G9871 or G9718;
	G9931<=G8931 or G9900;
	G9950<=G9901 or G9898 or G9779;
	G9951<=G9902 or G9899 or G9803;
	G9952<=G9944 or G9938 or G9817;
	G9953<=G9945 or G9939 or G9669;
	G9954<=G9946 or G9940 or G9781;
	G9955<=G9947 or G9941 or G9808;
	G9956<=G9948 or G9942 or G9815;
	G9957<=G9949 or G9943 or G9776;
	G9968<=I15171 or I15172;
	G9974<=I15176 or I15177;
	G9995<=I15199 or I15200;
	G10001<=I15204 or I15205;
	G10007<=I15209 or I15210;
	G10013<=I15214 or I15215;
	G10019<=I15219 or I15220;
	G10025<=I15224 or I15225;
	G10336<=G10230 or G9572;
	G10339<=G10232 or G9556;
	G10401<=G9317 or G10291;
	G10402<=G10295 or G9554;
	G10405<=G10297 or G9530;
	G10408<=G10298 or G9553;
	G10411<=G10299 or G9529;
	G10414<=G10300 or G9534;
	G10417<=G10301 or G9527;
	G10484<=G9317 or G10400;
	G10485<=G9317 or G10376;
	G10489<=G4961 or G10367;
	G10497<=G5052 or G10396;
	G10500<=G4157 or G10442;
	G10501<=G4161 or G10445;
	G10502<=G4169 or G10365;
	G10521<=I16148 or I16149;
	G10529<=I16160 or I16161;
	G10533<=G4933 or G10449;
	G10544<=G5511 or G10495;
	G10549<=G4951 or G10451;
	G10550<=G4942 or G10450;
	G10554<=G4097 or G10503;
	G10555<=G4103 or G10504;
	G10556<=G4115 or G10506;
	G10557<=G4123 or G10508;
	G10558<=G4126 or G10510;
	G10559<=G4141 or G10512;
	G10564<=G10560 or G7368;
	G10567<=G10514 or G7378;
	G10635<=G10622 or G7732;
	G10639<=G10623 or G7734;
	G10643<=G10624 or G7736;
	G10646<=G10625 or G7739;
	G10649<=G10626 or G7741;
	G10652<=G10627 or G7743;
	G10655<=G10561 or G7389;
	G10658<=G10595 or G7674;
	G10663<=G10237 or G10581;
	G10664<=G10240 or G10582;
	G10702<=G10562 or G3877;
	G10707<=G5545 or G10686;
	G10711<=G5547 or G10690;
	G10712<=G10662 or G9531;
	G10717<=G6235 or G10705;
	G10718<=G6238 or G10706;
	G10719<=G10303 or G10666;
	G10720<=G10304 or G10667;
	G10721<=G10306 or G10669;
	G10722<=G10308 or G10671;
	G10723<=G4952 or G10633;
	G10724<=G10312 or G10672;
	G10725<=G4962 or G10634;
	G10726<=G10316 or G10673;
	G10727<=G4969 or G10638;
	G10728<=G4973 or G10642;
	G10732<=G4358 or G10661;
	G10733<=G5227 or G10674;
	G10744<=G10600 or G10668 or I16427;
	G10765<=G5492 or G10680;
	G10767<=G5500 or G10681;
	G10770<=G5525 or G10682;
	G10771<=G5533 or G10684;
	G10773<=G5540 or G10685;
	G10776<=G5544 or G10758;
	G10791<=G6186 or G10762;
	G10793<=G6194 or G10763;
	G10795<=G6199 or G10764;
	G10797<=G6206 or G10766;
	G10798<=G6217 or G10768;
	G10799<=G6225 or G10769;
	G10800<=G6245 or G10772;
	G10805<=G10759 or G10760;
	G10807<=G10701 or G10761;
	G10855<=G6075 or G10736;
	G10856<=G6083 or G10737;
	G10857<=G6090 or G10738;
	G10858<=G5501 or G10741;
	G10859<=G5512 or G10742;
	G10860<=G5513 or G10743;
	G10861<=G5523 or G10745;
	G10862<=G5524 or G10746;
	G10863<=G5531 or G10750;
	G10864<=G5532 or G10751;
	G10865<=G5538 or G10752;
	G10866<=G5539 or G10753;
	G10898<=G4220 or G10777;
	G10923<=G10778 or G10715;
	G10936<=G5170 or G10808;
	G11058<=G10933 or G5280;
	G11201<=G11152 or G11011;
	G11217<=G11144 or G11005;
	G11219<=G11145 or G11006;
	G11221<=G11146 or G11007;
	G11223<=G11147 or G11008;
	G11225<=G11149 or G11009;
	G11227<=G11151 or G11010;
	G11229<=G11154 or G11012;
	G11231<=G11156 or G11013;
	G11232<=G11158 or G11015;
	G11233<=G11085 or G10946;
	G11246<=G11094 or G10948;
	G11247<=G11097 or G10949;
	G11249<=G6162 or G11143;
	G11252<=G11099 or G10969;
	G11256<=G11186 or G11018;
	G11257<=G11234 or G11019;
	G11258<=G11235 or G11020;
	G11259<=G11236 or G11021;
	G11260<=G11237 or G11022;
	G11261<=G11238 or G11023;
	G11262<=G11240 or G11024;
	G11263<=G11187 or G11025;
	G11264<=G11188 or G11026;
	G11265<=G11189 or G11027;
	G11266<=G11190 or G11028;
	G11267<=G11192 or G11029;
	G11268<=G11194 or G11030;
	G11269<=G11196 or G11031;
	G11270<=G11198 or G11032;
	G11275<=G11248 or G11148;
	G11278<=G11253 or G11150;
	G11280<=G11254 or G11153;
	G11285<=G11255 or G11161;
	G11286<=G10670 or G11209;
	G11288<=G11204 or G11070;
	G11293<=G11211 or G10818;
	G11294<=G6576 or G11210;
	G11298<=G11212 or G11087;
	G11300<=G11213 or G11091;
	G11303<=G11214 or G11092;
	G11305<=G11215 or G11093;
	G11306<=G11216 or G11095;
	G11308<=G11218 or G11098;
	G11310<=G11220 or G11100;
	G11312<=G11222 or G11101;
	G11314<=G11224 or G11102;
	G11316<=G11226 or G11103;
	G11318<=G11228 or G11104;
	G11321<=G11230 or G11105;
	G11324<=G11271 or G11164;
	G11325<=G11295 or G11165;
	G11326<=G11296 or G11166;
	G11327<=G11297 or G11167;
	G11328<=G11299 or G11168;
	G11329<=G11302 or G11169;
	G11330<=G11304 or G11170;
	G11331<=G11272 or G11171;
	G11332<=G11273 or G11172;
	G11333<=G11274 or G11173;
	G11334<=G11277 or G11174;
	G11335<=G11279 or G11175;
	G11336<=G11281 or G11176;
	G11337<=G11282 or G11177;
	G11338<=G11283 or G11178;
	G11430<=G11387 or G4006;
	G11443<=G7130 or G11407;
	G11478<=G6532 or G11455;
	G11481<=G6624 or G11458;
	G11482<=G6628 or G11459;
	G11483<=G6633 or G11460;
	G11484<=G6639 or G11461;
	G11485<=G6646 or G11462;
	G11486<=G6654 or G11463;
	G11487<=G6662 or G11464;
	G11488<=G6671 or G11465;
	G11579<=G5123 or G11551;
	G11580<=G11413 or G11544;
	G11602<=G11581 or G11552;
	G11603<=G11582 or G11553;
	G11604<=G11583 or G11554;
	G11605<=G11584 or G11555;
	G11606<=G11585 or G11556;
	G11607<=G11586 or G11557;
	G11608<=G11587 or G11558;
	G11609<=G11588 or G11559;
	G11610<=G11589 or G11560;
	G11612<=G11599 or G11590;
	G11613<=G11600 or G11591;
	G11615<=G11601 or G11592;
	G11624<=G11595 or G11571;
	G11625<=G6535 or G11597;
	G11647<=G6622 or G11637;
	I5351<=G1145 or G1141 or G1137 or G1133;
	I5352<=G1129 or G1125 or G1121 or G1117;
	I5357<=G1265 or G1260 or G1255 or G1250;
	I5358<=G1245 or G1240 or G1235 or G1275;
	I5363<=G1149 or G1153 or G1157 or G1160;
	I5366<=G1280 or G1284 or G1292 or G1296;
	I5570<=G416 or G411 or G406 or G401;
	I5571<=G396 or G391 or G386 or G426;
	I5576<=G431 or G435 or G440 or G444;
	I5599<=G516 or G511 or G506 or G501;
	I5600<=G496 or G491 or G486 or G481;
	I5626<=G521 or G525 or G530 or G534;
	I5629<=G845 or G841 or G837;
	I5649<=G1499 or G1486 or G1482;
	I5804<=G2111 or G2109 or G2106 or G2104;
	I5805<=G2102 or G2099 or G2096 or G2088;
	I6350<=G2445 or G2437 or G2433 or G2419;
	I6351<=G2405 or G2389 or G2380 or G2372;
	I14582<=G8995 or G9205 or G9192;
	I14585<=G8995 or G9205 or G9192;
	I14596<=G8995 or G9205 or G9192;
	I14602<=G8995 or G9205 or G9192;
	I14607<=G8995 or G9205 or G9192;
	I14751<=G8995 or G9205 or G9192;
	I14776<=G8995 or G9205 or G9192;
	I14779<=G8995 or G9205 or G9192;
	I14822<=G9597 or G9604 or G9582;
	I14827<=G9603 or G9614 or G9584;
	I14831<=G9613 or G9622 or G9586;
	I14835<=G9621 or G9645 or G9588;
	I14855<=G9583 or G9593 or G9601 or G9596;
	I14858<=G9585 or G9595 or G9610 or G9602;
	I14862<=G9587 or G9600 or G9611;
	I14866<=G9590 or G9609 or G9619;
	I15033<=G7853 or G9804 or G9624 or G9785;
	I15039<=G7853 or G9809 or G9624 or G9785;
	I15042<=G7853 or G9686 or G9624 or G9785;
	I15045<=G7853 or G9676 or G9624 or G9785;
	I15048<=G7853 or G9683 or G9624 or G9785;
	I15051<=G7853 or G9673 or G9624 or G9785;
	I15054<=G7853 or G9782 or G9624 or G9785;
	I15057<=G7853 or G9680 or G9624 or G9785;
	I15171<=G8175 or G9909 or G9896 or G9835;
	I15172<=G9843 or G9959 or G9861 or G9874;
	I15176<=G8176 or G9910 or G9897 or G9836;
	I15177<=G9844 or G9960 or G9863 or G9876;
	I15199<=G8167 or G9903 or G9932 or G9828;
	I15200<=G9837 or G9962 or G9848 or G9880;
	I15204<=G8168 or G9904 or G9933 or G9829;
	I15205<=G9838 or G9963 or G9850 or G9878;
	I15209<=G8169 or G9905 or G9934 or G9830;
	I15210<=G9839 or G9964 or G9852 or G9882;
	I15214<=G8170 or G9906 or G9935 or G9831;
	I15215<=G9840 or G9965 or G9854 or G9879;
	I15219<=G8172 or G9907 or G9936 or G9833;
	I15220<=G9841 or G9966 or G9857 or G9877;
	I15224<=G8174 or G9908 or G9937 or G9834;
	I15225<=G9842 or G9967 or G9859 or G9881;
	I16148<=G10386 or G10384 or G10476 or G10474;
	I16149<=G10472 or G10470 or G10468 or G10467;
	I16160<=G10394 or G10392 or G10482 or G10481;
	I16161<=G10479 or G10478 or G10477 or G10475;
	I16427<=G10683 or G10608 or G10604;
	G2459<= not (G1645 or G1642 or G1651 or G1648);
	G2478<= not (G1610 or G1737);
	G2791<= not (G2187 or G750);
	G2807<= not (G22 or G2320);
	G2862<= not (G2315 or G2305);
	G2863<= not (G2316 or G2309);
	G3107<= not (G2501 or G2499);
	G3118<= not (G2521 or G2514);
	G3462<= not (G2187 or G2795);
	G3879<= not (G3141 or G2354 or G2353);
	G4076<= not (G1707 or G2864);
	G4122<= not (G3291 or G2410 or G2538);
	G4218<= not (G3292 or G2593 or G3784 or G3776);
	G4227<= not (G3292 or G3793 or G2586 or G2579);
	G4234<= not (G3292 or G3793 or G2586 or G3776);
	G4251<= not (G3292 or G3793 or G3784 or G2579);
	G4259<= not (G3292 or G3793 or G3784 or G3776);
	G4267<= not (G3800 or G2593 or G2586 or G2579);
	G4276<= not (G4065 or G3261 or G2500);
	G4278<= not (G3800 or G2593 or G2586 or G3776);
	G4286<= not (G3800 or G2593 or G3784 or G2579);
	G4455<= not (G3543 or G3419 or G3408);
	G4572<= not (G3419 or G3408 or G3628);
	G4601<= not (G3077 or G2669 or G2662 or G3479);
	G4605<= not (G3077 or G2669 or G3485 or G2655);
	G4607<= not (G3077 or G2669 or G3485 or G3479);
	G4613<= not (G3077 or G3491 or G2662 or G2655);
	G4616<= not (G3077 or G3491 or G2662 or G3479);
	G4619<= not (G3077 or G3491 or G3485 or G2655);
	G4630<= not (G3077 or G3491 or G3485 or G3479);
	G4639<= not (G3501 or G2669 or G2662 or G2655);
	G4672<= not (G3501 or G2669 or G2662 or G3479);
	G4677<= not (G3501 or G2669 or G3485 or G2655);
	G4873<= not (G3292 or G2593 or G2586 or G3776);
	G4879<= not (G3292 or G2593 or G3784 or G2579);
	G4974<= not (G4502 or G3714);
	G5034<= not (G3524 or G4593);
	G5186<= not (G2047 or G4401);
	G5345<= not (G2754 or G4835);
	G5350<= not (G4163 or G4872);
	G5360<= not (G2071 or G4225);
	G5392<= not (G3369 or G4258);
	G5556<= not (G4787 or G2695 or G2299 or G2031);
	G5573<= not (G4117 or G4432);
	G5763<= not (G5350 or G5345);
	G5780<= not (G2112 or G4921);
	G5859<= not (G3362 or G4943);
	G5938<= not (G2764 or G4988);
	G5999<= not (G2753 or G4953);
	G6023<= not (G2763 or G4975);
	G6032<= not (G3430 or G5039);
	G6037<= not (G3305 or G5614);
	G6155<= not (G4974 or G2864);
	G6355<= not (G6032 or G6023);
	G6392<= not (G5859 or G5938);
	G8303<= not (G8209 or G4811);
	G9361<= not (G9010 or G9240 or G9223 or I14582);
	G9362<= not (G9010 or G9240 or G9223 or I14585);
	G9387<= not (G9010 or G9240 or G9223 or I14596);
	G9391<= not (G9010 or G9240 or G9223 or I14602);
	G9410<= not (G9010 or G9240 or G9223 or I14607);
	G9416<= not (G9052 or G9030);
	G9421<= not (G9052 or G9030);
	G9423<= not (G9052 or G9030);
	G9426<= not (G9052 or G9030);
	G9489<= not (G9052 or G9030);
	G9506<= not (G9052 or G9030);
	G9589<= not (G9125 or G9173 or G9151);
	G9591<= not (G9125 or G9151);
	G9605<= not (G9125 or G9111 or G9173 or G9151);
	G9606<= not (G9125 or G9111 or G9173 or G9151);
	G9615<= not (G9052 or G9030);
	G9616<= not (G9010 or G9240 or G9223 or I14751);
	G9646<= not (G9125 or G9151);
	G9647<= not (G9125 or G9111 or G9173 or G9151);
	G9654<= not (G9125 or G9173);
	G9655<= not (G9010 or G9240 or G9223 or I14776);
	G9656<= not (G9010 or G9240 or G9223 or I14779);
	G9667<= not (G9125 or G9111 or G9173 or G9151);
	G9669<= not (G9392 or G9367);
	G9746<= not (G9454 or G9274 or G9292);
	G9750<= not (G9454 or G9274 or G9292);
	G9757<= not (G9454 or G9274 or G9292);
	G9758<= not (G9454 or G9274 or G9292);
	G9759<= not (G9454 or G9274 or G9292);
	G9776<= not (G9392 or G9367);
	G9779<= not (G9392 or G9367);
	G9781<= not (G9392 or G9367);
	G9803<= not (G9392 or G9367);
	G9808<= not (G9392 or G9367);
	G9815<= not (G9392 or G9367);
	G9817<= not (G9392 or G9367);
	G9874<= not (G9519 or G9536 or G9579 or I15033);
	G9876<= not (G9522 or G9536 or G9576 or I15039);
	G9877<= not (G9512 or G9536 or G9569 or I15042);
	G9878<= not (G9754 or G9536 or G9560 or I15045);
	G9879<= not (G9747 or G9536 or G9566 or I15048);
	G9880<= not (G9751 or G9536 or G9557 or I15051);
	G9881<= not (G9516 or G9536 or G9573 or I15054);
	G9882<= not (G9742 or G9536 or G9563 or I15057);
	G10239<= not (G9317 or G10179);
	G10285<= not (G10276 or G3566);
	G10286<= not (G10271 or G3463);
	G10287<= not (G10275 or G3463);
	G10291<= not (G10247 or G3113);
	G10322<= not (G9317 or G10272);
	G10324<= not (G9317 or G10244);
	G10358<= not (G10226 or G4620);
	G10359<= not (G10227 or G4620);
	G10360<= not (G10277 or G3566);
	G10362<= not (G10228 or G3507);
	G10363<= not (G10355 or G3566);
	G10364<= not (G10327 or G3744);
	G10368<= not (G10342 or G3463);
	G10370<= not (G10343 or G3463);
	G10371<= not (G10344 or G3463);
	G10372<= not (G10345 or G3463);
	G10373<= not (G10346 or G3463);
	G10374<= not (G10347 or G3463);
	G10375<= not (G10288 or G3463);
	G10376<= not (G10323 or G3113);
	G10381<= not (G10310 or G2998);
	G10382<= not (G10314 or G2998);
	G10383<= not (G10318 or G2998);
	G10385<= not (G10321 or G2998);
	G10420<= not (G10329 or G3744);
	G10422<= not (G10289 or G4620);
	G10423<= not (G10290 or G4620);
	G10424<= not (G10292 or G4620);
	G10425<= not (G10293 or G4620);
	G10426<= not (G10294 or G4620);
	G10427<= not (G10296 or G4620);
	G10428<= not (G10335 or G4620);
	G10429<= not (G10326 or G3507);
	G10430<= not (G10349 or G3566);
	G10432<= not (G10350 or G3566);
	G10433<= not (G10330 or G3507);
	G10434<= not (G10352 or G3566);
	G10435<= not (G10332 or G3507);
	G10436<= not (G10354 or G3566);
	G10438<= not (G10356 or G3566);
	G10441<= not (G10351 or G3566);
	G10443<= not (G10353 or G3566);
	G10522<= not (G10486 or G10239);
	G10562<= not (G10483 or G10529);
	G10563<= not (G10539 or G10322);
	G10570<= not (G10542 or G10324);
	G10594<= not (G10480 or G10521);
	G10849<= not (G10739 or G3903);
	G11077<= not (G10970 or G10971);
	G11480<= not (G11456 or G4567);
end RTL;
